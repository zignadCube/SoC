-------------------------------------------------------------------------------
-- File         : nios_siso.vhd
-- Description  : nios_sios top level, automatically generated
-- Author       : Sabih Gerez, University of Twente
-- Creation date: August 7, 2015 (header added)
-------------------------------------------------------------------------------
-- $Rev: 1$
-- $Author: gerezsh$
-- $Date: Thu Sep 29 11:57:46 CEST 2022$
-- $Log$
-------------------------------------------------------------------------------

-- nios_siso.vhd

-- Generated using ACDS version 15.0 145

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios_siso is
  port (
    clk_clk              : in  std_logic                     := '0';             --           clk.clk
    clk_out_export       : out std_logic;                                        --       clk_out.export
    rst_reset_n          : in  std_logic                     := '0';             --           rst.reset_n
    siso_data_in_export  : in  std_logic_vector(15 downto 0) := (others => '0'); --  siso_data_in.export
    siso_data_out_export : out std_logic_vector(15 downto 0);                    -- siso_data_out.export
    siso_ready_export    : out std_logic;                                        --    siso_ready.export
    siso_req_export      : out std_logic;                                        --      siso_req.export
    stop_sim_export      : out std_logic                                         --      stop_sim.export
  );
end entity nios_siso;

architecture rtl of nios_siso is
  component gp_custom is
    port (
      clk           : in  std_logic                     := 'X';             -- clk
      resetn        : in  std_logic                     := 'X';             -- reset_n
      avs_addr      : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
      avs_read      : in  std_logic                     := 'X';             -- read
      avs_readdata  : out std_logic_vector(31 downto 0);                    -- readdata
      avs_write     : in  std_logic                     := 'X';             -- write
      avs_writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
      siso_req      : out std_logic;                                        -- export
      siso_ready    : out std_logic;                                        -- export
      siso_data_in  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- export
      siso_data_out : out std_logic_vector(15 downto 0);                    -- export
      clk_out       : out std_logic;                                        -- export
      stop_sim      : out std_logic                                         -- export
    );
  end component gp_custom;

  component nios_siso_jtag_uart_0 is
    port (
      clk            : in  std_logic                     := 'X';             -- clk
      rst_n          : in  std_logic                     := 'X';             -- reset_n
      av_chipselect  : in  std_logic                     := 'X';             -- chipselect
      av_address     : in  std_logic                     := 'X';             -- address
      av_read_n      : in  std_logic                     := 'X';             -- read_n
      av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
      av_write_n     : in  std_logic                     := 'X';             -- write_n
      av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
      av_waitrequest : out std_logic;                                        -- waitrequest
      av_irq         : out std_logic                                         -- irq
    );
  end component nios_siso_jtag_uart_0;

  component nios_siso_nios2_gen2 is
    port (
      clk                                 : in  std_logic                     := 'X';             -- clk
      reset_n                             : in  std_logic                     := 'X';             -- reset_n
      reset_req                           : in  std_logic                     := 'X';             -- reset_req
      d_address                           : out std_logic_vector(17 downto 0);                    -- address
      d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
      d_read                              : out std_logic;                                        -- read
      d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
      d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
      d_write                             : out std_logic;                                        -- write
      d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
      debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
      i_address                           : out std_logic_vector(17 downto 0);                    -- address
      i_read                              : out std_logic;                                        -- read
      i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
      i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
      irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
      debug_reset_request                 : out std_logic;                                        -- reset
      debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
      debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
      debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
      debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
      debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
      debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
      debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
      debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
      dummy_ci_port                       : out std_logic                                         -- readra
    );
  end component nios_siso_nios2_gen2;

  component nios_siso_on_chip_ra is
    port (
      clk        : in  std_logic                     := 'X';             -- clk
      address    : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
      clken      : in  std_logic                     := 'X';             -- clken
      chipselect : in  std_logic                     := 'X';             -- chipselect
      write      : in  std_logic                     := 'X';             -- write
      readdata   : out std_logic_vector(31 downto 0);                    -- readdata
      writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
      byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
      reset      : in  std_logic                     := 'X';             -- reset
      reset_req  : in  std_logic                     := 'X'              -- reset_req
    );
  end component nios_siso_on_chip_ra;

  component nios_siso_mm_interconnect_0 is
    port (
      clk_0_clk_clk                                : in  std_logic                     := 'X';             -- clk
      nios2_gen2_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
      nios2_gen2_data_master_address               : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
      nios2_gen2_data_master_waitrequest           : out std_logic;                                        -- waitrequest
      nios2_gen2_data_master_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
      nios2_gen2_data_master_read                  : in  std_logic                     := 'X';             -- read
      nios2_gen2_data_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
      nios2_gen2_data_master_write                 : in  std_logic                     := 'X';             -- write
      nios2_gen2_data_master_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
      nios2_gen2_data_master_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
      nios2_gen2_instruction_master_address        : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
      nios2_gen2_instruction_master_waitrequest    : out std_logic;                                        -- waitrequest
      nios2_gen2_instruction_master_read           : in  std_logic                     := 'X';             -- read
      nios2_gen2_instruction_master_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
      gp_custom_0_avalon_slave_address             : out std_logic_vector(5 downto 0);                     -- address
      gp_custom_0_avalon_slave_write               : out std_logic;                                        -- write
      gp_custom_0_avalon_slave_read                : out std_logic;                                        -- read
      gp_custom_0_avalon_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
      gp_custom_0_avalon_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
      jtag_uart_0_avalon_jtag_slave_address        : out std_logic_vector(0 downto 0);                     -- address
      jtag_uart_0_avalon_jtag_slave_write          : out std_logic;                                        -- write
      jtag_uart_0_avalon_jtag_slave_read           : out std_logic;                                        -- read
      jtag_uart_0_avalon_jtag_slave_readdata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
      jtag_uart_0_avalon_jtag_slave_writedata      : out std_logic_vector(31 downto 0);                    -- writedata
      jtag_uart_0_avalon_jtag_slave_waitrequest    : in  std_logic                     := 'X';             -- waitrequest
      jtag_uart_0_avalon_jtag_slave_chipselect     : out std_logic;                                        -- chipselect
      nios2_gen2_debug_mem_slave_address           : out std_logic_vector(8 downto 0);                     -- address
      nios2_gen2_debug_mem_slave_write             : out std_logic;                                        -- write
      nios2_gen2_debug_mem_slave_read              : out std_logic;                                        -- read
      nios2_gen2_debug_mem_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
      nios2_gen2_debug_mem_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
      nios2_gen2_debug_mem_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
      nios2_gen2_debug_mem_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
      nios2_gen2_debug_mem_slave_debugaccess       : out std_logic;                                        -- debugaccess
      on_chip_ra_s1_address                        : out std_logic_vector(13 downto 0);                    -- address
      on_chip_ra_s1_write                          : out std_logic;                                        -- write
      on_chip_ra_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
      on_chip_ra_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
      on_chip_ra_s1_byteenable                     : out std_logic_vector(3 downto 0);                     -- byteenable
      on_chip_ra_s1_chipselect                     : out std_logic;                                        -- chipselect
      on_chip_ra_s1_clken                          : out std_logic                                         -- clken
    );
  end component nios_siso_mm_interconnect_0;

  component nios_siso_irq_mapper is
    port (
      clk           : in  std_logic                     := 'X'; -- clk
      reset         : in  std_logic                     := 'X'; -- reset
      receiver0_irq : in  std_logic                     := 'X'; -- irq
      sender_irq    : out std_logic_vector(31 downto 0)         -- irq
    );
  end component nios_siso_irq_mapper;

  component altera_reset_controller is
    generic (
      NUM_RESET_INPUTS          : integer := 6;
      OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
      SYNC_DEPTH                : integer := 2;
      RESET_REQUEST_PRESENT     : integer := 0;
      RESET_REQ_WAIT_TIME       : integer := 1;
      MIN_RST_ASSERTION_TIME    : integer := 3;
      RESET_REQ_EARLY_DSRT_TIME : integer := 1;
      USE_RESET_REQUEST_IN0     : integer := 0;
      USE_RESET_REQUEST_IN1     : integer := 0;
      USE_RESET_REQUEST_IN2     : integer := 0;
      USE_RESET_REQUEST_IN3     : integer := 0;
      USE_RESET_REQUEST_IN4     : integer := 0;
      USE_RESET_REQUEST_IN5     : integer := 0;
      USE_RESET_REQUEST_IN6     : integer := 0;
      USE_RESET_REQUEST_IN7     : integer := 0;
      USE_RESET_REQUEST_IN8     : integer := 0;
      USE_RESET_REQUEST_IN9     : integer := 0;
      USE_RESET_REQUEST_IN10    : integer := 0;
      USE_RESET_REQUEST_IN11    : integer := 0;
      USE_RESET_REQUEST_IN12    : integer := 0;
      USE_RESET_REQUEST_IN13    : integer := 0;
      USE_RESET_REQUEST_IN14    : integer := 0;
      USE_RESET_REQUEST_IN15    : integer := 0;
      ADAPT_RESET_REQUEST       : integer := 0
    );
    port (
      reset_in0      : in  std_logic := 'X'; -- reset
      clk            : in  std_logic := 'X'; -- clk
      reset_out      : out std_logic;        -- reset
      reset_req      : out std_logic;        -- reset_req
      reset_req_in0  : in  std_logic := 'X'; -- reset_req
      reset_in1      : in  std_logic := 'X'; -- reset
      reset_req_in1  : in  std_logic := 'X'; -- reset_req
      reset_in2      : in  std_logic := 'X'; -- reset
      reset_req_in2  : in  std_logic := 'X'; -- reset_req
      reset_in3      : in  std_logic := 'X'; -- reset
      reset_req_in3  : in  std_logic := 'X'; -- reset_req
      reset_in4      : in  std_logic := 'X'; -- reset
      reset_req_in4  : in  std_logic := 'X'; -- reset_req
      reset_in5      : in  std_logic := 'X'; -- reset
      reset_req_in5  : in  std_logic := 'X'; -- reset_req
      reset_in6      : in  std_logic := 'X'; -- reset
      reset_req_in6  : in  std_logic := 'X'; -- reset_req
      reset_in7      : in  std_logic := 'X'; -- reset
      reset_req_in7  : in  std_logic := 'X'; -- reset_req
      reset_in8      : in  std_logic := 'X'; -- reset
      reset_req_in8  : in  std_logic := 'X'; -- reset_req
      reset_in9      : in  std_logic := 'X'; -- reset
      reset_req_in9  : in  std_logic := 'X'; -- reset_req
      reset_in10     : in  std_logic := 'X'; -- reset
      reset_req_in10 : in  std_logic := 'X'; -- reset_req
      reset_in11     : in  std_logic := 'X'; -- reset
      reset_req_in11 : in  std_logic := 'X'; -- reset_req
      reset_in12     : in  std_logic := 'X'; -- reset
      reset_req_in12 : in  std_logic := 'X'; -- reset_req
      reset_in13     : in  std_logic := 'X'; -- reset
      reset_req_in13 : in  std_logic := 'X'; -- reset_req
      reset_in14     : in  std_logic := 'X'; -- reset
      reset_req_in14 : in  std_logic := 'X'; -- reset_req
      reset_in15     : in  std_logic := 'X'; -- reset
      reset_req_in15 : in  std_logic := 'X'  -- reset_req
    );
  end component altera_reset_controller;

  signal nios2_gen2_data_master_readdata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_data_master_readdata -> nios2_gen2:d_readdata
  signal nios2_gen2_data_master_waitrequest                              : std_logic;                     -- mm_interconnect_0:nios2_gen2_data_master_waitrequest -> nios2_gen2:d_waitrequest
  signal nios2_gen2_data_master_debugaccess                              : std_logic;                     -- nios2_gen2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_data_master_debugaccess
  signal nios2_gen2_data_master_address                                  : std_logic_vector(17 downto 0); -- nios2_gen2:d_address -> mm_interconnect_0:nios2_gen2_data_master_address
  signal nios2_gen2_data_master_byteenable                               : std_logic_vector(3 downto 0);  -- nios2_gen2:d_byteenable -> mm_interconnect_0:nios2_gen2_data_master_byteenable
  signal nios2_gen2_data_master_read                                     : std_logic;                     -- nios2_gen2:d_read -> mm_interconnect_0:nios2_gen2_data_master_read
  signal nios2_gen2_data_master_write                                    : std_logic;                     -- nios2_gen2:d_write -> mm_interconnect_0:nios2_gen2_data_master_write
  signal nios2_gen2_data_master_writedata                                : std_logic_vector(31 downto 0); -- nios2_gen2:d_writedata -> mm_interconnect_0:nios2_gen2_data_master_writedata
  signal nios2_gen2_instruction_master_readdata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_instruction_master_readdata -> nios2_gen2:i_readdata
  signal nios2_gen2_instruction_master_waitrequest                       : std_logic;                     -- mm_interconnect_0:nios2_gen2_instruction_master_waitrequest -> nios2_gen2:i_waitrequest
  signal nios2_gen2_instruction_master_address                           : std_logic_vector(17 downto 0); -- nios2_gen2:i_address -> mm_interconnect_0:nios2_gen2_instruction_master_address
  signal nios2_gen2_instruction_master_read                              : std_logic;                     -- nios2_gen2:i_read -> mm_interconnect_0:nios2_gen2_instruction_master_read
  signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
  signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
  signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
  signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
  signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
  signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
  signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
  signal mm_interconnect_0_gp_custom_0_avalon_slave_readdata             : std_logic_vector(31 downto 0); -- gp_custom_0:avs_readdata -> mm_interconnect_0:gp_custom_0_avalon_slave_readdata
  signal mm_interconnect_0_gp_custom_0_avalon_slave_address              : std_logic_vector(5 downto 0);  -- mm_interconnect_0:gp_custom_0_avalon_slave_address -> gp_custom_0:avs_addr
  signal mm_interconnect_0_gp_custom_0_avalon_slave_read                 : std_logic;                     -- mm_interconnect_0:gp_custom_0_avalon_slave_read -> gp_custom_0:avs_read
  signal mm_interconnect_0_gp_custom_0_avalon_slave_write                : std_logic;                     -- mm_interconnect_0:gp_custom_0_avalon_slave_write -> gp_custom_0:avs_write
  signal mm_interconnect_0_gp_custom_0_avalon_slave_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:gp_custom_0_avalon_slave_writedata -> gp_custom_0:avs_writedata
  signal mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata           : std_logic_vector(31 downto 0); -- nios2_gen2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_debug_mem_slave_readdata
  signal mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest        : std_logic;                     -- nios2_gen2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_debug_mem_slave_waitrequest
  signal mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess        : std_logic;                     -- mm_interconnect_0:nios2_gen2_debug_mem_slave_debugaccess -> nios2_gen2:debug_mem_slave_debugaccess
  signal mm_interconnect_0_nios2_gen2_debug_mem_slave_address            : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_gen2_debug_mem_slave_address -> nios2_gen2:debug_mem_slave_address
  signal mm_interconnect_0_nios2_gen2_debug_mem_slave_read               : std_logic;                     -- mm_interconnect_0:nios2_gen2_debug_mem_slave_read -> nios2_gen2:debug_mem_slave_read
  signal mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_gen2_debug_mem_slave_byteenable -> nios2_gen2:debug_mem_slave_byteenable
  signal mm_interconnect_0_nios2_gen2_debug_mem_slave_write              : std_logic;                     -- mm_interconnect_0:nios2_gen2_debug_mem_slave_write -> nios2_gen2:debug_mem_slave_write
  signal mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_debug_mem_slave_writedata -> nios2_gen2:debug_mem_slave_writedata
  signal mm_interconnect_0_on_chip_ra_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:on_chip_ra_s1_chipselect -> on_chip_ra:chipselect
  signal mm_interconnect_0_on_chip_ra_s1_readdata                        : std_logic_vector(31 downto 0); -- on_chip_ra:readdata -> mm_interconnect_0:on_chip_ra_s1_readdata
  signal mm_interconnect_0_on_chip_ra_s1_address                         : std_logic_vector(13 downto 0); -- mm_interconnect_0:on_chip_ra_s1_address -> on_chip_ra:address
  signal mm_interconnect_0_on_chip_ra_s1_byteenable                      : std_logic_vector(3 downto 0);  -- mm_interconnect_0:on_chip_ra_s1_byteenable -> on_chip_ra:byteenable
  signal mm_interconnect_0_on_chip_ra_s1_write                           : std_logic;                     -- mm_interconnect_0:on_chip_ra_s1_write -> on_chip_ra:write
  signal mm_interconnect_0_on_chip_ra_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:on_chip_ra_s1_writedata -> on_chip_ra:writedata
  signal mm_interconnect_0_on_chip_ra_s1_clken                           : std_logic;                     -- mm_interconnect_0:on_chip_ra_s1_clken -> on_chip_ra:clken
  signal irq_mapper_receiver0_irq                                        : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
  signal nios2_gen2_irq_irq                                              : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_gen2:irq
  signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_gen2_reset_reset_bridge_in_reset_reset, on_chip_ra:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
  signal rst_controller_reset_out_reset_req                              : std_logic;                     -- rst_controller:reset_req -> [nios2_gen2:reset_req, on_chip_ra:reset_req, rst_translator:reset_req_in]
  signal rst_reset_n_ports_inv                                           : std_logic;                     -- rst_reset_n:inv -> rst_controller:reset_in0
  signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
  signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
  signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> [gp_custom_0:resetn, jtag_uart_0:rst_n, nios2_gen2:reset_n]

begin

  gp_custom_0 : component gp_custom
    port map (
      clk           => clk_clk,                                              --         clock.clk
      resetn        => rst_controller_reset_out_reset_ports_inv,             --    reset_sink.reset_n
      avs_addr      => mm_interconnect_0_gp_custom_0_avalon_slave_address,   --  avalon_slave.address
      avs_read      => mm_interconnect_0_gp_custom_0_avalon_slave_read,      --              .read
      avs_readdata  => mm_interconnect_0_gp_custom_0_avalon_slave_readdata,  --              .readdata
      avs_write     => mm_interconnect_0_gp_custom_0_avalon_slave_write,     --              .write
      avs_writedata => mm_interconnect_0_gp_custom_0_avalon_slave_writedata, --              .writedata
      siso_req      => siso_req_export,                                      --      siso_req.export
      siso_ready    => siso_ready_export,                                    --    siso_ready.export
      siso_data_in  => siso_data_in_export,                                  --  siso_data_in.export
      siso_data_out => siso_data_out_export,                                 -- siso_data_out.export
      clk_out       => clk_out_export,                                       --       clk_out.export
      stop_sim      => stop_sim_export                                       --      stop_sim.export
    );

  jtag_uart_0 : component nios_siso_jtag_uart_0
    port map (
      clk            => clk_clk,                                                         --               clk.clk
      rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
      av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
      av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
      av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
      av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
      av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
      av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
      av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
      av_irq         => irq_mapper_receiver0_irq                                         --               irq.irq
    );

  nios2_gen2 : component nios_siso_nios2_gen2
    port map (
      clk                                 => clk_clk,                                                  --                       clk.clk
      reset_n                             => rst_controller_reset_out_reset_ports_inv,                 --                     reset.reset_n
      reset_req                           => rst_controller_reset_out_reset_req,                       --                          .reset_req
      d_address                           => nios2_gen2_data_master_address,                           --               data_master.address
      d_byteenable                        => nios2_gen2_data_master_byteenable,                        --                          .byteenable
      d_read                              => nios2_gen2_data_master_read,                              --                          .read
      d_readdata                          => nios2_gen2_data_master_readdata,                          --                          .readdata
      d_waitrequest                       => nios2_gen2_data_master_waitrequest,                       --                          .waitrequest
      d_write                             => nios2_gen2_data_master_write,                             --                          .write
      d_writedata                         => nios2_gen2_data_master_writedata,                         --                          .writedata
      debug_mem_slave_debugaccess_to_roms => nios2_gen2_data_master_debugaccess,                       --                          .debugaccess
      i_address                           => nios2_gen2_instruction_master_address,                    --        instruction_master.address
      i_read                              => nios2_gen2_instruction_master_read,                       --                          .read
      i_readdata                          => nios2_gen2_instruction_master_readdata,                   --                          .readdata
      i_waitrequest                       => nios2_gen2_instruction_master_waitrequest,                --                          .waitrequest
      irq                                 => nios2_gen2_irq_irq,                                       --                       irq.irq
      debug_reset_request                 => open,                                                     --       debug_reset_request.reset
      debug_mem_slave_address             => mm_interconnect_0_nios2_gen2_debug_mem_slave_address,     --           debug_mem_slave.address
      debug_mem_slave_byteenable          => mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable,  --                          .byteenable
      debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess, --                          .debugaccess
      debug_mem_slave_read                => mm_interconnect_0_nios2_gen2_debug_mem_slave_read,        --                          .read
      debug_mem_slave_readdata            => mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata,    --                          .readdata
      debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest, --                          .waitrequest
      debug_mem_slave_write               => mm_interconnect_0_nios2_gen2_debug_mem_slave_write,       --                          .write
      debug_mem_slave_writedata           => mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata,   --                          .writedata
      dummy_ci_port                       => open                                                      -- custom_instruction_master.readra
    );

  on_chip_ra : component nios_siso_on_chip_ra
    port map (
      clk        => clk_clk,                                    --   clk1.clk
      address    => mm_interconnect_0_on_chip_ra_s1_address,    --     s1.address
      clken      => mm_interconnect_0_on_chip_ra_s1_clken,      --       .clken
      chipselect => mm_interconnect_0_on_chip_ra_s1_chipselect, --       .chipselect
      write      => mm_interconnect_0_on_chip_ra_s1_write,      --       .write
      readdata   => mm_interconnect_0_on_chip_ra_s1_readdata,   --       .readdata
      writedata  => mm_interconnect_0_on_chip_ra_s1_writedata,  --       .writedata
      byteenable => mm_interconnect_0_on_chip_ra_s1_byteenable, --       .byteenable
      reset      => rst_controller_reset_out_reset,             -- reset1.reset
      reset_req  => rst_controller_reset_out_reset_req          --       .reset_req
    );

  mm_interconnect_0 : component nios_siso_mm_interconnect_0
    port map (
      clk_0_clk_clk                                => clk_clk,                                                     --                              clk_0_clk.clk
      nios2_gen2_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                              -- nios2_gen2_reset_reset_bridge_in_reset.reset
      nios2_gen2_data_master_address               => nios2_gen2_data_master_address,                              --                 nios2_gen2_data_master.address
      nios2_gen2_data_master_waitrequest           => nios2_gen2_data_master_waitrequest,                          --                                       .waitrequest
      nios2_gen2_data_master_byteenable            => nios2_gen2_data_master_byteenable,                           --                                       .byteenable
      nios2_gen2_data_master_read                  => nios2_gen2_data_master_read,                                 --                                       .read
      nios2_gen2_data_master_readdata              => nios2_gen2_data_master_readdata,                             --                                       .readdata
      nios2_gen2_data_master_write                 => nios2_gen2_data_master_write,                                --                                       .write
      nios2_gen2_data_master_writedata             => nios2_gen2_data_master_writedata,                            --                                       .writedata
      nios2_gen2_data_master_debugaccess           => nios2_gen2_data_master_debugaccess,                          --                                       .debugaccess
      nios2_gen2_instruction_master_address        => nios2_gen2_instruction_master_address,                       --          nios2_gen2_instruction_master.address
      nios2_gen2_instruction_master_waitrequest    => nios2_gen2_instruction_master_waitrequest,                   --                                       .waitrequest
      nios2_gen2_instruction_master_read           => nios2_gen2_instruction_master_read,                          --                                       .read
      nios2_gen2_instruction_master_readdata       => nios2_gen2_instruction_master_readdata,                      --                                       .readdata
      gp_custom_0_avalon_slave_address             => mm_interconnect_0_gp_custom_0_avalon_slave_address,          --               gp_custom_0_avalon_slave.address
      gp_custom_0_avalon_slave_write               => mm_interconnect_0_gp_custom_0_avalon_slave_write,            --                                       .write
      gp_custom_0_avalon_slave_read                => mm_interconnect_0_gp_custom_0_avalon_slave_read,             --                                       .read
      gp_custom_0_avalon_slave_readdata            => mm_interconnect_0_gp_custom_0_avalon_slave_readdata,         --                                       .readdata
      gp_custom_0_avalon_slave_writedata           => mm_interconnect_0_gp_custom_0_avalon_slave_writedata,        --                                       .writedata
      jtag_uart_0_avalon_jtag_slave_address        => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,     --          jtag_uart_0_avalon_jtag_slave.address
      jtag_uart_0_avalon_jtag_slave_write          => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,       --                                       .write
      jtag_uart_0_avalon_jtag_slave_read           => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,        --                                       .read
      jtag_uart_0_avalon_jtag_slave_readdata       => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,    --                                       .readdata
      jtag_uart_0_avalon_jtag_slave_writedata      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,   --                                       .writedata
      jtag_uart_0_avalon_jtag_slave_waitrequest    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest, --                                       .waitrequest
      jtag_uart_0_avalon_jtag_slave_chipselect     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,  --                                       .chipselect
      nios2_gen2_debug_mem_slave_address           => mm_interconnect_0_nios2_gen2_debug_mem_slave_address,        --             nios2_gen2_debug_mem_slave.address
      nios2_gen2_debug_mem_slave_write             => mm_interconnect_0_nios2_gen2_debug_mem_slave_write,          --                                       .write
      nios2_gen2_debug_mem_slave_read              => mm_interconnect_0_nios2_gen2_debug_mem_slave_read,           --                                       .read
      nios2_gen2_debug_mem_slave_readdata          => mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata,       --                                       .readdata
      nios2_gen2_debug_mem_slave_writedata         => mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata,      --                                       .writedata
      nios2_gen2_debug_mem_slave_byteenable        => mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable,     --                                       .byteenable
      nios2_gen2_debug_mem_slave_waitrequest       => mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest,    --                                       .waitrequest
      nios2_gen2_debug_mem_slave_debugaccess       => mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess,    --                                       .debugaccess
      on_chip_ra_s1_address                        => mm_interconnect_0_on_chip_ra_s1_address,                     --                          on_chip_ra_s1.address
      on_chip_ra_s1_write                          => mm_interconnect_0_on_chip_ra_s1_write,                       --                                       .write
      on_chip_ra_s1_readdata                       => mm_interconnect_0_on_chip_ra_s1_readdata,                    --                                       .readdata
      on_chip_ra_s1_writedata                      => mm_interconnect_0_on_chip_ra_s1_writedata,                   --                                       .writedata
      on_chip_ra_s1_byteenable                     => mm_interconnect_0_on_chip_ra_s1_byteenable,                  --                                       .byteenable
      on_chip_ra_s1_chipselect                     => mm_interconnect_0_on_chip_ra_s1_chipselect,                  --                                       .chipselect
      on_chip_ra_s1_clken                          => mm_interconnect_0_on_chip_ra_s1_clken                        --                                       .clken
    );

  irq_mapper : component nios_siso_irq_mapper
    port map (
      clk           => clk_clk,                        --       clk.clk
      reset         => rst_controller_reset_out_reset, -- clk_reset.reset
      receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
      sender_irq    => nios2_gen2_irq_irq              --    sender.irq
    );

  rst_controller : component altera_reset_controller
    generic map (
      NUM_RESET_INPUTS          => 1,
      OUTPUT_RESET_SYNC_EDGES   => "deassert",
      SYNC_DEPTH                => 2,
      RESET_REQUEST_PRESENT     => 1,
      RESET_REQ_WAIT_TIME       => 1,
      MIN_RST_ASSERTION_TIME    => 3,
      RESET_REQ_EARLY_DSRT_TIME => 1,
      USE_RESET_REQUEST_IN0     => 0,
      USE_RESET_REQUEST_IN1     => 0,
      USE_RESET_REQUEST_IN2     => 0,
      USE_RESET_REQUEST_IN3     => 0,
      USE_RESET_REQUEST_IN4     => 0,
      USE_RESET_REQUEST_IN5     => 0,
      USE_RESET_REQUEST_IN6     => 0,
      USE_RESET_REQUEST_IN7     => 0,
      USE_RESET_REQUEST_IN8     => 0,
      USE_RESET_REQUEST_IN9     => 0,
      USE_RESET_REQUEST_IN10    => 0,
      USE_RESET_REQUEST_IN11    => 0,
      USE_RESET_REQUEST_IN12    => 0,
      USE_RESET_REQUEST_IN13    => 0,
      USE_RESET_REQUEST_IN14    => 0,
      USE_RESET_REQUEST_IN15    => 0,
      ADAPT_RESET_REQUEST       => 0
    )
    port map (
      reset_in0      => rst_reset_n_ports_inv,              -- reset_in0.reset
      clk            => clk_clk,                            --       clk.clk
      reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
      reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
      reset_req_in0  => '0',                                -- (terminated)
      reset_in1      => '0',                                -- (terminated)
      reset_req_in1  => '0',                                -- (terminated)
      reset_in2      => '0',                                -- (terminated)
      reset_req_in2  => '0',                                -- (terminated)
      reset_in3      => '0',                                -- (terminated)
      reset_req_in3  => '0',                                -- (terminated)
      reset_in4      => '0',                                -- (terminated)
      reset_req_in4  => '0',                                -- (terminated)
      reset_in5      => '0',                                -- (terminated)
      reset_req_in5  => '0',                                -- (terminated)
      reset_in6      => '0',                                -- (terminated)
      reset_req_in6  => '0',                                -- (terminated)
      reset_in7      => '0',                                -- (terminated)
      reset_req_in7  => '0',                                -- (terminated)
      reset_in8      => '0',                                -- (terminated)
      reset_req_in8  => '0',                                -- (terminated)
      reset_in9      => '0',                                -- (terminated)
      reset_req_in9  => '0',                                -- (terminated)
      reset_in10     => '0',                                -- (terminated)
      reset_req_in10 => '0',                                -- (terminated)
      reset_in11     => '0',                                -- (terminated)
      reset_req_in11 => '0',                                -- (terminated)
      reset_in12     => '0',                                -- (terminated)
      reset_req_in12 => '0',                                -- (terminated)
      reset_in13     => '0',                                -- (terminated)
      reset_req_in13 => '0',                                -- (terminated)
      reset_in14     => '0',                                -- (terminated)
      reset_req_in14 => '0',                                -- (terminated)
      reset_in15     => '0',                                -- (terminated)
      reset_req_in15 => '0'                                 -- (terminated)
    );

  rst_reset_n_ports_inv <= not rst_reset_n;

  mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

  mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

  rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of nios_siso
