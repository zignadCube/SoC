
library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

package CONV_PACK_gp_custom is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_gp_custom;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_gp_custom.all;

architecture flat_filter_none_5 of gp_custom is

   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component MUXB2DL
      port( A0, A1, SL : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AO21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN4D1
      port( A1, A2, A3, A4 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component AO22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2DL
      port( A0, A1, SL : in std_logic;  Z : out std_logic);
   end component;
   
   component AO31D1
      port( A1, A2, A3, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22M10D1
      port( B1, B2, A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3M1D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211D1
      port( A1, A2, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2D1
      port( A0, A1, SL : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFRPQ1
      port( D, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component DFERPQ1
      port( D, CEB, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFSPQ1
      port( D, CK, SB : in std_logic;  Q : out std_logic);
   end component;
   
   component OAI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI32D1
      port( A1, A2, A3, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   signal N62, N63, N64, avs_readdata_31_port, avs_readdata_30_port, 
      avs_readdata_29_port, avs_readdata_28_port, avs_readdata_27_port, 
      avs_readdata_26_port, avs_readdata_25_port, avs_readdata_24_port, 
      avs_readdata_23_port, avs_readdata_22_port, avs_readdata_21_port, 
      avs_readdata_20_port, avs_readdata_19_port, avs_readdata_18_port, 
      avs_readdata_17_port, avs_readdata_16_port, avs_readdata_15_port, 
      avs_readdata_14_port, avs_readdata_13_port, avs_readdata_12_port, 
      avs_readdata_11_port, avs_readdata_10_port, avs_readdata_9_port, 
      avs_readdata_8_port, avs_readdata_7_port, avs_readdata_6_port, 
      avs_readdata_5_port, avs_readdata_4_port, avs_readdata_3_port, 
      avs_readdata_2_port, avs_readdata_1_port, avs_readdata_0_port, 
      stop_sim_port, out_buf_255_port, out_buf_254_port, out_buf_253_port, 
      out_buf_252_port, out_buf_251_port, out_buf_250_port, out_buf_249_port, 
      out_buf_248_port, out_buf_247_port, out_buf_246_port, out_buf_245_port, 
      out_buf_244_port, out_buf_243_port, out_buf_242_port, out_buf_241_port, 
      out_buf_240_port, out_buf_239_port, out_buf_238_port, out_buf_237_port, 
      out_buf_236_port, out_buf_235_port, out_buf_234_port, out_buf_233_port, 
      out_buf_232_port, out_buf_231_port, out_buf_230_port, out_buf_229_port, 
      out_buf_228_port, out_buf_227_port, out_buf_226_port, out_buf_225_port, 
      out_buf_224_port, out_buf_223_port, out_buf_222_port, out_buf_221_port, 
      out_buf_220_port, out_buf_219_port, out_buf_218_port, out_buf_217_port, 
      out_buf_216_port, out_buf_215_port, out_buf_214_port, out_buf_213_port, 
      out_buf_212_port, out_buf_211_port, out_buf_210_port, out_buf_209_port, 
      out_buf_208_port, out_buf_207_port, out_buf_206_port, out_buf_205_port, 
      out_buf_204_port, out_buf_203_port, out_buf_202_port, out_buf_201_port, 
      out_buf_200_port, out_buf_199_port, out_buf_198_port, out_buf_197_port, 
      out_buf_196_port, out_buf_195_port, out_buf_194_port, out_buf_193_port, 
      out_buf_192_port, out_buf_191_port, out_buf_190_port, out_buf_189_port, 
      out_buf_188_port, out_buf_187_port, out_buf_186_port, out_buf_185_port, 
      out_buf_184_port, out_buf_183_port, out_buf_182_port, out_buf_181_port, 
      out_buf_180_port, out_buf_179_port, out_buf_178_port, out_buf_177_port, 
      out_buf_176_port, out_buf_175_port, out_buf_174_port, out_buf_173_port, 
      out_buf_172_port, out_buf_171_port, out_buf_170_port, out_buf_169_port, 
      out_buf_168_port, out_buf_167_port, out_buf_166_port, out_buf_165_port, 
      out_buf_164_port, out_buf_163_port, out_buf_162_port, out_buf_161_port, 
      out_buf_160_port, out_buf_159_port, out_buf_158_port, out_buf_157_port, 
      out_buf_156_port, out_buf_155_port, out_buf_154_port, out_buf_153_port, 
      out_buf_152_port, out_buf_151_port, out_buf_150_port, out_buf_149_port, 
      out_buf_148_port, out_buf_147_port, out_buf_146_port, out_buf_145_port, 
      out_buf_144_port, out_buf_143_port, out_buf_142_port, out_buf_141_port, 
      out_buf_140_port, out_buf_139_port, out_buf_138_port, out_buf_137_port, 
      out_buf_136_port, out_buf_135_port, out_buf_134_port, out_buf_133_port, 
      out_buf_132_port, out_buf_131_port, out_buf_130_port, out_buf_129_port, 
      out_buf_128_port, out_buf_127_port, out_buf_126_port, out_buf_125_port, 
      out_buf_124_port, out_buf_123_port, out_buf_122_port, out_buf_121_port, 
      out_buf_120_port, out_buf_119_port, out_buf_118_port, out_buf_117_port, 
      out_buf_116_port, out_buf_115_port, out_buf_114_port, out_buf_113_port, 
      out_buf_112_port, out_buf_111_port, out_buf_110_port, out_buf_109_port, 
      out_buf_108_port, out_buf_107_port, out_buf_106_port, out_buf_105_port, 
      out_buf_104_port, out_buf_103_port, out_buf_102_port, out_buf_101_port, 
      out_buf_100_port, out_buf_99_port, out_buf_98_port, out_buf_97_port, 
      out_buf_96_port, out_buf_95_port, out_buf_94_port, out_buf_93_port, 
      out_buf_92_port, out_buf_91_port, out_buf_90_port, out_buf_89_port, 
      out_buf_88_port, out_buf_87_port, out_buf_86_port, out_buf_85_port, 
      out_buf_84_port, out_buf_83_port, out_buf_82_port, out_buf_81_port, 
      out_buf_80_port, out_buf_79_port, out_buf_78_port, out_buf_77_port, 
      out_buf_76_port, out_buf_75_port, out_buf_74_port, out_buf_73_port, 
      out_buf_72_port, out_buf_71_port, out_buf_70_port, out_buf_69_port, 
      out_buf_68_port, out_buf_67_port, out_buf_66_port, out_buf_65_port, 
      out_buf_64_port, out_buf_63_port, out_buf_62_port, out_buf_61_port, 
      out_buf_60_port, out_buf_59_port, out_buf_58_port, out_buf_57_port, 
      out_buf_56_port, out_buf_55_port, out_buf_54_port, out_buf_53_port, 
      out_buf_52_port, out_buf_51_port, out_buf_50_port, out_buf_49_port, 
      out_buf_48_port, out_buf_47_port, out_buf_46_port, out_buf_45_port, 
      out_buf_44_port, out_buf_43_port, out_buf_42_port, out_buf_41_port, 
      out_buf_40_port, out_buf_39_port, out_buf_38_port, out_buf_37_port, 
      out_buf_36_port, out_buf_35_port, out_buf_34_port, out_buf_33_port, 
      out_buf_32_port, out_buf_31_port, out_buf_30_port, out_buf_29_port, 
      out_buf_28_port, out_buf_27_port, out_buf_26_port, out_buf_25_port, 
      out_buf_24_port, out_buf_23_port, out_buf_22_port, out_buf_21_port, 
      out_buf_20_port, out_buf_19_port, out_buf_18_port, out_buf_17_port, 
      out_buf_16_port, out_buf_15_port, out_buf_14_port, out_buf_13_port, 
      out_buf_12_port, out_buf_11_port, out_buf_10_port, out_buf_9_port, 
      out_buf_8_port, out_buf_7_port, out_buf_6_port, out_buf_5_port, 
      out_buf_4_port, out_buf_3_port, out_buf_2_port, out_buf_1_port, 
      out_buf_0_port, coeff_memory_0_31, coeff_memory_0_30, coeff_memory_0_29, 
      coeff_memory_0_28, coeff_memory_0_27, coeff_memory_0_26, 
      coeff_memory_0_25, coeff_memory_0_24, coeff_memory_0_23, 
      coeff_memory_0_22, coeff_memory_0_21, coeff_memory_0_20, 
      coeff_memory_0_19, coeff_memory_0_18, coeff_memory_0_17, 
      coeff_memory_0_16, coeff_memory_0_15, coeff_memory_0_14, 
      coeff_memory_0_13, coeff_memory_0_12, coeff_memory_0_11, 
      coeff_memory_0_10, coeff_memory_0_9, coeff_memory_0_8, coeff_memory_0_7, 
      coeff_memory_0_6, coeff_memory_0_5, coeff_memory_0_4, coeff_memory_0_3, 
      coeff_memory_0_2, coeff_memory_0_1, coeff_memory_0_0, coeff_memory_1_31, 
      coeff_memory_1_30, coeff_memory_1_29, coeff_memory_1_28, 
      coeff_memory_1_27, coeff_memory_1_26, coeff_memory_1_25, 
      coeff_memory_1_24, coeff_memory_1_23, coeff_memory_1_22, 
      coeff_memory_1_21, coeff_memory_1_20, coeff_memory_1_19, 
      coeff_memory_1_18, coeff_memory_1_17, coeff_memory_1_16, 
      coeff_memory_1_15, coeff_memory_1_14, coeff_memory_1_13, 
      coeff_memory_1_12, coeff_memory_1_11, coeff_memory_1_10, coeff_memory_1_9
      , coeff_memory_1_8, coeff_memory_1_7, coeff_memory_1_6, coeff_memory_1_5,
      coeff_memory_1_4, coeff_memory_1_3, coeff_memory_1_2, coeff_memory_1_1, 
      coeff_memory_1_0, coeff_memory_2_31, coeff_memory_2_30, coeff_memory_2_29
      , coeff_memory_2_28, coeff_memory_2_27, coeff_memory_2_26, 
      coeff_memory_2_25, coeff_memory_2_24, coeff_memory_2_23, 
      coeff_memory_2_22, coeff_memory_2_21, coeff_memory_2_20, 
      coeff_memory_2_19, coeff_memory_2_18, coeff_memory_2_17, 
      coeff_memory_2_16, coeff_memory_2_15, coeff_memory_2_14, 
      coeff_memory_2_13, coeff_memory_2_12, coeff_memory_2_11, 
      coeff_memory_2_10, coeff_memory_2_9, coeff_memory_2_8, coeff_memory_2_7, 
      coeff_memory_2_6, coeff_memory_2_5, coeff_memory_2_4, coeff_memory_2_3, 
      coeff_memory_2_2, coeff_memory_2_1, coeff_memory_2_0, coeff_memory_3_31, 
      coeff_memory_3_30, coeff_memory_3_29, coeff_memory_3_28, 
      coeff_memory_3_27, coeff_memory_3_26, coeff_memory_3_25, 
      coeff_memory_3_24, coeff_memory_3_23, coeff_memory_3_22, 
      coeff_memory_3_21, coeff_memory_3_20, coeff_memory_3_19, 
      coeff_memory_3_18, coeff_memory_3_17, coeff_memory_3_16, 
      coeff_memory_3_15, coeff_memory_3_14, coeff_memory_3_13, 
      coeff_memory_3_12, coeff_memory_3_11, coeff_memory_3_10, coeff_memory_3_9
      , coeff_memory_3_8, coeff_memory_3_7, coeff_memory_3_6, coeff_memory_3_5,
      coeff_memory_3_4, coeff_memory_3_3, coeff_memory_3_2, coeff_memory_3_1, 
      coeff_memory_3_0, coeff_memory_4_31, coeff_memory_4_30, coeff_memory_4_29
      , coeff_memory_4_28, coeff_memory_4_27, coeff_memory_4_26, 
      coeff_memory_4_25, coeff_memory_4_24, coeff_memory_4_23, 
      coeff_memory_4_22, coeff_memory_4_21, coeff_memory_4_20, 
      coeff_memory_4_19, coeff_memory_4_18, coeff_memory_4_17, 
      coeff_memory_4_16, coeff_memory_4_15, coeff_memory_4_14, 
      coeff_memory_4_13, coeff_memory_4_12, coeff_memory_4_11, 
      coeff_memory_4_10, coeff_memory_4_9, coeff_memory_4_8, coeff_memory_4_7, 
      coeff_memory_4_6, coeff_memory_4_5, coeff_memory_4_4, coeff_memory_4_3, 
      coeff_memory_4_2, coeff_memory_4_1, coeff_memory_4_0, 
      operand_regs_255_port, operand_regs_254_port, operand_regs_253_port, 
      operand_regs_252_port, operand_regs_251_port, operand_regs_250_port, 
      operand_regs_249_port, operand_regs_248_port, operand_regs_247_port, 
      operand_regs_246_port, operand_regs_245_port, operand_regs_244_port, 
      operand_regs_243_port, operand_regs_242_port, operand_regs_241_port, 
      operand_regs_240_port, operand_regs_239_port, operand_regs_238_port, 
      operand_regs_237_port, operand_regs_236_port, operand_regs_235_port, 
      operand_regs_234_port, operand_regs_233_port, operand_regs_232_port, 
      operand_regs_231_port, operand_regs_230_port, operand_regs_229_port, 
      operand_regs_228_port, operand_regs_227_port, operand_regs_226_port, 
      operand_regs_225_port, operand_regs_224_port, operand_regs_223_port, 
      operand_regs_222_port, operand_regs_221_port, operand_regs_220_port, 
      operand_regs_219_port, operand_regs_218_port, operand_regs_217_port, 
      operand_regs_216_port, operand_regs_215_port, operand_regs_214_port, 
      operand_regs_213_port, operand_regs_212_port, operand_regs_211_port, 
      operand_regs_210_port, operand_regs_209_port, operand_regs_208_port, 
      operand_regs_207_port, operand_regs_206_port, operand_regs_205_port, 
      operand_regs_204_port, operand_regs_203_port, operand_regs_202_port, 
      operand_regs_201_port, operand_regs_200_port, operand_regs_199_port, 
      operand_regs_198_port, operand_regs_197_port, operand_regs_196_port, 
      operand_regs_195_port, operand_regs_194_port, operand_regs_193_port, 
      operand_regs_192_port, operand_regs_191_port, operand_regs_190_port, 
      operand_regs_189_port, operand_regs_188_port, operand_regs_187_port, 
      operand_regs_186_port, operand_regs_185_port, operand_regs_184_port, 
      operand_regs_183_port, operand_regs_182_port, operand_regs_181_port, 
      operand_regs_180_port, operand_regs_179_port, operand_regs_178_port, 
      operand_regs_177_port, operand_regs_176_port, operand_regs_175_port, 
      operand_regs_174_port, operand_regs_173_port, operand_regs_172_port, 
      operand_regs_171_port, operand_regs_170_port, operand_regs_169_port, 
      operand_regs_168_port, operand_regs_167_port, operand_regs_166_port, 
      operand_regs_165_port, operand_regs_164_port, operand_regs_163_port, 
      operand_regs_162_port, operand_regs_161_port, operand_regs_160_port, 
      operand_regs_159_port, operand_regs_158_port, operand_regs_157_port, 
      operand_regs_156_port, operand_regs_155_port, operand_regs_154_port, 
      operand_regs_153_port, operand_regs_152_port, operand_regs_151_port, 
      operand_regs_150_port, operand_regs_149_port, operand_regs_148_port, 
      operand_regs_147_port, operand_regs_146_port, operand_regs_145_port, 
      operand_regs_144_port, operand_regs_143_port, operand_regs_142_port, 
      operand_regs_141_port, operand_regs_140_port, operand_regs_139_port, 
      operand_regs_138_port, operand_regs_137_port, operand_regs_136_port, 
      operand_regs_135_port, operand_regs_134_port, operand_regs_133_port, 
      operand_regs_132_port, operand_regs_131_port, operand_regs_130_port, 
      operand_regs_129_port, operand_regs_128_port, operand_regs_127_port, 
      operand_regs_126_port, operand_regs_125_port, operand_regs_124_port, 
      operand_regs_123_port, operand_regs_122_port, operand_regs_121_port, 
      operand_regs_120_port, operand_regs_119_port, operand_regs_118_port, 
      operand_regs_117_port, operand_regs_116_port, operand_regs_115_port, 
      operand_regs_114_port, operand_regs_113_port, operand_regs_112_port, 
      operand_regs_111_port, operand_regs_110_port, operand_regs_109_port, 
      operand_regs_108_port, operand_regs_107_port, operand_regs_106_port, 
      operand_regs_105_port, operand_regs_104_port, operand_regs_103_port, 
      operand_regs_102_port, operand_regs_101_port, operand_regs_100_port, 
      operand_regs_99_port, operand_regs_98_port, operand_regs_97_port, 
      operand_regs_96_port, operand_regs_95_port, operand_regs_94_port, 
      operand_regs_93_port, operand_regs_92_port, operand_regs_91_port, 
      operand_regs_90_port, operand_regs_89_port, operand_regs_88_port, 
      operand_regs_87_port, operand_regs_86_port, operand_regs_85_port, 
      operand_regs_84_port, operand_regs_83_port, operand_regs_82_port, 
      operand_regs_81_port, operand_regs_80_port, operand_regs_79_port, 
      operand_regs_78_port, operand_regs_77_port, operand_regs_76_port, 
      operand_regs_75_port, operand_regs_74_port, operand_regs_73_port, 
      operand_regs_72_port, operand_regs_71_port, operand_regs_70_port, 
      operand_regs_69_port, operand_regs_68_port, operand_regs_67_port, 
      operand_regs_66_port, operand_regs_65_port, operand_regs_64_port, 
      operand_regs_63_port, operand_regs_62_port, operand_regs_61_port, 
      operand_regs_60_port, operand_regs_59_port, operand_regs_58_port, 
      operand_regs_57_port, operand_regs_56_port, operand_regs_55_port, 
      operand_regs_54_port, operand_regs_53_port, operand_regs_52_port, 
      operand_regs_51_port, operand_regs_50_port, operand_regs_49_port, 
      operand_regs_48_port, operand_regs_47_port, operand_regs_46_port, 
      operand_regs_45_port, operand_regs_44_port, operand_regs_43_port, 
      operand_regs_42_port, operand_regs_41_port, operand_regs_40_port, 
      operand_regs_39_port, operand_regs_38_port, operand_regs_37_port, 
      operand_regs_36_port, operand_regs_35_port, operand_regs_34_port, 
      operand_regs_33_port, operand_regs_32_port, operand_regs_31_port, 
      operand_regs_30_port, operand_regs_29_port, operand_regs_28_port, 
      operand_regs_27_port, operand_regs_26_port, operand_regs_25_port, 
      operand_regs_24_port, operand_regs_23_port, operand_regs_22_port, 
      operand_regs_21_port, operand_regs_20_port, operand_regs_19_port, 
      operand_regs_18_port, operand_regs_17_port, operand_regs_16_port, 
      operand_regs_15_port, operand_regs_14_port, operand_regs_13_port, 
      operand_regs_12_port, operand_regs_11_port, operand_regs_10_port, 
      operand_regs_9_port, operand_regs_8_port, operand_regs_7_port, 
      operand_regs_6_port, operand_regs_5_port, operand_regs_4_port, 
      operand_regs_3_port, operand_regs_2_port, operand_regs_1_port, 
      operand_regs_0_port, in_trigger, out_trigger, coeff_load, operand_load, 
      read_comp_res, filt_mult_inputs, N66, comp_res_159_port, 
      comp_res_158_port, comp_res_157_port, comp_res_156_port, 
      comp_res_155_port, comp_res_154_port, comp_res_153_port, 
      comp_res_152_port, comp_res_151_port, comp_res_150_port, 
      comp_res_149_port, comp_res_148_port, comp_res_147_port, 
      comp_res_146_port, comp_res_145_port, comp_res_144_port, 
      comp_res_143_port, comp_res_142_port, comp_res_141_port, 
      comp_res_140_port, comp_res_139_port, comp_res_138_port, 
      comp_res_137_port, comp_res_136_port, comp_res_135_port, 
      comp_res_134_port, comp_res_133_port, comp_res_132_port, 
      comp_res_131_port, comp_res_130_port, comp_res_129_port, 
      comp_res_128_port, comp_res_127_port, comp_res_126_port, 
      comp_res_125_port, comp_res_124_port, comp_res_123_port, 
      comp_res_122_port, comp_res_121_port, comp_res_120_port, 
      comp_res_119_port, comp_res_118_port, comp_res_117_port, 
      comp_res_116_port, comp_res_115_port, comp_res_114_port, 
      comp_res_113_port, comp_res_112_port, comp_res_111_port, 
      comp_res_110_port, comp_res_109_port, comp_res_108_port, 
      comp_res_107_port, comp_res_106_port, comp_res_105_port, 
      comp_res_104_port, comp_res_103_port, comp_res_102_port, 
      comp_res_101_port, comp_res_100_port, comp_res_99_port, comp_res_98_port,
      comp_res_97_port, comp_res_96_port, comp_res_95_port, comp_res_94_port, 
      comp_res_93_port, comp_res_92_port, comp_res_91_port, comp_res_90_port, 
      comp_res_89_port, comp_res_88_port, comp_res_87_port, comp_res_86_port, 
      comp_res_85_port, comp_res_84_port, comp_res_83_port, comp_res_82_port, 
      comp_res_81_port, comp_res_80_port, comp_res_79_port, comp_res_78_port, 
      comp_res_77_port, comp_res_76_port, comp_res_75_port, comp_res_74_port, 
      comp_res_73_port, comp_res_72_port, comp_res_71_port, comp_res_70_port, 
      comp_res_69_port, comp_res_68_port, comp_res_67_port, comp_res_66_port, 
      comp_res_65_port, comp_res_64_port, comp_res_63_port, comp_res_62_port, 
      comp_res_61_port, comp_res_60_port, comp_res_59_port, comp_res_58_port, 
      comp_res_57_port, comp_res_56_port, comp_res_55_port, comp_res_54_port, 
      comp_res_53_port, comp_res_52_port, comp_res_51_port, comp_res_50_port, 
      comp_res_49_port, comp_res_48_port, comp_res_47_port, comp_res_46_port, 
      comp_res_45_port, comp_res_44_port, comp_res_43_port, comp_res_42_port, 
      comp_res_41_port, comp_res_40_port, comp_res_39_port, comp_res_38_port, 
      comp_res_37_port, comp_res_36_port, comp_res_35_port, comp_res_34_port, 
      comp_res_33_port, comp_res_32_port, comp_res_31_port, comp_res_30_port, 
      comp_res_29_port, comp_res_28_port, comp_res_27_port, comp_res_26_port, 
      comp_res_25_port, comp_res_24_port, comp_res_23_port, comp_res_22_port, 
      comp_res_21_port, comp_res_20_port, comp_res_19_port, comp_res_18_port, 
      comp_res_17_port, comp_res_16_port, comp_res_15_port, comp_res_14_port, 
      comp_res_13_port, comp_res_12_port, comp_res_11_port, comp_res_10_port, 
      comp_res_9_port, comp_res_8_port, comp_res_7_port, comp_res_6_port, 
      comp_res_5_port, comp_res_4_port, comp_res_3_port, comp_res_2_port, 
      comp_res_1_port, comp_res_0_port, N1978, N1979, N1980, N1981, N1982, 
      N1983, N1984, N1985, N1986, N1987, N1988, N1989, N1990, N1991, N1992, 
      N1993, N1994, N1995, N1996, N1997, N1998, N1999, N2000, N2001, N2002, 
      N2003, N2004, N2005, N2006, N2007, N2008, N2009, in_buf_255_port, 
      in_buf_254_port, in_buf_253_port, in_buf_252_port, in_buf_251_port, 
      in_buf_250_port, in_buf_249_port, in_buf_248_port, in_buf_247_port, 
      in_buf_246_port, in_buf_245_port, in_buf_244_port, in_buf_243_port, 
      in_buf_242_port, in_buf_241_port, in_buf_240_port, in_buf_239_port, 
      in_buf_238_port, in_buf_237_port, in_buf_236_port, in_buf_235_port, 
      in_buf_234_port, in_buf_233_port, in_buf_232_port, in_buf_231_port, 
      in_buf_230_port, in_buf_229_port, in_buf_228_port, in_buf_227_port, 
      in_buf_226_port, in_buf_225_port, in_buf_224_port, in_buf_223_port, 
      in_buf_222_port, in_buf_221_port, in_buf_220_port, in_buf_219_port, 
      in_buf_218_port, in_buf_217_port, in_buf_216_port, in_buf_215_port, 
      in_buf_214_port, in_buf_213_port, in_buf_212_port, in_buf_211_port, 
      in_buf_210_port, in_buf_209_port, in_buf_208_port, in_buf_207_port, 
      in_buf_206_port, in_buf_205_port, in_buf_204_port, in_buf_203_port, 
      in_buf_202_port, in_buf_201_port, in_buf_200_port, in_buf_199_port, 
      in_buf_198_port, in_buf_197_port, in_buf_196_port, in_buf_195_port, 
      in_buf_194_port, in_buf_193_port, in_buf_192_port, in_buf_191_port, 
      in_buf_190_port, in_buf_189_port, in_buf_188_port, in_buf_187_port, 
      in_buf_186_port, in_buf_185_port, in_buf_184_port, in_buf_183_port, 
      in_buf_182_port, in_buf_181_port, in_buf_180_port, in_buf_179_port, 
      in_buf_178_port, in_buf_177_port, in_buf_176_port, in_buf_175_port, 
      in_buf_174_port, in_buf_173_port, in_buf_172_port, in_buf_171_port, 
      in_buf_170_port, in_buf_169_port, in_buf_168_port, in_buf_167_port, 
      in_buf_166_port, in_buf_165_port, in_buf_164_port, in_buf_163_port, 
      in_buf_162_port, in_buf_161_port, in_buf_160_port, in_buf_159_port, 
      in_buf_158_port, in_buf_157_port, in_buf_156_port, in_buf_155_port, 
      in_buf_154_port, in_buf_153_port, in_buf_152_port, in_buf_151_port, 
      in_buf_150_port, in_buf_149_port, in_buf_148_port, in_buf_147_port, 
      in_buf_146_port, in_buf_145_port, in_buf_144_port, in_buf_143_port, 
      in_buf_142_port, in_buf_141_port, in_buf_140_port, in_buf_139_port, 
      in_buf_138_port, in_buf_137_port, in_buf_136_port, in_buf_135_port, 
      in_buf_134_port, in_buf_133_port, in_buf_132_port, in_buf_131_port, 
      in_buf_130_port, in_buf_129_port, in_buf_128_port, in_buf_127_port, 
      in_buf_126_port, in_buf_125_port, in_buf_124_port, in_buf_123_port, 
      in_buf_122_port, in_buf_121_port, in_buf_120_port, in_buf_119_port, 
      in_buf_118_port, in_buf_117_port, in_buf_116_port, in_buf_115_port, 
      in_buf_114_port, in_buf_113_port, in_buf_112_port, in_buf_111_port, 
      in_buf_110_port, in_buf_109_port, in_buf_108_port, in_buf_107_port, 
      in_buf_106_port, in_buf_105_port, in_buf_104_port, in_buf_103_port, 
      in_buf_102_port, in_buf_101_port, in_buf_100_port, in_buf_99_port, 
      in_buf_98_port, in_buf_97_port, in_buf_96_port, in_buf_95_port, 
      in_buf_94_port, in_buf_93_port, in_buf_92_port, in_buf_91_port, 
      in_buf_90_port, in_buf_89_port, in_buf_88_port, in_buf_87_port, 
      in_buf_86_port, in_buf_85_port, in_buf_84_port, in_buf_83_port, 
      in_buf_82_port, in_buf_81_port, in_buf_80_port, in_buf_79_port, 
      in_buf_78_port, in_buf_77_port, in_buf_76_port, in_buf_75_port, 
      in_buf_74_port, in_buf_73_port, in_buf_72_port, in_buf_71_port, 
      in_buf_70_port, in_buf_69_port, in_buf_68_port, in_buf_67_port, 
      in_buf_66_port, in_buf_65_port, in_buf_64_port, in_buf_63_port, 
      in_buf_62_port, in_buf_61_port, in_buf_60_port, in_buf_59_port, 
      in_buf_58_port, in_buf_57_port, in_buf_56_port, in_buf_55_port, 
      in_buf_54_port, in_buf_53_port, in_buf_52_port, in_buf_51_port, 
      in_buf_50_port, in_buf_49_port, in_buf_48_port, in_buf_47_port, 
      in_buf_46_port, in_buf_45_port, in_buf_44_port, in_buf_43_port, 
      in_buf_42_port, in_buf_41_port, in_buf_40_port, in_buf_39_port, 
      in_buf_38_port, in_buf_37_port, in_buf_36_port, in_buf_35_port, 
      in_buf_34_port, in_buf_33_port, in_buf_32_port, in_buf_31_port, 
      in_buf_30_port, in_buf_29_port, in_buf_28_port, in_buf_27_port, 
      in_buf_26_port, in_buf_25_port, in_buf_24_port, in_buf_23_port, 
      in_buf_22_port, in_buf_21_port, in_buf_20_port, in_buf_19_port, 
      in_buf_18_port, in_buf_17_port, in_buf_16_port, in_buf_15_port, 
      in_buf_14_port, in_buf_13_port, in_buf_12_port, in_buf_11_port, 
      in_buf_10_port, in_buf_9_port, in_buf_8_port, in_buf_7_port, 
      in_buf_6_port, in_buf_5_port, in_buf_4_port, in_buf_3_port, in_buf_2_port
      , in_buf_1_port, in_buf_0_port, N2010, N2011, N2012, N2013, N2014, N2015,
      N2016, N2017, N2018, N2019, N2020, N2021, N2022, N2023, N2024, N2025, 
      N2026, N2027, N2028, N2029, N2030, N2031, N2032, N2033, N2034, N2035, 
      N2036, N2037, N2038, N2039, N2040, N2041, in_busy, out_busy, 
      in_counter_2_port, in_counter_1_port, in_counter_0_port, odd, odd1, N2850
      , N2851, N2852, N2853, N2854, N2855, N2856, N2857, N2858, N2859, N2860, 
      N2861, N2862, N2863, N2864, N2865, N2867, N2868, N2869, N2870, N2871, 
      N2872, N2873, N2874, N2875, N2876, N2877, N2878, N2879, N2880, N2881, 
      N2882, N2888, N2889, N2890, N2891, N2892, N2893, N2894, N2895, N2896, 
      N2897, N2898, N2899, N2900, N2901, N2902, N2903, N2913, N2914, N2915, 
      N2916, N2917, N2918, N2919, N2920, N2921, N2922, N2923, N2924, N2925, 
      N2926, N2927, N2928, N2929, N2930, N2931, N2932, N2933, N2934, N2935, 
      N2936, N2937, N2938, N2939, N2940, N2941, N2942, N2943, N2944, N2945, 
      N2946, N2947, N2948, N2949, N2950, N2951, N2952, N2953, N2954, N2955, 
      N2956, N2957, N2958, N2959, N2960, N2961, N2962, N2963, N2964, N2965, 
      N2966, N2967, N2968, N2969, N2970, N2971, N2972, N2973, N2974, N2975, 
      N2976, N2977, N2978, N2979, N2980, N2981, N2982, N2983, N2984, N2985, 
      N2986, N2987, N2988, N2989, N2990, N2991, N2992, N2993, N2994, N2995, 
      N2996, N2997, N2998, N2999, N3000, N3001, N3002, N3003, N3004, N3005, 
      N3006, N3007, N3008, N3009, N3010, N3011, N3012, N3013, N3014, N3015, 
      N3016, N3017, N3018, N3019, N3020, N3021, N3022, N3023, N3024, N3025, 
      N3026, N3027, N3028, N3029, N3030, N3031, N3032, N3033, N3034, N3035, 
      N3036, N3037, N3038, N3039, N3040, N3041, N3042, N3043, N3044, N3045, 
      N3046, N3047, N3048, N3049, N3050, N3051, N3052, N3053, N3054, N3055, 
      N3056, N3057, N3058, N3059, N3060, N3061, N3062, N3063, N3064, N3065, 
      N3066, N3067, N3068, N3069, N3070, N3071, N3072, N3073, N3074, N3075, 
      N3076, N3077, N3078, N3079, N3080, N3081, N3082, N3083, N3084, N3085, 
      N3086, N3087, N3088, N3089, N3090, N3091, N3092, N3093, N3094, N3095, 
      N3096, N3097, N3098, N3099, N3100, N3101, N3102, N3103, N3104, N3105, 
      N3106, N3107, N3108, N3109, N3110, N3111, N3112, N3113, N3114, N3115, 
      N3116, N3117, N3118, N3119, N3120, N3121, N3122, N3123, N3124, N3125, 
      N3126, N3127, N3128, N3129, N3130, N3131, N3132, N3133, N3134, N3135, 
      N3136, N3137, N3138, N3139, N3140, N3141, N3142, N3143, N3144, N3145, 
      N3146, N3147, N3148, N3149, N3150, N3151, N3152, N3153, N3154, N3155, 
      N3156, N3157, N3158, N3159, N3160, N3161, N3162, N3163, N3164, N3165, 
      N3166, N3167, N3168, N3233, N3234, N3235, N3236, N3237, N3238, N3239, 
      N3240, N3241, N3242, N3243, N3244, N3245, N3246, N3247, N3248, N3249, 
      N3250, N3251, N3252, N3253, N3254, N3255, N3256, N3257, N3258, N3259, 
      N3260, N3261, N3262, N3263, N3264, N3265, N3266, N3267, N3268, N3269, 
      N3270, N3271, N3272, N3273, N3274, N3275, N3276, N3277, N3278, N3279, 
      N3280, N3281, N3282, N3283, N3284, N3285, N3286, N3287, N3288, N3289, 
      N3290, N3291, N3292, N3293, N3294, N3295, N3296, N3297, N3298, N3299, 
      N3300, N3301, N3302, N3303, N3304, N3305, N3306, N3307, N3308, N3309, 
      N3310, N3311, N3312, N3313, N3314, N3315, N3316, N3317, N3318, N3319, 
      N3320, N3321, N3322, N3323, N3324, N3325, N3326, N3327, N3328, N3329, 
      N3330, N3331, N3332, N3333, N3334, N3335, N3336, N3337, N3338, N3339, 
      N3340, N3341, N3342, N3343, N3344, N3345, N3346, N3347, N3348, N3349, 
      N3350, N3351, N3352, N3353, N3354, N3355, N3356, N3357, N3358, N3359, 
      N3360, N3361, N3362, N3363, N3364, N3365, N3366, N3367, N3368, N3369, 
      N3370, N3371, N3372, N3373, N3374, N3375, N3376, N3377, N3378, N3379, 
      N3380, N3381, N3382, N3383, N3384, N3385, N3386, N3387, N3388, N3389, 
      N3390, N3391, N3392, n4, n5, n10, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n5900, n6000, n6100, 
      n6300, n6400, n65, n70, n72, n73, n74, n76, n77, n78, n79, n81, n84, n85,
      n86, n87, n88, n89, n91, n92, n95, n96, n100, n101, n104, n110, n111, 
      n114, n115, n118, n119, n120, n154, n155, n156, n157, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n201, n202, n203, n204, n205, n206, n207, n208, 
      n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, 
      n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, 
      n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, 
      n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, 
      n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, 
      n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, 
      n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
      n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, 
      n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, 
      n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, 
      n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, 
      n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, 
      n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, 
      n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, 
      n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, 
      n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, 
      n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, 
      n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, 
      n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, 
      n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, 
      n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, 
      n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, 
      n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, 
      n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, 
      n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, 
      n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, 
      n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
      n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, 
      n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, 
      n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, 
      n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
      n581, n582, n583, n584, n585, n586, n587, n588, n589, n5901, n591, n592, 
      n593, n594, n595, n596, n597, n598, n599, n6001, n601, n602, n603, n604, 
      n605, n606, n607, n608, n609, n6101, n611, n612, n613, n614, n615, n616, 
      n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, 
      n629, n6301, n631, n632, n633, n634, n635, n636, n637, n638, n639, n6401,
      n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, 
      n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, 
      n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, 
      n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, 
      n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, 
      n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, 
      n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, 
      n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, 
      n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, 
      n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, 
      n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, 
      n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, 
      n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, 
      n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, 
      n809, n810, n811, n812, n813, n_1160, n_1161, n_1162, n_1163, n_1164, 
      n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, 
      n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, 
      n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, 
      n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, 
      n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, 
      n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, 
      n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, 
      n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, 
      n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, 
      n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, 
      n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, 
      n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, 
      n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, 
      n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, 
      n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, 
      n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, 
      n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, 
      n_1318, n_1319, mult_21_C241_n1549, mult_21_C241_n1548, 
      mult_21_C241_n1547, mult_21_C241_n1546, mult_21_C241_n1545, 
      mult_21_C241_n1544, mult_21_C241_n1543, mult_21_C241_n1542, 
      mult_21_C241_n1541, mult_21_C241_n1540, mult_21_C241_n1539, 
      mult_21_C241_n1538, mult_21_C241_n1537, mult_21_C241_n1536, 
      mult_21_C241_n1535, mult_21_C241_n1534, mult_21_C241_n1533, 
      mult_21_C241_n1532, mult_21_C241_n1531, mult_21_C241_n1530, 
      mult_21_C241_n1529, mult_21_C241_n1528, mult_21_C241_n1527, 
      mult_21_C241_n1526, mult_21_C241_n1525, mult_21_C241_n1524, 
      mult_21_C241_n1523, mult_21_C241_n1522, mult_21_C241_n1521, 
      mult_21_C241_n1519, mult_21_C241_n1518, mult_21_C241_n1517, 
      mult_21_C241_n1368, mult_21_C241_n1367, mult_21_C241_n1366, 
      mult_21_C241_n1365, mult_21_C241_n1364, mult_21_C241_n1363, 
      mult_21_C241_n1362, mult_21_C241_n1361, mult_21_C241_n1360, 
      mult_21_C241_n1359, mult_21_C241_n1358, mult_21_C241_n1357, 
      mult_21_C241_n1356, mult_21_C241_n1355, mult_21_C241_n1354, 
      mult_21_C241_n1353, mult_21_C241_n1352, mult_21_C241_n1351, 
      mult_21_C241_n1350, mult_21_C241_n1349, mult_21_C241_n1348, 
      mult_21_C241_n1347, mult_21_C241_n1346, mult_21_C241_n1345, 
      mult_21_C241_n1344, mult_21_C241_n1343, mult_21_C241_n1342, 
      mult_21_C241_n1341, mult_21_C241_n1340, mult_21_C241_n1339, 
      mult_21_C241_n1338, mult_21_C241_n1337, mult_21_C241_n1336, 
      mult_21_C241_n1335, mult_21_C241_n1334, mult_21_C241_n1333, 
      mult_21_C241_n1332, mult_21_C241_n1331, mult_21_C241_n1330, 
      mult_21_C241_n1329, mult_21_C241_n1328, mult_21_C241_n1327, 
      mult_21_C241_n1326, mult_21_C241_n1325, mult_21_C241_n1324, 
      mult_21_C241_n1323, mult_21_C241_n1322, mult_21_C241_n1321, 
      mult_21_C241_n1320, mult_21_C241_n1319, mult_21_C241_n1318, 
      mult_21_C241_n1317, mult_21_C241_n1316, mult_21_C241_n1315, 
      mult_21_C241_n1314, mult_21_C241_n1313, mult_21_C241_n1312, 
      mult_21_C241_n1311, mult_21_C241_n1310, mult_21_C241_n1309, 
      mult_21_C241_n1308, mult_21_C241_n1307, mult_21_C241_n1306, 
      mult_21_C241_n1305, mult_21_C241_n1304, mult_21_C241_n1303, 
      mult_21_C241_n1302, mult_21_C241_n1301, mult_21_C241_n1300, 
      mult_21_C241_n1299, mult_21_C241_n1298, mult_21_C241_n1297, 
      mult_21_C241_n1296, mult_21_C241_n1295, mult_21_C241_n1294, 
      mult_21_C241_n1293, mult_21_C241_n1292, mult_21_C241_n1291, 
      mult_21_C241_n1290, mult_21_C241_n1289, mult_21_C241_n1288, 
      mult_21_C241_n1287, mult_21_C241_n1286, mult_21_C241_n1285, 
      mult_21_C241_n1284, mult_21_C241_n1283, mult_21_C241_n1282, 
      mult_21_C241_n1281, mult_21_C241_n1280, mult_21_C241_n1279, 
      mult_21_C241_n1278, mult_21_C241_n1277, mult_21_C241_n1276, 
      mult_21_C241_n1275, mult_21_C241_n1274, mult_21_C241_n1273, 
      mult_21_C241_n1272, mult_21_C241_n1271, mult_21_C241_n1270, 
      mult_21_C241_n1269, mult_21_C241_n1268, mult_21_C241_n1267, 
      mult_21_C241_n1266, mult_21_C241_n1265, mult_21_C241_n1264, 
      mult_21_C241_n1263, mult_21_C241_n1262, mult_21_C241_n1261, 
      mult_21_C241_n1260, mult_21_C241_n1259, mult_21_C241_n1258, 
      mult_21_C241_n1257, mult_21_C241_n1256, mult_21_C241_n1255, 
      mult_21_C241_n1254, mult_21_C241_n1253, mult_21_C241_n1252, 
      mult_21_C241_n1251, mult_21_C241_n1250, mult_21_C241_n1249, 
      mult_21_C241_n1248, mult_21_C241_n1247, mult_21_C241_n1246, 
      mult_21_C241_n1245, mult_21_C241_n1244, mult_21_C241_n1243, 
      mult_21_C241_n1242, mult_21_C241_n1241, mult_21_C241_n1240, 
      mult_21_C241_n1239, mult_21_C241_n1238, mult_21_C241_n1237, 
      mult_21_C241_n1236, mult_21_C241_n1235, mult_21_C241_n1234, 
      mult_21_C241_n1233, mult_21_C241_n1232, mult_21_C241_n1231, 
      mult_21_C241_n1230, mult_21_C241_n1229, mult_21_C241_n1228, 
      mult_21_C241_n1227, mult_21_C241_n1226, mult_21_C241_n1225, 
      mult_21_C241_n1224, mult_21_C241_n1223, mult_21_C241_n1222, 
      mult_21_C241_n1221, mult_21_C241_n1220, mult_21_C241_n1219, 
      mult_21_C241_n1218, mult_21_C241_n1217, mult_21_C241_n1216, 
      mult_21_C241_n1215, mult_21_C241_n1214, mult_21_C241_n1213, 
      mult_21_C241_n1212, mult_21_C241_n1211, mult_21_C241_n1210, 
      mult_21_C241_n1209, mult_21_C241_n1208, mult_21_C241_n1207, 
      mult_21_C241_n1206, mult_21_C241_n1205, mult_21_C241_n1204, 
      mult_21_C241_n1203, mult_21_C241_n1202, mult_21_C241_n1201, 
      mult_21_C241_n1200, mult_21_C241_n1199, mult_21_C241_n1198, 
      mult_21_C241_n1197, mult_21_C241_n1196, mult_21_C241_n1195, 
      mult_21_C241_n1194, mult_21_C241_n1193, mult_21_C241_n1192, 
      mult_21_C241_n1191, mult_21_C241_n1190, mult_21_C241_n1189, 
      mult_21_C241_n1188, mult_21_C241_n1187, mult_21_C241_n1186, 
      mult_21_C241_n1185, mult_21_C241_n1184, mult_21_C241_n1183, 
      mult_21_C241_n1182, mult_21_C241_n1181, mult_21_C241_n1180, 
      mult_21_C241_n1179, mult_21_C241_n1178, mult_21_C241_n1177, 
      mult_21_C241_n1176, mult_21_C241_n1175, mult_21_C241_n1174, 
      mult_21_C241_n1173, mult_21_C241_n1172, mult_21_C241_n1171, 
      mult_21_C241_n1170, mult_21_C241_n1169, mult_21_C241_n1168, 
      mult_21_C241_n1167, mult_21_C241_n1166, mult_21_C241_n1165, 
      mult_21_C241_n1164, mult_21_C241_n1163, mult_21_C241_n1162, 
      mult_21_C241_n1161, mult_21_C241_n1160, mult_21_C241_n1159, 
      mult_21_C241_n1158, mult_21_C241_n1157, mult_21_C241_n1156, 
      mult_21_C241_n1155, mult_21_C241_n1154, mult_21_C241_n1153, 
      mult_21_C241_n1152, mult_21_C241_n1151, mult_21_C241_n1150, 
      mult_21_C241_n1149, mult_21_C241_n1148, mult_21_C241_n1147, 
      mult_21_C241_n1146, mult_21_C241_n1145, mult_21_C241_n1144, 
      mult_21_C241_n1143, mult_21_C241_n1142, mult_21_C241_n1141, 
      mult_21_C241_n1140, mult_21_C241_n1139, mult_21_C241_n1138, 
      mult_21_C241_n1137, mult_21_C241_n1136, mult_21_C241_n1135, 
      mult_21_C241_n1134, mult_21_C241_n1133, mult_21_C241_n1132, 
      mult_21_C241_n1131, mult_21_C241_n1130, mult_21_C241_n1129, 
      mult_21_C241_n1128, mult_21_C241_n1127, mult_21_C241_n1126, 
      mult_21_C241_n1125, mult_21_C241_n1124, mult_21_C241_n1123, 
      mult_21_C241_n1122, mult_21_C241_n1121, mult_21_C241_n1120, 
      mult_21_C241_n1119, mult_21_C241_n1118, mult_21_C241_n1117, 
      mult_21_C241_n1116, mult_21_C241_n1115, mult_21_C241_n1114, 
      mult_21_C241_n1113, mult_21_C241_n1112, mult_21_C241_n1111, 
      mult_21_C241_n1110, mult_21_C241_n1109, mult_21_C241_n1108, 
      mult_21_C241_n1107, mult_21_C241_n1106, mult_21_C241_n1105, 
      mult_21_C241_n1104, mult_21_C241_n1103, mult_21_C241_n1102, 
      mult_21_C241_n1101, mult_21_C241_n1100, mult_21_C241_n1099, 
      mult_21_C241_n1098, mult_21_C241_n1097, mult_21_C241_n1096, 
      mult_21_C241_n1095, mult_21_C241_n1094, mult_21_C241_n1093, 
      mult_21_C241_n1092, mult_21_C241_n1091, mult_21_C241_n1090, 
      mult_21_C241_n1089, mult_21_C241_n1088, mult_21_C241_n1087, 
      mult_21_C241_n1086, mult_21_C241_n1085, mult_21_C241_n1084, 
      mult_21_C241_n1083, mult_21_C241_n1082, mult_21_C241_n1081, 
      mult_21_C241_n1080, mult_21_C241_n1079, mult_21_C241_n1078, 
      mult_21_C241_n1077, mult_21_C241_n1076, mult_21_C241_n1075, 
      mult_21_C241_n1074, mult_21_C241_n1073, mult_21_C241_n1072, 
      mult_21_C241_n1071, mult_21_C241_n1070, mult_21_C241_n1069, 
      mult_21_C241_n1068, mult_21_C241_n1067, mult_21_C241_n1066, 
      mult_21_C241_n1065, mult_21_C241_n1064, mult_21_C241_n1063, 
      mult_21_C241_n1062, mult_21_C241_n1061, mult_21_C241_n1060, 
      mult_21_C241_n1059, mult_21_C241_n1058, mult_21_C241_n1057, 
      mult_21_C241_n1056, mult_21_C241_n1055, mult_21_C241_n1054, 
      mult_21_C241_n1053, mult_21_C241_n1052, mult_21_C241_n1051, 
      mult_21_C241_n1050, mult_21_C241_n1049, mult_21_C241_n1048, 
      mult_21_C241_n1047, mult_21_C241_n1046, mult_21_C241_n1045, 
      mult_21_C241_n1044, mult_21_C241_n1043, mult_21_C241_n1042, 
      mult_21_C241_n1041, mult_21_C241_n1040, mult_21_C241_n1039, 
      mult_21_C241_n1038, mult_21_C241_n1037, mult_21_C241_n1036, 
      mult_21_C241_n1035, mult_21_C241_n1034, mult_21_C241_n1033, 
      mult_21_C241_n1032, mult_21_C241_n1031, mult_21_C241_n1030, 
      mult_21_C241_n1029, mult_21_C241_n1028, mult_21_C241_n1027, 
      mult_21_C241_n1026, mult_21_C241_n1025, mult_21_C241_n1024, 
      mult_21_C241_n1023, mult_21_C241_n1022, mult_21_C241_n1021, 
      mult_21_C241_n1020, mult_21_C241_n1019, mult_21_C241_n1018, 
      mult_21_C241_n1017, mult_21_C241_n1016, mult_21_C241_n1015, 
      mult_21_C241_n1014, mult_21_C241_n1013, mult_21_C241_n1012, 
      mult_21_C241_n1011, mult_21_C241_n1010, mult_21_C241_n1009, 
      mult_21_C241_n1008, mult_21_C241_n1007, mult_21_C241_n1006, 
      mult_21_C241_n1005, mult_21_C241_n1004, mult_21_C241_n1003, 
      mult_21_C241_n1002, mult_21_C241_n1001, mult_21_C241_n1000, 
      mult_21_C241_n999, mult_21_C241_n998, mult_21_C241_n997, 
      mult_21_C241_n996, mult_21_C241_n995, mult_21_C241_n994, 
      mult_21_C241_n993, mult_21_C241_n992, mult_21_C241_n991, 
      mult_21_C241_n990, mult_21_C241_n989, mult_21_C241_n988, 
      mult_21_C241_n987, mult_21_C241_n986, mult_21_C241_n985, 
      mult_21_C241_n984, mult_21_C241_n983, mult_21_C241_n982, 
      mult_21_C241_n981, mult_21_C241_n980, mult_21_C241_n979, 
      mult_21_C241_n978, mult_21_C241_n977, mult_21_C241_n976, 
      mult_21_C241_n975, mult_21_C241_n974, mult_21_C241_n973, 
      mult_21_C241_n972, mult_21_C241_n971, mult_21_C241_n970, 
      mult_21_C241_n969, mult_21_C241_n968, mult_21_C241_n967, 
      mult_21_C241_n966, mult_21_C241_n965, mult_21_C241_n964, 
      mult_21_C241_n963, mult_21_C241_n962, mult_21_C241_n961, 
      mult_21_C241_n960, mult_21_C241_n959, mult_21_C241_n958, 
      mult_21_C241_n957, mult_21_C241_n956, mult_21_C241_n955, 
      mult_21_C241_n954, mult_21_C241_n953, mult_21_C241_n952, 
      mult_21_C241_n951, mult_21_C241_n950, mult_21_C241_n949, 
      mult_21_C241_n948, mult_21_C241_n947, mult_21_C241_n946, 
      mult_21_C241_n945, mult_21_C241_n944, mult_21_C241_n943, 
      mult_21_C241_n942, mult_21_C241_n941, mult_21_C241_n940, 
      mult_21_C241_n939, mult_21_C241_n938, mult_21_C241_n937, 
      mult_21_C241_n936, mult_21_C241_n935, mult_21_C241_n934, 
      mult_21_C241_n933, mult_21_C241_n932, mult_21_C241_n931, 
      mult_21_C241_n930, mult_21_C241_n929, mult_21_C241_n928, 
      mult_21_C241_n927, mult_21_C241_n926, mult_21_C241_n925, 
      mult_21_C241_n924, mult_21_C241_n923, mult_21_C241_n922, 
      mult_21_C241_n921, mult_21_C241_n920, mult_21_C241_n919, 
      mult_21_C241_n918, mult_21_C241_n917, mult_21_C241_n916, 
      mult_21_C241_n915, mult_21_C241_n914, mult_21_C241_n913, 
      mult_21_C241_n912, mult_21_C241_n911, mult_21_C241_n910, 
      mult_21_C241_n909, mult_21_C241_n908, mult_21_C241_n907, 
      mult_21_C241_n906, mult_21_C241_n905, mult_21_C241_n904, 
      mult_21_C241_n903, mult_21_C241_n902, mult_21_C241_n901, 
      mult_21_C241_n900, mult_21_C241_n899, mult_21_C241_n898, 
      mult_21_C241_n897, mult_21_C241_n896, mult_21_C241_n895, 
      mult_21_C241_n894, mult_21_C241_n893, mult_21_C241_n892, 
      mult_21_C241_n891, mult_21_C241_n890, mult_21_C241_n889, 
      mult_21_C241_n888, mult_21_C241_n887, mult_21_C241_n886, 
      mult_21_C241_n885, mult_21_C241_n884, mult_21_C241_n883, 
      mult_21_C241_n882, mult_21_C241_n881, mult_21_C241_n880, 
      mult_21_C241_n879, mult_21_C241_n878, mult_21_C241_n877, 
      mult_21_C241_n876, mult_21_C241_n875, mult_21_C241_n874, 
      mult_21_C241_n873, mult_21_C241_n872, mult_21_C241_n871, 
      mult_21_C241_n870, mult_21_C241_n869, mult_21_C241_n868, 
      mult_21_C241_n867, mult_21_C241_n866, mult_21_C241_n865, 
      mult_21_C241_n864, mult_21_C241_n863, mult_21_C241_n862, 
      mult_21_C241_n861, mult_21_C241_n860, mult_21_C241_n859, 
      mult_21_C241_n858, mult_21_C241_n857, mult_21_C241_n856, 
      mult_21_C241_n855, mult_21_C241_n854, mult_21_C241_n853, 
      mult_21_C241_n852, mult_21_C241_n851, mult_21_C241_n850, 
      mult_21_C241_n849, mult_21_C241_n848, mult_21_C241_n847, 
      mult_21_C241_n846, mult_21_C241_n845, mult_21_C241_n844, 
      mult_21_C241_n843, mult_21_C241_n842, mult_21_C241_n841, 
      mult_21_C241_n840, mult_21_C241_n839, mult_21_C241_n838, 
      mult_21_C241_n837, mult_21_C241_n836, mult_21_C241_n835, 
      mult_21_C241_n834, mult_21_C241_n833, mult_21_C241_n832, 
      mult_21_C241_n831, mult_21_C241_n830, mult_21_C241_n829, 
      mult_21_C241_n828, mult_21_C241_n827, mult_21_C241_n826, 
      mult_21_C241_n825, mult_21_C241_n824, mult_21_C241_n823, 
      mult_21_C241_n822, mult_21_C241_n821, mult_21_C241_n820, 
      mult_21_C241_n819, mult_21_C241_n818, mult_21_C241_n817, 
      mult_21_C241_n816, mult_21_C241_n815, mult_21_C241_n814, 
      mult_21_C241_n813, mult_21_C241_n812, mult_21_C241_n811, 
      mult_21_C241_n810, mult_21_C241_n809, mult_21_C241_n808, 
      mult_21_C241_n807, mult_21_C241_n806, mult_21_C241_n805, 
      mult_21_C241_n804, mult_21_C241_n803, mult_21_C241_n802, 
      mult_21_C241_n801, mult_21_C241_n800, mult_21_C241_n799, 
      mult_21_C241_n798, mult_21_C241_n797, mult_21_C241_n796, 
      mult_21_C241_n795, mult_21_C241_n794, mult_21_C241_n793, 
      mult_21_C241_n792, mult_21_C241_n791, mult_21_C241_n790, 
      mult_21_C241_n789, mult_21_C241_n788, mult_21_C241_n787, 
      mult_21_C241_n786, mult_21_C241_n785, mult_21_C241_n784, 
      mult_21_C241_n783, mult_21_C241_n782, mult_21_C241_n781, 
      mult_21_C241_n780, mult_21_C241_n779, mult_21_C241_n778, 
      mult_21_C241_n777, mult_21_C241_n776, mult_21_C241_n775, 
      mult_21_C241_n774, mult_21_C241_n773, mult_21_C241_n772, 
      mult_21_C241_n771, mult_21_C241_n770, mult_21_C241_n769, 
      mult_21_C241_n768, mult_21_C241_n767, mult_21_C241_n766, 
      mult_21_C241_n765, mult_21_C241_n764, mult_21_C241_n763, 
      mult_21_C241_n762, mult_21_C241_n761, mult_21_C241_n760, 
      mult_21_C241_n759, mult_21_C241_n758, mult_21_C241_n757, 
      mult_21_C241_n756, mult_21_C241_n755, mult_21_C241_n754, 
      mult_21_C241_n753, mult_21_C241_n752, mult_21_C241_n751, 
      mult_21_C241_n750, mult_21_C241_n749, mult_21_C241_n748, 
      mult_21_C241_n747, mult_21_C241_n746, mult_21_C241_n745, 
      mult_21_C241_n744, mult_21_C241_n743, mult_21_C241_n742, 
      mult_21_C241_n741, mult_21_C241_n740, mult_21_C241_n739, 
      mult_21_C241_n738, mult_21_C241_n737, mult_21_C241_n736, 
      mult_21_C241_n735, mult_21_C241_n734, mult_21_C241_n733, 
      mult_21_C241_n732, mult_21_C241_n731, mult_21_C241_n730, 
      mult_21_C241_n729, mult_21_C241_n728, mult_21_C241_n727, 
      mult_21_C241_n726, mult_21_C241_n725, mult_21_C241_n724, 
      mult_21_C241_n723, mult_21_C241_n722, mult_21_C241_n721, 
      mult_21_C241_n720, mult_21_C241_n719, mult_21_C241_n718, 
      mult_21_C241_n717, mult_21_C241_n716, mult_21_C241_n715, 
      mult_21_C241_n714, mult_21_C241_n713, mult_21_C241_n712, 
      mult_21_C241_n711, mult_21_C241_n710, mult_21_C241_n709, 
      mult_21_C241_n708, mult_21_C241_n707, mult_21_C241_n706, 
      mult_21_C241_n705, mult_21_C241_n704, mult_21_C241_n703, 
      mult_21_C241_n702, mult_21_C241_n701, mult_21_C241_n700, 
      mult_21_C241_n699, mult_21_C241_n698, mult_21_C241_n697, 
      mult_21_C241_n696, mult_21_C241_n695, mult_21_C241_n694, 
      mult_21_C241_n693, mult_21_C241_n692, mult_21_C241_n691, 
      mult_21_C241_n690, mult_21_C241_n689, mult_21_C241_n688, 
      mult_21_C241_n687, mult_21_C241_n686, mult_21_C241_n685, 
      mult_21_C241_n684, mult_21_C241_n683, mult_21_C241_n682, 
      mult_21_C241_n681, mult_21_C241_n680, mult_21_C241_n679, 
      mult_21_C241_n678, mult_21_C241_n677, mult_21_C241_n676, 
      mult_21_C241_n675, mult_21_C241_n674, mult_21_C241_n673, 
      mult_21_C241_n672, mult_21_C241_n671, mult_21_C241_n670, 
      mult_21_C241_n669, mult_21_C241_n668, mult_21_C241_n667, 
      mult_21_C241_n666, mult_21_C241_n665, mult_21_C241_n664, 
      mult_21_C241_n663, mult_21_C241_n662, mult_21_C241_n661, 
      mult_21_C241_n660, mult_21_C241_n659, mult_21_C241_n658, 
      mult_21_C241_n657, mult_21_C241_n656, mult_21_C241_n655, 
      mult_21_C241_n654, mult_21_C241_n653, mult_21_C241_n652, 
      mult_21_C241_n651, mult_21_C241_n650, mult_21_C241_n649, 
      mult_21_C241_n648, mult_21_C241_n647, mult_21_C241_n646, 
      mult_21_C241_n645, mult_21_C241_n644, mult_21_C241_n643, 
      mult_21_C241_n642, mult_21_C241_n641, mult_21_C241_n640, 
      mult_21_C241_n639, mult_21_C241_n638, mult_21_C241_n637, 
      mult_21_C241_n636, mult_21_C241_n635, mult_21_C241_n634, 
      mult_21_C241_n633, mult_21_C241_n632, mult_21_C241_n631, 
      mult_21_C241_n630, mult_21_C241_n629, mult_21_C241_n628, 
      mult_21_C241_n627, mult_21_C241_n626, mult_21_C241_n625, 
      mult_21_C241_n624, mult_21_C241_n623, mult_21_C241_n622, 
      mult_21_C241_n621, mult_21_C241_n620, mult_21_C241_n619, 
      mult_21_C241_n618, mult_21_C241_n617, mult_21_C241_n616, 
      mult_21_C241_n615, mult_21_C241_n614, mult_21_C241_n613, 
      mult_21_C241_n612, mult_21_C241_n611, mult_21_C241_n610, 
      mult_21_C241_n609, mult_21_C241_n608, mult_21_C241_n607, 
      mult_21_C241_n606, mult_21_C241_n605, mult_21_C241_n604, 
      mult_21_C241_n603, mult_21_C241_n602, mult_21_C241_n601, 
      mult_21_C241_n600, mult_21_C241_n599, mult_21_C241_n598, 
      mult_21_C241_n597, mult_21_C241_n596, mult_21_C241_n595, 
      mult_21_C241_n594, mult_21_C241_n593, mult_21_C241_n592, 
      mult_21_C241_n591, mult_21_C241_n590, mult_21_C241_n589, 
      mult_21_C241_n588, mult_21_C241_n587, mult_21_C241_n586, 
      mult_21_C241_n585, mult_21_C241_n584, mult_21_C241_n583, 
      mult_21_C241_n582, mult_21_C241_n581, mult_21_C241_n580, 
      mult_21_C241_n579, mult_21_C241_n578, mult_21_C241_n577, 
      mult_21_C241_n576, mult_21_C241_n575, mult_21_C241_n574, 
      mult_21_C241_n573, mult_21_C241_n572, mult_21_C241_n571, 
      mult_21_C241_n570, mult_21_C241_n569, mult_21_C241_n568, 
      mult_21_C241_n567, mult_21_C241_n566, mult_21_C241_n565, 
      mult_21_C241_n564, mult_21_C241_n563, mult_21_C241_n562, 
      mult_21_C241_n561, mult_21_C241_n560, mult_21_C241_n559, 
      mult_21_C241_n558, mult_21_C241_n557, mult_21_C241_n556, 
      mult_21_C241_n555, mult_21_C241_n554, mult_21_C241_n553, 
      mult_21_C241_n552, mult_21_C241_n551, mult_21_C241_n550, 
      mult_21_C241_n549, mult_21_C241_n548, mult_21_C241_n547, 
      mult_21_C241_n546, mult_21_C241_n545, mult_21_C241_n544, 
      mult_21_C241_n543, mult_21_C241_n542, mult_21_C241_n541, 
      mult_21_C241_n540, mult_21_C241_n539, mult_21_C241_n538, 
      mult_21_C241_n537, mult_21_C241_n536, mult_21_C241_n535, 
      mult_21_C241_n534, mult_21_C241_n533, mult_21_C241_n532, 
      mult_21_C241_n531, mult_21_C241_n530, mult_21_C241_n529, 
      mult_21_C241_n528, mult_21_C241_n527, mult_21_C241_n526, 
      mult_21_C241_n525, mult_21_C241_n524, mult_21_C241_n523, 
      mult_21_C241_n522, mult_21_C241_n521, mult_21_C241_n520, 
      mult_21_C241_n519, mult_21_C241_n518, mult_21_C241_n517, 
      mult_21_C241_n516, mult_21_C241_n515, mult_21_C241_n514, 
      mult_21_C241_n513, mult_21_C241_n512, mult_21_C241_n511, 
      mult_21_C241_n510, mult_21_C241_n509, mult_21_C241_n508, 
      mult_21_C241_n507, mult_21_C241_n506, mult_21_C241_n505, 
      mult_21_C241_n504, mult_21_C241_n503, mult_21_C241_n502, 
      mult_21_C241_n501, mult_21_C241_n500, mult_21_C241_n499, 
      mult_21_C241_n498, mult_21_C241_n497, mult_21_C241_n496, 
      mult_21_C241_n495, mult_21_C241_n494, mult_21_C241_n493, 
      mult_21_C241_n492, mult_21_C241_n491, mult_21_C241_n490, 
      mult_21_C241_n489, mult_21_C241_n488, mult_21_C241_n487, 
      mult_21_C241_n486, mult_21_C241_n485, mult_21_C241_n484, 
      mult_21_C241_n483, mult_21_C241_n482, mult_21_C241_n481, 
      mult_21_C241_n480, mult_21_C241_n479, mult_21_C241_n478, 
      mult_21_C241_n477, mult_21_C241_n476, mult_21_C241_n475, 
      mult_21_C241_n474, mult_21_C241_n473, mult_21_C241_n472, 
      mult_21_C241_n471, mult_21_C241_n470, mult_21_C241_n469, 
      mult_21_C241_n468, mult_21_C241_n467, mult_21_C241_n466, 
      mult_21_C241_n465, mult_21_C241_n464, mult_21_C241_n463, 
      mult_21_C241_n462, mult_21_C241_n461, mult_21_C241_n460, 
      mult_21_C241_n459, mult_21_C241_n458, mult_21_C241_n457, 
      mult_21_C241_n456, mult_21_C241_n455, mult_21_C241_n454, 
      mult_21_C241_n453, mult_21_C241_n452, mult_21_C241_n451, 
      mult_21_C241_n450, mult_21_C241_n449, mult_21_C241_n448, 
      mult_21_C241_n447, mult_21_C241_n446, mult_21_C241_n445, 
      mult_21_C241_n444, mult_21_C241_n443, mult_21_C241_n442, 
      mult_21_C241_n441, mult_21_C241_n440, mult_21_C241_n439, 
      mult_21_C241_n438, mult_21_C241_n437, mult_21_C241_n436, 
      mult_21_C241_n435, mult_21_C241_n434, mult_21_C241_n433, 
      mult_21_C241_n432, mult_21_C241_n431, mult_21_C241_n430, 
      mult_21_C241_n429, mult_21_C241_n428, mult_21_C241_n427, 
      mult_21_C241_n426, mult_21_C241_n425, mult_21_C241_n424, 
      mult_21_C241_n423, mult_21_C241_n422, mult_21_C241_n421, 
      mult_21_C241_n420, mult_21_C241_n419, mult_21_C241_n418, 
      mult_21_C241_n417, mult_21_C241_n416, mult_21_C241_n415, 
      mult_21_C241_n414, mult_21_C241_n413, mult_21_C241_n412, 
      mult_21_C241_n411, mult_21_C241_n410, mult_21_C241_n409, 
      mult_21_C241_n408, mult_21_C241_n407, mult_21_C241_n406, 
      mult_21_C241_n405, mult_21_C241_n404, mult_21_C241_n403, 
      mult_21_C241_n402, mult_21_C241_n401, mult_21_C241_n400, 
      mult_21_C241_n399, mult_21_C241_n398, mult_21_C241_n397, 
      mult_21_C241_n396, mult_21_C241_n395, mult_21_C241_n394, 
      mult_21_C241_n393, mult_21_C241_n392, mult_21_C241_n391, 
      mult_21_C241_n390, mult_21_C241_n389, mult_21_C241_n388, 
      mult_21_C241_n387, mult_21_C241_n386, mult_21_C241_n385, 
      mult_21_C241_n384, mult_21_C241_n383, mult_21_C241_n382, 
      mult_21_C241_n381, mult_21_C241_n380, mult_21_C241_n379, 
      mult_21_C241_n378, mult_21_C241_n377, mult_21_C241_n376, 
      mult_21_C241_n375, mult_21_C241_n374, mult_21_C241_n373, 
      mult_21_C241_n372, mult_21_C241_n371, mult_21_C241_n370, 
      mult_21_C241_n369, mult_21_C241_n368, mult_21_C241_n367, 
      mult_21_C241_n366, mult_21_C241_n365, mult_21_C241_n364, 
      mult_21_C241_n363, mult_21_C241_n362, mult_21_C241_n361, 
      mult_21_C241_n360, mult_21_C241_n359, mult_21_C241_n358, 
      mult_21_C241_n357, mult_21_C241_n356, mult_21_C241_n355, 
      mult_21_C241_n354, mult_21_C241_n353, mult_21_C241_n352, 
      mult_21_C241_n351, mult_21_C241_n350, mult_21_C241_n349, 
      mult_21_C241_n348, mult_21_C241_n347, mult_21_C241_n346, 
      mult_21_C241_n345, mult_21_C241_n344, mult_21_C241_n343, 
      mult_21_C241_n342, mult_21_C241_n341, mult_21_C241_n340, 
      mult_21_C241_n339, mult_21_C241_n338, mult_21_C241_n337, 
      mult_21_C241_n336, mult_21_C241_n335, mult_21_C241_n334, 
      mult_21_C241_n333, mult_21_C241_n332, mult_21_C241_n331, 
      mult_21_C241_n330, mult_21_C241_n329, mult_21_C241_n326, 
      mult_21_C241_n324, mult_21_C241_n323, mult_21_C241_n322, 
      mult_21_C241_n319, mult_21_C241_n318, mult_21_C241_n315, 
      mult_21_C241_n314, mult_21_C241_n313, mult_21_C241_n312, 
      mult_21_C241_n310, mult_21_C241_n305, mult_21_C241_n303, 
      mult_21_C241_n302, mult_21_C241_n301, mult_21_C241_n297, 
      mult_21_C241_n296, mult_21_C241_n295, mult_21_C241_n294, 
      mult_21_C241_n293, mult_21_C241_n289, mult_21_C241_n288, 
      mult_21_C241_n287, mult_21_C241_n286, mult_21_C241_n285, 
      mult_21_C241_n284, mult_21_C241_n283, mult_21_C241_n282, 
      mult_21_C241_n281, mult_21_C241_n280, mult_21_C241_n279, 
      mult_21_C241_n278, mult_21_C241_n277, mult_21_C241_n276, 
      mult_21_C241_n275, mult_21_C241_n273, mult_21_C241_n271, 
      mult_21_C241_n270, mult_21_C241_n268, mult_21_C241_n266, 
      mult_21_C241_n265, mult_21_C241_n264, mult_21_C241_n263, 
      mult_21_C241_n262, mult_21_C241_n261, mult_21_C241_n260, 
      mult_21_C241_n259, mult_21_C241_n258, mult_21_C241_n257, 
      mult_21_C241_n256, mult_21_C241_n255, mult_21_C241_n254, 
      mult_21_C241_n253, mult_21_C241_n251, mult_21_C241_n249, 
      mult_21_C241_n248, mult_21_C241_n246, mult_21_C241_n244, 
      mult_21_C241_n243, mult_21_C241_n242, mult_21_C241_n241, 
      mult_21_C241_n240, mult_21_C241_n239, mult_21_C241_n238, 
      mult_21_C241_n237, mult_21_C241_n236, mult_21_C241_n235, 
      mult_21_C241_n234, mult_21_C241_n233, mult_21_C241_n232, 
      mult_21_C241_n231, mult_21_C241_n230, mult_21_C241_n229, 
      mult_21_C241_n227, mult_21_C241_n226, mult_21_C241_n225, 
      mult_21_C241_n224, mult_21_C241_n223, mult_21_C241_n222, 
      mult_21_C241_n221, mult_21_C241_n219, mult_21_C241_n217, 
      mult_21_C241_n216, mult_21_C241_n215, mult_21_C241_n214, 
      mult_21_C241_n211, mult_21_C241_n209, mult_21_C241_n208, 
      mult_21_C241_n207, mult_21_C241_n206, mult_21_C241_n204, 
      mult_21_C241_n202, mult_21_C241_n201, mult_21_C241_n200, 
      mult_21_C241_n199, mult_21_C241_n197, mult_21_C241_n195, 
      mult_21_C241_n194, mult_21_C241_n190, mult_21_C241_n189, 
      mult_21_C241_n188, mult_21_C241_n187, mult_21_C241_n185, 
      mult_21_C241_n184, mult_21_C241_n183, mult_21_C241_n182, 
      mult_21_C241_n181, mult_21_C241_n180, mult_21_C241_n179, 
      mult_21_C241_n178, mult_21_C241_n176, mult_21_C241_n175, 
      mult_21_C241_n174, mult_21_C241_n173, mult_21_C241_n172, 
      mult_21_C241_n171, mult_21_C241_n170, mult_21_C241_n169, 
      mult_21_C241_n168, mult_21_C241_n167, mult_21_C241_n166, 
      mult_21_C241_n165, mult_21_C241_n164, mult_21_C241_n163, 
      mult_21_C241_n162, mult_21_C241_n161, mult_21_C241_n160, 
      mult_21_C241_n159, mult_21_C241_n158, mult_21_C241_n157, 
      mult_21_C241_n156, mult_21_C241_n155, mult_21_C241_n106, 
      mult_21_C241_n105, mult_21_C241_n104, mult_21_C241_n103, 
      mult_21_C241_n101, mult_21_C241_n99, mult_21_C241_n98, mult_21_C241_n96, 
      mult_21_C241_n94, mult_21_C241_n93, mult_21_C241_n91, mult_21_C241_n89, 
      mult_21_C241_n88, mult_21_C241_n86, mult_21_C241_n84, mult_21_C241_n83, 
      mult_21_C241_n81, mult_21_C241_n79, mult_21_C241_n78, mult_21_C241_n76, 
      mult_21_C241_n73, mult_21_C241_n71, mult_21_C241_n69, mult_21_C241_n66, 
      mult_21_C241_n63, mult_21_C241_n61, mult_21_C241_n58, mult_21_C241_n56, 
      mult_21_C241_n53, mult_21_C241_n50, mult_21_C241_n48, mult_21_C241_n45, 
      mult_21_C241_n42, mult_21_C241_n38, mult_21_C241_n30, mult_21_C241_n22, 
      mult_21_C241_n14, mult_21_C241_n8, mult_21_C241_n6, mult_21_C241_n3, 
      mult_21_C243_n1546, mult_21_C243_n1545, mult_21_C243_n1544, 
      mult_21_C243_n1543, mult_21_C243_n1542, mult_21_C243_n1541, 
      mult_21_C243_n1540, mult_21_C243_n1539, mult_21_C243_n1538, 
      mult_21_C243_n1537, mult_21_C243_n1536, mult_21_C243_n1535, 
      mult_21_C243_n1534, mult_21_C243_n1533, mult_21_C243_n1532, 
      mult_21_C243_n1531, mult_21_C243_n1530, mult_21_C243_n1529, 
      mult_21_C243_n1528, mult_21_C243_n1527, mult_21_C243_n1526, 
      mult_21_C243_n1525, mult_21_C243_n1524, mult_21_C243_n1523, 
      mult_21_C243_n1522, mult_21_C243_n1521, mult_21_C243_n1519, 
      mult_21_C243_n1518, mult_21_C243_n1517, mult_21_C243_n1368, 
      mult_21_C243_n1367, mult_21_C243_n1366, mult_21_C243_n1365, 
      mult_21_C243_n1364, mult_21_C243_n1363, mult_21_C243_n1362, 
      mult_21_C243_n1361, mult_21_C243_n1360, mult_21_C243_n1359, 
      mult_21_C243_n1358, mult_21_C243_n1357, mult_21_C243_n1356, 
      mult_21_C243_n1355, mult_21_C243_n1354, mult_21_C243_n1353, 
      mult_21_C243_n1352, mult_21_C243_n1351, mult_21_C243_n1350, 
      mult_21_C243_n1349, mult_21_C243_n1348, mult_21_C243_n1347, 
      mult_21_C243_n1346, mult_21_C243_n1345, mult_21_C243_n1344, 
      mult_21_C243_n1343, mult_21_C243_n1342, mult_21_C243_n1341, 
      mult_21_C243_n1340, mult_21_C243_n1339, mult_21_C243_n1338, 
      mult_21_C243_n1337, mult_21_C243_n1336, mult_21_C243_n1335, 
      mult_21_C243_n1334, mult_21_C243_n1333, mult_21_C243_n1332, 
      mult_21_C243_n1331, mult_21_C243_n1330, mult_21_C243_n1329, 
      mult_21_C243_n1328, mult_21_C243_n1327, mult_21_C243_n1326, 
      mult_21_C243_n1325, mult_21_C243_n1324, mult_21_C243_n1323, 
      mult_21_C243_n1322, mult_21_C243_n1321, mult_21_C243_n1320, 
      mult_21_C243_n1319, mult_21_C243_n1318, mult_21_C243_n1317, 
      mult_21_C243_n1316, mult_21_C243_n1315, mult_21_C243_n1314, 
      mult_21_C243_n1313, mult_21_C243_n1312, mult_21_C243_n1311, 
      mult_21_C243_n1310, mult_21_C243_n1309, mult_21_C243_n1308, 
      mult_21_C243_n1307, mult_21_C243_n1306, mult_21_C243_n1305, 
      mult_21_C243_n1304, mult_21_C243_n1303, mult_21_C243_n1302, 
      mult_21_C243_n1301, mult_21_C243_n1300, mult_21_C243_n1299, 
      mult_21_C243_n1298, mult_21_C243_n1297, mult_21_C243_n1296, 
      mult_21_C243_n1295, mult_21_C243_n1294, mult_21_C243_n1293, 
      mult_21_C243_n1292, mult_21_C243_n1291, mult_21_C243_n1290, 
      mult_21_C243_n1289, mult_21_C243_n1288, mult_21_C243_n1287, 
      mult_21_C243_n1286, mult_21_C243_n1285, mult_21_C243_n1284, 
      mult_21_C243_n1283, mult_21_C243_n1282, mult_21_C243_n1281, 
      mult_21_C243_n1280, mult_21_C243_n1279, mult_21_C243_n1278, 
      mult_21_C243_n1277, mult_21_C243_n1276, mult_21_C243_n1275, 
      mult_21_C243_n1274, mult_21_C243_n1273, mult_21_C243_n1272, 
      mult_21_C243_n1271, mult_21_C243_n1270, mult_21_C243_n1269, 
      mult_21_C243_n1268, mult_21_C243_n1267, mult_21_C243_n1266, 
      mult_21_C243_n1265, mult_21_C243_n1264, mult_21_C243_n1263, 
      mult_21_C243_n1262, mult_21_C243_n1261, mult_21_C243_n1260, 
      mult_21_C243_n1259, mult_21_C243_n1258, mult_21_C243_n1257, 
      mult_21_C243_n1256, mult_21_C243_n1255, mult_21_C243_n1254, 
      mult_21_C243_n1253, mult_21_C243_n1252, mult_21_C243_n1251, 
      mult_21_C243_n1250, mult_21_C243_n1249, mult_21_C243_n1248, 
      mult_21_C243_n1247, mult_21_C243_n1246, mult_21_C243_n1245, 
      mult_21_C243_n1244, mult_21_C243_n1243, mult_21_C243_n1242, 
      mult_21_C243_n1241, mult_21_C243_n1240, mult_21_C243_n1239, 
      mult_21_C243_n1238, mult_21_C243_n1237, mult_21_C243_n1236, 
      mult_21_C243_n1235, mult_21_C243_n1234, mult_21_C243_n1233, 
      mult_21_C243_n1232, mult_21_C243_n1231, mult_21_C243_n1230, 
      mult_21_C243_n1229, mult_21_C243_n1228, mult_21_C243_n1227, 
      mult_21_C243_n1226, mult_21_C243_n1225, mult_21_C243_n1224, 
      mult_21_C243_n1223, mult_21_C243_n1222, mult_21_C243_n1221, 
      mult_21_C243_n1220, mult_21_C243_n1219, mult_21_C243_n1218, 
      mult_21_C243_n1217, mult_21_C243_n1216, mult_21_C243_n1215, 
      mult_21_C243_n1214, mult_21_C243_n1213, mult_21_C243_n1212, 
      mult_21_C243_n1211, mult_21_C243_n1210, mult_21_C243_n1209, 
      mult_21_C243_n1208, mult_21_C243_n1207, mult_21_C243_n1206, 
      mult_21_C243_n1205, mult_21_C243_n1204, mult_21_C243_n1203, 
      mult_21_C243_n1202, mult_21_C243_n1201, mult_21_C243_n1200, 
      mult_21_C243_n1199, mult_21_C243_n1198, mult_21_C243_n1197, 
      mult_21_C243_n1196, mult_21_C243_n1195, mult_21_C243_n1194, 
      mult_21_C243_n1193, mult_21_C243_n1192, mult_21_C243_n1191, 
      mult_21_C243_n1190, mult_21_C243_n1189, mult_21_C243_n1188, 
      mult_21_C243_n1187, mult_21_C243_n1186, mult_21_C243_n1185, 
      mult_21_C243_n1184, mult_21_C243_n1183, mult_21_C243_n1182, 
      mult_21_C243_n1181, mult_21_C243_n1180, mult_21_C243_n1179, 
      mult_21_C243_n1178, mult_21_C243_n1177, mult_21_C243_n1176, 
      mult_21_C243_n1175, mult_21_C243_n1174, mult_21_C243_n1173, 
      mult_21_C243_n1172, mult_21_C243_n1171, mult_21_C243_n1170, 
      mult_21_C243_n1169, mult_21_C243_n1168, mult_21_C243_n1167, 
      mult_21_C243_n1166, mult_21_C243_n1165, mult_21_C243_n1164, 
      mult_21_C243_n1163, mult_21_C243_n1162, mult_21_C243_n1161, 
      mult_21_C243_n1160, mult_21_C243_n1159, mult_21_C243_n1158, 
      mult_21_C243_n1157, mult_21_C243_n1156, mult_21_C243_n1155, 
      mult_21_C243_n1154, mult_21_C243_n1153, mult_21_C243_n1152, 
      mult_21_C243_n1151, mult_21_C243_n1150, mult_21_C243_n1149, 
      mult_21_C243_n1148, mult_21_C243_n1147, mult_21_C243_n1146, 
      mult_21_C243_n1145, mult_21_C243_n1144, mult_21_C243_n1143, 
      mult_21_C243_n1142, mult_21_C243_n1141, mult_21_C243_n1140, 
      mult_21_C243_n1139, mult_21_C243_n1138, mult_21_C243_n1137, 
      mult_21_C243_n1136, mult_21_C243_n1135, mult_21_C243_n1134, 
      mult_21_C243_n1133, mult_21_C243_n1132, mult_21_C243_n1131, 
      mult_21_C243_n1130, mult_21_C243_n1129, mult_21_C243_n1128, 
      mult_21_C243_n1127, mult_21_C243_n1126, mult_21_C243_n1125, 
      mult_21_C243_n1124, mult_21_C243_n1123, mult_21_C243_n1122, 
      mult_21_C243_n1121, mult_21_C243_n1120, mult_21_C243_n1119, 
      mult_21_C243_n1118, mult_21_C243_n1117, mult_21_C243_n1116, 
      mult_21_C243_n1115, mult_21_C243_n1114, mult_21_C243_n1113, 
      mult_21_C243_n1112, mult_21_C243_n1111, mult_21_C243_n1110, 
      mult_21_C243_n1109, mult_21_C243_n1108, mult_21_C243_n1107, 
      mult_21_C243_n1106, mult_21_C243_n1105, mult_21_C243_n1104, 
      mult_21_C243_n1103, mult_21_C243_n1102, mult_21_C243_n1101, 
      mult_21_C243_n1100, mult_21_C243_n1099, mult_21_C243_n1098, 
      mult_21_C243_n1097, mult_21_C243_n1096, mult_21_C243_n1095, 
      mult_21_C243_n1094, mult_21_C243_n1093, mult_21_C243_n1092, 
      mult_21_C243_n1091, mult_21_C243_n1090, mult_21_C243_n1089, 
      mult_21_C243_n1088, mult_21_C243_n1087, mult_21_C243_n1086, 
      mult_21_C243_n1085, mult_21_C243_n1084, mult_21_C243_n1083, 
      mult_21_C243_n1082, mult_21_C243_n1081, mult_21_C243_n1080, 
      mult_21_C243_n1079, mult_21_C243_n1078, mult_21_C243_n1077, 
      mult_21_C243_n1076, mult_21_C243_n1075, mult_21_C243_n1074, 
      mult_21_C243_n1073, mult_21_C243_n1072, mult_21_C243_n1071, 
      mult_21_C243_n1070, mult_21_C243_n1069, mult_21_C243_n1068, 
      mult_21_C243_n1067, mult_21_C243_n1066, mult_21_C243_n1065, 
      mult_21_C243_n1064, mult_21_C243_n1063, mult_21_C243_n1062, 
      mult_21_C243_n1061, mult_21_C243_n1060, mult_21_C243_n1059, 
      mult_21_C243_n1058, mult_21_C243_n1057, mult_21_C243_n1056, 
      mult_21_C243_n1055, mult_21_C243_n1054, mult_21_C243_n1053, 
      mult_21_C243_n1052, mult_21_C243_n1051, mult_21_C243_n1050, 
      mult_21_C243_n1049, mult_21_C243_n1048, mult_21_C243_n1047, 
      mult_21_C243_n1046, mult_21_C243_n1045, mult_21_C243_n1044, 
      mult_21_C243_n1043, mult_21_C243_n1042, mult_21_C243_n1041, 
      mult_21_C243_n1040, mult_21_C243_n1039, mult_21_C243_n1038, 
      mult_21_C243_n1037, mult_21_C243_n1036, mult_21_C243_n1035, 
      mult_21_C243_n1034, mult_21_C243_n1033, mult_21_C243_n1032, 
      mult_21_C243_n1031, mult_21_C243_n1030, mult_21_C243_n1029, 
      mult_21_C243_n1028, mult_21_C243_n1027, mult_21_C243_n1026, 
      mult_21_C243_n1025, mult_21_C243_n1024, mult_21_C243_n1023, 
      mult_21_C243_n1022, mult_21_C243_n1021, mult_21_C243_n1020, 
      mult_21_C243_n1019, mult_21_C243_n1018, mult_21_C243_n1017, 
      mult_21_C243_n1016, mult_21_C243_n1015, mult_21_C243_n1014, 
      mult_21_C243_n1013, mult_21_C243_n1012, mult_21_C243_n1011, 
      mult_21_C243_n1010, mult_21_C243_n1009, mult_21_C243_n1008, 
      mult_21_C243_n1007, mult_21_C243_n1006, mult_21_C243_n1005, 
      mult_21_C243_n1004, mult_21_C243_n1003, mult_21_C243_n1002, 
      mult_21_C243_n1001, mult_21_C243_n1000, mult_21_C243_n999, 
      mult_21_C243_n998, mult_21_C243_n997, mult_21_C243_n996, 
      mult_21_C243_n995, mult_21_C243_n994, mult_21_C243_n993, 
      mult_21_C243_n992, mult_21_C243_n991, mult_21_C243_n990, 
      mult_21_C243_n989, mult_21_C243_n988, mult_21_C243_n987, 
      mult_21_C243_n986, mult_21_C243_n985, mult_21_C243_n984, 
      mult_21_C243_n983, mult_21_C243_n982, mult_21_C243_n981, 
      mult_21_C243_n980, mult_21_C243_n979, mult_21_C243_n978, 
      mult_21_C243_n977, mult_21_C243_n976, mult_21_C243_n975, 
      mult_21_C243_n974, mult_21_C243_n973, mult_21_C243_n972, 
      mult_21_C243_n971, mult_21_C243_n970, mult_21_C243_n969, 
      mult_21_C243_n968, mult_21_C243_n967, mult_21_C243_n966, 
      mult_21_C243_n965, mult_21_C243_n964, mult_21_C243_n963, 
      mult_21_C243_n962, mult_21_C243_n961, mult_21_C243_n960, 
      mult_21_C243_n959, mult_21_C243_n958, mult_21_C243_n957, 
      mult_21_C243_n956, mult_21_C243_n955, mult_21_C243_n954, 
      mult_21_C243_n953, mult_21_C243_n952, mult_21_C243_n951, 
      mult_21_C243_n950, mult_21_C243_n949, mult_21_C243_n948, 
      mult_21_C243_n947, mult_21_C243_n946, mult_21_C243_n945, 
      mult_21_C243_n944, mult_21_C243_n943, mult_21_C243_n942, 
      mult_21_C243_n941, mult_21_C243_n940, mult_21_C243_n939, 
      mult_21_C243_n938, mult_21_C243_n937, mult_21_C243_n936, 
      mult_21_C243_n935, mult_21_C243_n934, mult_21_C243_n933, 
      mult_21_C243_n932, mult_21_C243_n931, mult_21_C243_n930, 
      mult_21_C243_n929, mult_21_C243_n928, mult_21_C243_n927, 
      mult_21_C243_n926, mult_21_C243_n925, mult_21_C243_n924, 
      mult_21_C243_n923, mult_21_C243_n922, mult_21_C243_n921, 
      mult_21_C243_n920, mult_21_C243_n919, mult_21_C243_n918, 
      mult_21_C243_n917, mult_21_C243_n916, mult_21_C243_n915, 
      mult_21_C243_n914, mult_21_C243_n913, mult_21_C243_n912, 
      mult_21_C243_n911, mult_21_C243_n910, mult_21_C243_n909, 
      mult_21_C243_n908, mult_21_C243_n907, mult_21_C243_n906, 
      mult_21_C243_n905, mult_21_C243_n904, mult_21_C243_n903, 
      mult_21_C243_n902, mult_21_C243_n901, mult_21_C243_n900, 
      mult_21_C243_n899, mult_21_C243_n898, mult_21_C243_n897, 
      mult_21_C243_n896, mult_21_C243_n895, mult_21_C243_n894, 
      mult_21_C243_n893, mult_21_C243_n892, mult_21_C243_n891, 
      mult_21_C243_n890, mult_21_C243_n889, mult_21_C243_n888, 
      mult_21_C243_n887, mult_21_C243_n886, mult_21_C243_n885, 
      mult_21_C243_n884, mult_21_C243_n883, mult_21_C243_n882, 
      mult_21_C243_n881, mult_21_C243_n880, mult_21_C243_n879, 
      mult_21_C243_n878, mult_21_C243_n877, mult_21_C243_n876, 
      mult_21_C243_n875, mult_21_C243_n874, mult_21_C243_n873, 
      mult_21_C243_n872, mult_21_C243_n871, mult_21_C243_n870, 
      mult_21_C243_n869, mult_21_C243_n868, mult_21_C243_n867, 
      mult_21_C243_n866, mult_21_C243_n865, mult_21_C243_n864, 
      mult_21_C243_n863, mult_21_C243_n862, mult_21_C243_n861, 
      mult_21_C243_n860, mult_21_C243_n859, mult_21_C243_n858, 
      mult_21_C243_n857, mult_21_C243_n856, mult_21_C243_n855, 
      mult_21_C243_n854, mult_21_C243_n853, mult_21_C243_n852, 
      mult_21_C243_n851, mult_21_C243_n850, mult_21_C243_n849, 
      mult_21_C243_n848, mult_21_C243_n847, mult_21_C243_n846, 
      mult_21_C243_n845, mult_21_C243_n844, mult_21_C243_n843, 
      mult_21_C243_n842, mult_21_C243_n841, mult_21_C243_n840, 
      mult_21_C243_n839, mult_21_C243_n838, mult_21_C243_n837, 
      mult_21_C243_n836, mult_21_C243_n835, mult_21_C243_n834, 
      mult_21_C243_n833, mult_21_C243_n832, mult_21_C243_n831, 
      mult_21_C243_n830, mult_21_C243_n829, mult_21_C243_n828, 
      mult_21_C243_n827, mult_21_C243_n826, mult_21_C243_n825, 
      mult_21_C243_n824, mult_21_C243_n823, mult_21_C243_n822, 
      mult_21_C243_n821, mult_21_C243_n820, mult_21_C243_n819, 
      mult_21_C243_n818, mult_21_C243_n817, mult_21_C243_n816, 
      mult_21_C243_n815, mult_21_C243_n814, mult_21_C243_n813, 
      mult_21_C243_n812, mult_21_C243_n811, mult_21_C243_n810, 
      mult_21_C243_n809, mult_21_C243_n808, mult_21_C243_n807, 
      mult_21_C243_n806, mult_21_C243_n805, mult_21_C243_n804, 
      mult_21_C243_n803, mult_21_C243_n802, mult_21_C243_n801, 
      mult_21_C243_n800, mult_21_C243_n799, mult_21_C243_n798, 
      mult_21_C243_n797, mult_21_C243_n796, mult_21_C243_n795, 
      mult_21_C243_n794, mult_21_C243_n793, mult_21_C243_n792, 
      mult_21_C243_n791, mult_21_C243_n790, mult_21_C243_n789, 
      mult_21_C243_n788, mult_21_C243_n787, mult_21_C243_n786, 
      mult_21_C243_n785, mult_21_C243_n784, mult_21_C243_n783, 
      mult_21_C243_n782, mult_21_C243_n781, mult_21_C243_n780, 
      mult_21_C243_n779, mult_21_C243_n778, mult_21_C243_n777, 
      mult_21_C243_n776, mult_21_C243_n775, mult_21_C243_n774, 
      mult_21_C243_n773, mult_21_C243_n772, mult_21_C243_n771, 
      mult_21_C243_n770, mult_21_C243_n769, mult_21_C243_n768, 
      mult_21_C243_n767, mult_21_C243_n766, mult_21_C243_n765, 
      mult_21_C243_n764, mult_21_C243_n763, mult_21_C243_n762, 
      mult_21_C243_n761, mult_21_C243_n760, mult_21_C243_n759, 
      mult_21_C243_n758, mult_21_C243_n757, mult_21_C243_n756, 
      mult_21_C243_n755, mult_21_C243_n754, mult_21_C243_n753, 
      mult_21_C243_n752, mult_21_C243_n751, mult_21_C243_n750, 
      mult_21_C243_n749, mult_21_C243_n748, mult_21_C243_n747, 
      mult_21_C243_n746, mult_21_C243_n745, mult_21_C243_n744, 
      mult_21_C243_n743, mult_21_C243_n742, mult_21_C243_n741, 
      mult_21_C243_n740, mult_21_C243_n739, mult_21_C243_n738, 
      mult_21_C243_n737, mult_21_C243_n736, mult_21_C243_n735, 
      mult_21_C243_n734, mult_21_C243_n733, mult_21_C243_n732, 
      mult_21_C243_n731, mult_21_C243_n730, mult_21_C243_n729, 
      mult_21_C243_n728, mult_21_C243_n727, mult_21_C243_n726, 
      mult_21_C243_n725, mult_21_C243_n724, mult_21_C243_n723, 
      mult_21_C243_n722, mult_21_C243_n721, mult_21_C243_n720, 
      mult_21_C243_n719, mult_21_C243_n718, mult_21_C243_n717, 
      mult_21_C243_n716, mult_21_C243_n715, mult_21_C243_n714, 
      mult_21_C243_n713, mult_21_C243_n712, mult_21_C243_n711, 
      mult_21_C243_n710, mult_21_C243_n709, mult_21_C243_n708, 
      mult_21_C243_n707, mult_21_C243_n706, mult_21_C243_n705, 
      mult_21_C243_n704, mult_21_C243_n703, mult_21_C243_n702, 
      mult_21_C243_n701, mult_21_C243_n700, mult_21_C243_n699, 
      mult_21_C243_n698, mult_21_C243_n697, mult_21_C243_n696, 
      mult_21_C243_n695, mult_21_C243_n694, mult_21_C243_n693, 
      mult_21_C243_n692, mult_21_C243_n691, mult_21_C243_n690, 
      mult_21_C243_n689, mult_21_C243_n688, mult_21_C243_n687, 
      mult_21_C243_n686, mult_21_C243_n685, mult_21_C243_n684, 
      mult_21_C243_n683, mult_21_C243_n682, mult_21_C243_n681, 
      mult_21_C243_n680, mult_21_C243_n679, mult_21_C243_n678, 
      mult_21_C243_n677, mult_21_C243_n676, mult_21_C243_n675, 
      mult_21_C243_n674, mult_21_C243_n673, mult_21_C243_n672, 
      mult_21_C243_n671, mult_21_C243_n670, mult_21_C243_n669, 
      mult_21_C243_n668, mult_21_C243_n667, mult_21_C243_n666, 
      mult_21_C243_n665, mult_21_C243_n664, mult_21_C243_n663, 
      mult_21_C243_n662, mult_21_C243_n661, mult_21_C243_n660, 
      mult_21_C243_n659, mult_21_C243_n658, mult_21_C243_n657, 
      mult_21_C243_n656, mult_21_C243_n655, mult_21_C243_n654, 
      mult_21_C243_n653, mult_21_C243_n652, mult_21_C243_n651, 
      mult_21_C243_n650, mult_21_C243_n649, mult_21_C243_n648, 
      mult_21_C243_n647, mult_21_C243_n646, mult_21_C243_n645, 
      mult_21_C243_n644, mult_21_C243_n643, mult_21_C243_n642, 
      mult_21_C243_n641, mult_21_C243_n640, mult_21_C243_n639, 
      mult_21_C243_n638, mult_21_C243_n637, mult_21_C243_n636, 
      mult_21_C243_n635, mult_21_C243_n634, mult_21_C243_n633, 
      mult_21_C243_n632, mult_21_C243_n631, mult_21_C243_n630, 
      mult_21_C243_n629, mult_21_C243_n628, mult_21_C243_n627, 
      mult_21_C243_n626, mult_21_C243_n625, mult_21_C243_n624, 
      mult_21_C243_n623, mult_21_C243_n622, mult_21_C243_n621, 
      mult_21_C243_n620, mult_21_C243_n619, mult_21_C243_n618, 
      mult_21_C243_n617, mult_21_C243_n616, mult_21_C243_n615, 
      mult_21_C243_n614, mult_21_C243_n613, mult_21_C243_n612, 
      mult_21_C243_n611, mult_21_C243_n610, mult_21_C243_n609, 
      mult_21_C243_n608, mult_21_C243_n607, mult_21_C243_n606, 
      mult_21_C243_n605, mult_21_C243_n604, mult_21_C243_n603, 
      mult_21_C243_n602, mult_21_C243_n601, mult_21_C243_n600, 
      mult_21_C243_n599, mult_21_C243_n598, mult_21_C243_n597, 
      mult_21_C243_n596, mult_21_C243_n595, mult_21_C243_n594, 
      mult_21_C243_n593, mult_21_C243_n592, mult_21_C243_n591, 
      mult_21_C243_n590, mult_21_C243_n589, mult_21_C243_n588, 
      mult_21_C243_n587, mult_21_C243_n586, mult_21_C243_n585, 
      mult_21_C243_n584, mult_21_C243_n583, mult_21_C243_n582, 
      mult_21_C243_n581, mult_21_C243_n580, mult_21_C243_n579, 
      mult_21_C243_n578, mult_21_C243_n577, mult_21_C243_n576, 
      mult_21_C243_n575, mult_21_C243_n574, mult_21_C243_n573, 
      mult_21_C243_n572, mult_21_C243_n571, mult_21_C243_n570, 
      mult_21_C243_n569, mult_21_C243_n568, mult_21_C243_n567, 
      mult_21_C243_n566, mult_21_C243_n565, mult_21_C243_n564, 
      mult_21_C243_n563, mult_21_C243_n562, mult_21_C243_n561, 
      mult_21_C243_n560, mult_21_C243_n559, mult_21_C243_n558, 
      mult_21_C243_n557, mult_21_C243_n556, mult_21_C243_n555, 
      mult_21_C243_n554, mult_21_C243_n553, mult_21_C243_n552, 
      mult_21_C243_n551, mult_21_C243_n550, mult_21_C243_n549, 
      mult_21_C243_n548, mult_21_C243_n547, mult_21_C243_n546, 
      mult_21_C243_n545, mult_21_C243_n544, mult_21_C243_n543, 
      mult_21_C243_n542, mult_21_C243_n541, mult_21_C243_n540, 
      mult_21_C243_n539, mult_21_C243_n538, mult_21_C243_n537, 
      mult_21_C243_n536, mult_21_C243_n535, mult_21_C243_n534, 
      mult_21_C243_n533, mult_21_C243_n532, mult_21_C243_n531, 
      mult_21_C243_n530, mult_21_C243_n529, mult_21_C243_n528, 
      mult_21_C243_n527, mult_21_C243_n526, mult_21_C243_n525, 
      mult_21_C243_n524, mult_21_C243_n523, mult_21_C243_n522, 
      mult_21_C243_n521, mult_21_C243_n520, mult_21_C243_n519, 
      mult_21_C243_n518, mult_21_C243_n517, mult_21_C243_n516, 
      mult_21_C243_n515, mult_21_C243_n514, mult_21_C243_n513, 
      mult_21_C243_n512, mult_21_C243_n511, mult_21_C243_n510, 
      mult_21_C243_n509, mult_21_C243_n508, mult_21_C243_n507, 
      mult_21_C243_n506, mult_21_C243_n505, mult_21_C243_n504, 
      mult_21_C243_n503, mult_21_C243_n502, mult_21_C243_n501, 
      mult_21_C243_n500, mult_21_C243_n499, mult_21_C243_n498, 
      mult_21_C243_n497, mult_21_C243_n496, mult_21_C243_n495, 
      mult_21_C243_n494, mult_21_C243_n493, mult_21_C243_n492, 
      mult_21_C243_n491, mult_21_C243_n490, mult_21_C243_n489, 
      mult_21_C243_n488, mult_21_C243_n487, mult_21_C243_n486, 
      mult_21_C243_n485, mult_21_C243_n484, mult_21_C243_n483, 
      mult_21_C243_n482, mult_21_C243_n481, mult_21_C243_n480, 
      mult_21_C243_n479, mult_21_C243_n478, mult_21_C243_n477, 
      mult_21_C243_n476, mult_21_C243_n475, mult_21_C243_n474, 
      mult_21_C243_n473, mult_21_C243_n472, mult_21_C243_n471, 
      mult_21_C243_n470, mult_21_C243_n469, mult_21_C243_n468, 
      mult_21_C243_n467, mult_21_C243_n466, mult_21_C243_n465, 
      mult_21_C243_n464, mult_21_C243_n463, mult_21_C243_n462, 
      mult_21_C243_n461, mult_21_C243_n460, mult_21_C243_n459, 
      mult_21_C243_n458, mult_21_C243_n457, mult_21_C243_n456, 
      mult_21_C243_n455, mult_21_C243_n454, mult_21_C243_n453, 
      mult_21_C243_n452, mult_21_C243_n451, mult_21_C243_n450, 
      mult_21_C243_n449, mult_21_C243_n448, mult_21_C243_n447, 
      mult_21_C243_n446, mult_21_C243_n445, mult_21_C243_n444, 
      mult_21_C243_n443, mult_21_C243_n442, mult_21_C243_n441, 
      mult_21_C243_n440, mult_21_C243_n439, mult_21_C243_n438, 
      mult_21_C243_n437, mult_21_C243_n436, mult_21_C243_n435, 
      mult_21_C243_n434, mult_21_C243_n433, mult_21_C243_n432, 
      mult_21_C243_n431, mult_21_C243_n430, mult_21_C243_n429, 
      mult_21_C243_n428, mult_21_C243_n427, mult_21_C243_n426, 
      mult_21_C243_n425, mult_21_C243_n424, mult_21_C243_n423, 
      mult_21_C243_n422, mult_21_C243_n421, mult_21_C243_n420, 
      mult_21_C243_n419, mult_21_C243_n418, mult_21_C243_n417, 
      mult_21_C243_n416, mult_21_C243_n415, mult_21_C243_n414, 
      mult_21_C243_n413, mult_21_C243_n412, mult_21_C243_n411, 
      mult_21_C243_n410, mult_21_C243_n409, mult_21_C243_n408, 
      mult_21_C243_n407, mult_21_C243_n406, mult_21_C243_n405, 
      mult_21_C243_n404, mult_21_C243_n403, mult_21_C243_n402, 
      mult_21_C243_n401, mult_21_C243_n400, mult_21_C243_n399, 
      mult_21_C243_n398, mult_21_C243_n397, mult_21_C243_n396, 
      mult_21_C243_n395, mult_21_C243_n394, mult_21_C243_n393, 
      mult_21_C243_n392, mult_21_C243_n391, mult_21_C243_n390, 
      mult_21_C243_n389, mult_21_C243_n388, mult_21_C243_n387, 
      mult_21_C243_n386, mult_21_C243_n385, mult_21_C243_n384, 
      mult_21_C243_n383, mult_21_C243_n382, mult_21_C243_n381, 
      mult_21_C243_n380, mult_21_C243_n379, mult_21_C243_n378, 
      mult_21_C243_n377, mult_21_C243_n376, mult_21_C243_n375, 
      mult_21_C243_n374, mult_21_C243_n373, mult_21_C243_n372, 
      mult_21_C243_n371, mult_21_C243_n370, mult_21_C243_n369, 
      mult_21_C243_n368, mult_21_C243_n367, mult_21_C243_n366, 
      mult_21_C243_n365, mult_21_C243_n364, mult_21_C243_n363, 
      mult_21_C243_n362, mult_21_C243_n361, mult_21_C243_n360, 
      mult_21_C243_n359, mult_21_C243_n358, mult_21_C243_n357, 
      mult_21_C243_n356, mult_21_C243_n355, mult_21_C243_n354, 
      mult_21_C243_n353, mult_21_C243_n352, mult_21_C243_n351, 
      mult_21_C243_n350, mult_21_C243_n349, mult_21_C243_n348, 
      mult_21_C243_n347, mult_21_C243_n346, mult_21_C243_n345, 
      mult_21_C243_n344, mult_21_C243_n343, mult_21_C243_n342, 
      mult_21_C243_n341, mult_21_C243_n340, mult_21_C243_n339, 
      mult_21_C243_n338, mult_21_C243_n337, mult_21_C243_n336, 
      mult_21_C243_n335, mult_21_C243_n334, mult_21_C243_n333, 
      mult_21_C243_n332, mult_21_C243_n331, mult_21_C243_n330, 
      mult_21_C243_n329, mult_21_C243_n326, mult_21_C243_n324, 
      mult_21_C243_n323, mult_21_C243_n322, mult_21_C243_n319, 
      mult_21_C243_n318, mult_21_C243_n315, mult_21_C243_n314, 
      mult_21_C243_n313, mult_21_C243_n312, mult_21_C243_n310, 
      mult_21_C243_n305, mult_21_C243_n303, mult_21_C243_n302, 
      mult_21_C243_n301, mult_21_C243_n297, mult_21_C243_n296, 
      mult_21_C243_n295, mult_21_C243_n294, mult_21_C243_n293, 
      mult_21_C243_n289, mult_21_C243_n288, mult_21_C243_n287, 
      mult_21_C243_n286, mult_21_C243_n285, mult_21_C243_n284, 
      mult_21_C243_n283, mult_21_C243_n282, mult_21_C243_n281, 
      mult_21_C243_n280, mult_21_C243_n279, mult_21_C243_n278, 
      mult_21_C243_n277, mult_21_C243_n276, mult_21_C243_n275, 
      mult_21_C243_n273, mult_21_C243_n271, mult_21_C243_n270, 
      mult_21_C243_n268, mult_21_C243_n266, mult_21_C243_n265, 
      mult_21_C243_n264, mult_21_C243_n263, mult_21_C243_n262, 
      mult_21_C243_n261, mult_21_C243_n260, mult_21_C243_n259, 
      mult_21_C243_n258, mult_21_C243_n257, mult_21_C243_n256, 
      mult_21_C243_n255, mult_21_C243_n254, mult_21_C243_n253, 
      mult_21_C243_n251, mult_21_C243_n249, mult_21_C243_n248, 
      mult_21_C243_n246, mult_21_C243_n244, mult_21_C243_n243, 
      mult_21_C243_n242, mult_21_C243_n241, mult_21_C243_n240, 
      mult_21_C243_n239, mult_21_C243_n238, mult_21_C243_n237, 
      mult_21_C243_n236, mult_21_C243_n235, mult_21_C243_n234, 
      mult_21_C243_n233, mult_21_C243_n232, mult_21_C243_n231, 
      mult_21_C243_n230, mult_21_C243_n229, mult_21_C243_n227, 
      mult_21_C243_n226, mult_21_C243_n225, mult_21_C243_n224, 
      mult_21_C243_n223, mult_21_C243_n222, mult_21_C243_n221, 
      mult_21_C243_n219, mult_21_C243_n217, mult_21_C243_n216, 
      mult_21_C243_n215, mult_21_C243_n214, mult_21_C243_n211, 
      mult_21_C243_n209, mult_21_C243_n208, mult_21_C243_n207, 
      mult_21_C243_n206, mult_21_C243_n204, mult_21_C243_n202, 
      mult_21_C243_n201, mult_21_C243_n200, mult_21_C243_n199, 
      mult_21_C243_n197, mult_21_C243_n195, mult_21_C243_n194, 
      mult_21_C243_n190, mult_21_C243_n189, mult_21_C243_n188, 
      mult_21_C243_n187, mult_21_C243_n185, mult_21_C243_n184, 
      mult_21_C243_n183, mult_21_C243_n182, mult_21_C243_n181, 
      mult_21_C243_n180, mult_21_C243_n179, mult_21_C243_n178, 
      mult_21_C243_n176, mult_21_C243_n175, mult_21_C243_n174, 
      mult_21_C243_n173, mult_21_C243_n172, mult_21_C243_n171, 
      mult_21_C243_n170, mult_21_C243_n169, mult_21_C243_n168, 
      mult_21_C243_n167, mult_21_C243_n166, mult_21_C243_n165, 
      mult_21_C243_n164, mult_21_C243_n163, mult_21_C243_n162, 
      mult_21_C243_n161, mult_21_C243_n160, mult_21_C243_n159, 
      mult_21_C243_n158, mult_21_C243_n157, mult_21_C243_n156, 
      mult_21_C243_n155, mult_21_C243_n106, mult_21_C243_n105, 
      mult_21_C243_n104, mult_21_C243_n103, mult_21_C243_n101, mult_21_C243_n99
      , mult_21_C243_n98, mult_21_C243_n96, mult_21_C243_n94, mult_21_C243_n93,
      mult_21_C243_n91, mult_21_C243_n89, mult_21_C243_n88, mult_21_C243_n86, 
      mult_21_C243_n84, mult_21_C243_n83, mult_21_C243_n81, mult_21_C243_n79, 
      mult_21_C243_n78, mult_21_C243_n76, mult_21_C243_n73, mult_21_C243_n71, 
      mult_21_C243_n69, mult_21_C243_n66, mult_21_C243_n63, mult_21_C243_n61, 
      mult_21_C243_n58, mult_21_C243_n56, mult_21_C243_n53, mult_21_C243_n50, 
      mult_21_C243_n48, mult_21_C243_n45, mult_21_C243_n42, mult_21_C243_n38, 
      mult_21_C243_n30, mult_21_C243_n22, mult_21_C243_n14, mult_21_C243_n8, 
      mult_21_C243_n6, mult_21_C243_n3, mult_21_C245_n1544, mult_21_C245_n1543,
      mult_21_C245_n1542, mult_21_C245_n1541, mult_21_C245_n1540, 
      mult_21_C245_n1539, mult_21_C245_n1538, mult_21_C245_n1537, 
      mult_21_C245_n1536, mult_21_C245_n1535, mult_21_C245_n1534, 
      mult_21_C245_n1533, mult_21_C245_n1532, mult_21_C245_n1531, 
      mult_21_C245_n1530, mult_21_C245_n1529, mult_21_C245_n1528, 
      mult_21_C245_n1527, mult_21_C245_n1526, mult_21_C245_n1525, 
      mult_21_C245_n1524, mult_21_C245_n1523, mult_21_C245_n1522, 
      mult_21_C245_n1521, mult_21_C245_n1519, mult_21_C245_n1518, 
      mult_21_C245_n1517, mult_21_C245_n1368, mult_21_C245_n1367, 
      mult_21_C245_n1366, mult_21_C245_n1365, mult_21_C245_n1364, 
      mult_21_C245_n1363, mult_21_C245_n1362, mult_21_C245_n1361, 
      mult_21_C245_n1360, mult_21_C245_n1359, mult_21_C245_n1358, 
      mult_21_C245_n1357, mult_21_C245_n1356, mult_21_C245_n1355, 
      mult_21_C245_n1354, mult_21_C245_n1353, mult_21_C245_n1352, 
      mult_21_C245_n1351, mult_21_C245_n1350, mult_21_C245_n1349, 
      mult_21_C245_n1348, mult_21_C245_n1347, mult_21_C245_n1346, 
      mult_21_C245_n1345, mult_21_C245_n1344, mult_21_C245_n1343, 
      mult_21_C245_n1342, mult_21_C245_n1341, mult_21_C245_n1340, 
      mult_21_C245_n1339, mult_21_C245_n1338, mult_21_C245_n1337, 
      mult_21_C245_n1336, mult_21_C245_n1335, mult_21_C245_n1334, 
      mult_21_C245_n1333, mult_21_C245_n1332, mult_21_C245_n1331, 
      mult_21_C245_n1330, mult_21_C245_n1329, mult_21_C245_n1328, 
      mult_21_C245_n1327, mult_21_C245_n1326, mult_21_C245_n1325, 
      mult_21_C245_n1324, mult_21_C245_n1323, mult_21_C245_n1322, 
      mult_21_C245_n1321, mult_21_C245_n1320, mult_21_C245_n1319, 
      mult_21_C245_n1318, mult_21_C245_n1317, mult_21_C245_n1316, 
      mult_21_C245_n1315, mult_21_C245_n1314, mult_21_C245_n1313, 
      mult_21_C245_n1312, mult_21_C245_n1311, mult_21_C245_n1310, 
      mult_21_C245_n1309, mult_21_C245_n1308, mult_21_C245_n1307, 
      mult_21_C245_n1306, mult_21_C245_n1305, mult_21_C245_n1304, 
      mult_21_C245_n1303, mult_21_C245_n1302, mult_21_C245_n1301, 
      mult_21_C245_n1300, mult_21_C245_n1299, mult_21_C245_n1298, 
      mult_21_C245_n1297, mult_21_C245_n1296, mult_21_C245_n1295, 
      mult_21_C245_n1294, mult_21_C245_n1293, mult_21_C245_n1292, 
      mult_21_C245_n1291, mult_21_C245_n1290, mult_21_C245_n1289, 
      mult_21_C245_n1288, mult_21_C245_n1287, mult_21_C245_n1286, 
      mult_21_C245_n1285, mult_21_C245_n1284, mult_21_C245_n1283, 
      mult_21_C245_n1282, mult_21_C245_n1281, mult_21_C245_n1280, 
      mult_21_C245_n1279, mult_21_C245_n1278, mult_21_C245_n1277, 
      mult_21_C245_n1276, mult_21_C245_n1275, mult_21_C245_n1274, 
      mult_21_C245_n1273, mult_21_C245_n1272, mult_21_C245_n1271, 
      mult_21_C245_n1270, mult_21_C245_n1269, mult_21_C245_n1268, 
      mult_21_C245_n1267, mult_21_C245_n1266, mult_21_C245_n1265, 
      mult_21_C245_n1264, mult_21_C245_n1263, mult_21_C245_n1262, 
      mult_21_C245_n1261, mult_21_C245_n1260, mult_21_C245_n1259, 
      mult_21_C245_n1258, mult_21_C245_n1257, mult_21_C245_n1256, 
      mult_21_C245_n1255, mult_21_C245_n1254, mult_21_C245_n1253, 
      mult_21_C245_n1252, mult_21_C245_n1251, mult_21_C245_n1250, 
      mult_21_C245_n1249, mult_21_C245_n1248, mult_21_C245_n1247, 
      mult_21_C245_n1246, mult_21_C245_n1245, mult_21_C245_n1244, 
      mult_21_C245_n1243, mult_21_C245_n1242, mult_21_C245_n1241, 
      mult_21_C245_n1240, mult_21_C245_n1239, mult_21_C245_n1238, 
      mult_21_C245_n1237, mult_21_C245_n1236, mult_21_C245_n1235, 
      mult_21_C245_n1234, mult_21_C245_n1233, mult_21_C245_n1232, 
      mult_21_C245_n1231, mult_21_C245_n1230, mult_21_C245_n1229, 
      mult_21_C245_n1228, mult_21_C245_n1227, mult_21_C245_n1226, 
      mult_21_C245_n1225, mult_21_C245_n1224, mult_21_C245_n1223, 
      mult_21_C245_n1222, mult_21_C245_n1221, mult_21_C245_n1220, 
      mult_21_C245_n1219, mult_21_C245_n1218, mult_21_C245_n1217, 
      mult_21_C245_n1216, mult_21_C245_n1215, mult_21_C245_n1214, 
      mult_21_C245_n1213, mult_21_C245_n1212, mult_21_C245_n1211, 
      mult_21_C245_n1210, mult_21_C245_n1209, mult_21_C245_n1208, 
      mult_21_C245_n1207, mult_21_C245_n1206, mult_21_C245_n1205, 
      mult_21_C245_n1204, mult_21_C245_n1203, mult_21_C245_n1202, 
      mult_21_C245_n1201, mult_21_C245_n1200, mult_21_C245_n1199, 
      mult_21_C245_n1198, mult_21_C245_n1197, mult_21_C245_n1196, 
      mult_21_C245_n1195, mult_21_C245_n1194, mult_21_C245_n1193, 
      mult_21_C245_n1192, mult_21_C245_n1191, mult_21_C245_n1190, 
      mult_21_C245_n1189, mult_21_C245_n1188, mult_21_C245_n1187, 
      mult_21_C245_n1186, mult_21_C245_n1185, mult_21_C245_n1184, 
      mult_21_C245_n1183, mult_21_C245_n1182, mult_21_C245_n1181, 
      mult_21_C245_n1180, mult_21_C245_n1179, mult_21_C245_n1178, 
      mult_21_C245_n1177, mult_21_C245_n1176, mult_21_C245_n1175, 
      mult_21_C245_n1174, mult_21_C245_n1173, mult_21_C245_n1172, 
      mult_21_C245_n1171, mult_21_C245_n1170, mult_21_C245_n1169, 
      mult_21_C245_n1168, mult_21_C245_n1167, mult_21_C245_n1166, 
      mult_21_C245_n1165, mult_21_C245_n1164, mult_21_C245_n1163, 
      mult_21_C245_n1162, mult_21_C245_n1161, mult_21_C245_n1160, 
      mult_21_C245_n1159, mult_21_C245_n1158, mult_21_C245_n1157, 
      mult_21_C245_n1156, mult_21_C245_n1155, mult_21_C245_n1154, 
      mult_21_C245_n1153, mult_21_C245_n1152, mult_21_C245_n1151, 
      mult_21_C245_n1150, mult_21_C245_n1149, mult_21_C245_n1148, 
      mult_21_C245_n1147, mult_21_C245_n1146, mult_21_C245_n1145, 
      mult_21_C245_n1144, mult_21_C245_n1143, mult_21_C245_n1142, 
      mult_21_C245_n1141, mult_21_C245_n1140, mult_21_C245_n1139, 
      mult_21_C245_n1138, mult_21_C245_n1137, mult_21_C245_n1136, 
      mult_21_C245_n1135, mult_21_C245_n1134, mult_21_C245_n1133, 
      mult_21_C245_n1132, mult_21_C245_n1131, mult_21_C245_n1130, 
      mult_21_C245_n1129, mult_21_C245_n1128, mult_21_C245_n1127, 
      mult_21_C245_n1126, mult_21_C245_n1125, mult_21_C245_n1124, 
      mult_21_C245_n1123, mult_21_C245_n1122, mult_21_C245_n1121, 
      mult_21_C245_n1120, mult_21_C245_n1119, mult_21_C245_n1118, 
      mult_21_C245_n1117, mult_21_C245_n1116, mult_21_C245_n1115, 
      mult_21_C245_n1114, mult_21_C245_n1113, mult_21_C245_n1112, 
      mult_21_C245_n1111, mult_21_C245_n1110, mult_21_C245_n1109, 
      mult_21_C245_n1108, mult_21_C245_n1107, mult_21_C245_n1106, 
      mult_21_C245_n1105, mult_21_C245_n1104, mult_21_C245_n1103, 
      mult_21_C245_n1102, mult_21_C245_n1101, mult_21_C245_n1100, 
      mult_21_C245_n1099, mult_21_C245_n1098, mult_21_C245_n1097, 
      mult_21_C245_n1096, mult_21_C245_n1095, mult_21_C245_n1094, 
      mult_21_C245_n1093, mult_21_C245_n1092, mult_21_C245_n1091, 
      mult_21_C245_n1090, mult_21_C245_n1089, mult_21_C245_n1088, 
      mult_21_C245_n1087, mult_21_C245_n1086, mult_21_C245_n1085, 
      mult_21_C245_n1084, mult_21_C245_n1083, mult_21_C245_n1082, 
      mult_21_C245_n1081, mult_21_C245_n1080, mult_21_C245_n1079, 
      mult_21_C245_n1078, mult_21_C245_n1077, mult_21_C245_n1076, 
      mult_21_C245_n1075, mult_21_C245_n1074, mult_21_C245_n1073, 
      mult_21_C245_n1072, mult_21_C245_n1071, mult_21_C245_n1070, 
      mult_21_C245_n1069, mult_21_C245_n1068, mult_21_C245_n1067, 
      mult_21_C245_n1066, mult_21_C245_n1065, mult_21_C245_n1064, 
      mult_21_C245_n1063, mult_21_C245_n1062, mult_21_C245_n1061, 
      mult_21_C245_n1060, mult_21_C245_n1059, mult_21_C245_n1058, 
      mult_21_C245_n1057, mult_21_C245_n1056, mult_21_C245_n1055, 
      mult_21_C245_n1054, mult_21_C245_n1053, mult_21_C245_n1052, 
      mult_21_C245_n1051, mult_21_C245_n1050, mult_21_C245_n1049, 
      mult_21_C245_n1048, mult_21_C245_n1047, mult_21_C245_n1046, 
      mult_21_C245_n1045, mult_21_C245_n1044, mult_21_C245_n1043, 
      mult_21_C245_n1042, mult_21_C245_n1041, mult_21_C245_n1040, 
      mult_21_C245_n1039, mult_21_C245_n1038, mult_21_C245_n1037, 
      mult_21_C245_n1036, mult_21_C245_n1035, mult_21_C245_n1034, 
      mult_21_C245_n1033, mult_21_C245_n1032, mult_21_C245_n1031, 
      mult_21_C245_n1030, mult_21_C245_n1029, mult_21_C245_n1028, 
      mult_21_C245_n1027, mult_21_C245_n1026, mult_21_C245_n1025, 
      mult_21_C245_n1024, mult_21_C245_n1023, mult_21_C245_n1022, 
      mult_21_C245_n1021, mult_21_C245_n1020, mult_21_C245_n1019, 
      mult_21_C245_n1018, mult_21_C245_n1017, mult_21_C245_n1016, 
      mult_21_C245_n1015, mult_21_C245_n1014, mult_21_C245_n1013, 
      mult_21_C245_n1012, mult_21_C245_n1011, mult_21_C245_n1010, 
      mult_21_C245_n1009, mult_21_C245_n1008, mult_21_C245_n1007, 
      mult_21_C245_n1006, mult_21_C245_n1005, mult_21_C245_n1004, 
      mult_21_C245_n1003, mult_21_C245_n1002, mult_21_C245_n1001, 
      mult_21_C245_n1000, mult_21_C245_n999, mult_21_C245_n998, 
      mult_21_C245_n997, mult_21_C245_n996, mult_21_C245_n995, 
      mult_21_C245_n994, mult_21_C245_n993, mult_21_C245_n992, 
      mult_21_C245_n991, mult_21_C245_n990, mult_21_C245_n989, 
      mult_21_C245_n988, mult_21_C245_n987, mult_21_C245_n986, 
      mult_21_C245_n985, mult_21_C245_n984, mult_21_C245_n983, 
      mult_21_C245_n982, mult_21_C245_n981, mult_21_C245_n980, 
      mult_21_C245_n979, mult_21_C245_n978, mult_21_C245_n977, 
      mult_21_C245_n976, mult_21_C245_n975, mult_21_C245_n974, 
      mult_21_C245_n973, mult_21_C245_n972, mult_21_C245_n971, 
      mult_21_C245_n970, mult_21_C245_n969, mult_21_C245_n968, 
      mult_21_C245_n967, mult_21_C245_n966, mult_21_C245_n965, 
      mult_21_C245_n964, mult_21_C245_n963, mult_21_C245_n962, 
      mult_21_C245_n961, mult_21_C245_n960, mult_21_C245_n959, 
      mult_21_C245_n958, mult_21_C245_n957, mult_21_C245_n956, 
      mult_21_C245_n955, mult_21_C245_n954, mult_21_C245_n953, 
      mult_21_C245_n952, mult_21_C245_n951, mult_21_C245_n950, 
      mult_21_C245_n949, mult_21_C245_n948, mult_21_C245_n947, 
      mult_21_C245_n946, mult_21_C245_n945, mult_21_C245_n944, 
      mult_21_C245_n943, mult_21_C245_n942, mult_21_C245_n941, 
      mult_21_C245_n940, mult_21_C245_n939, mult_21_C245_n938, 
      mult_21_C245_n937, mult_21_C245_n936, mult_21_C245_n935, 
      mult_21_C245_n934, mult_21_C245_n933, mult_21_C245_n932, 
      mult_21_C245_n931, mult_21_C245_n930, mult_21_C245_n929, 
      mult_21_C245_n928, mult_21_C245_n927, mult_21_C245_n926, 
      mult_21_C245_n925, mult_21_C245_n924, mult_21_C245_n923, 
      mult_21_C245_n922, mult_21_C245_n921, mult_21_C245_n920, 
      mult_21_C245_n919, mult_21_C245_n918, mult_21_C245_n917, 
      mult_21_C245_n916, mult_21_C245_n915, mult_21_C245_n914, 
      mult_21_C245_n913, mult_21_C245_n912, mult_21_C245_n911, 
      mult_21_C245_n910, mult_21_C245_n909, mult_21_C245_n908, 
      mult_21_C245_n907, mult_21_C245_n906, mult_21_C245_n905, 
      mult_21_C245_n904, mult_21_C245_n903, mult_21_C245_n902, 
      mult_21_C245_n901, mult_21_C245_n900, mult_21_C245_n899, 
      mult_21_C245_n898, mult_21_C245_n897, mult_21_C245_n896, 
      mult_21_C245_n895, mult_21_C245_n894, mult_21_C245_n893, 
      mult_21_C245_n892, mult_21_C245_n891, mult_21_C245_n890, 
      mult_21_C245_n889, mult_21_C245_n888, mult_21_C245_n887, 
      mult_21_C245_n886, mult_21_C245_n885, mult_21_C245_n884, 
      mult_21_C245_n883, mult_21_C245_n882, mult_21_C245_n881, 
      mult_21_C245_n880, mult_21_C245_n879, mult_21_C245_n878, 
      mult_21_C245_n877, mult_21_C245_n876, mult_21_C245_n875, 
      mult_21_C245_n874, mult_21_C245_n873, mult_21_C245_n872, 
      mult_21_C245_n871, mult_21_C245_n870, mult_21_C245_n869, 
      mult_21_C245_n868, mult_21_C245_n867, mult_21_C245_n866, 
      mult_21_C245_n865, mult_21_C245_n864, mult_21_C245_n863, 
      mult_21_C245_n862, mult_21_C245_n861, mult_21_C245_n860, 
      mult_21_C245_n859, mult_21_C245_n858, mult_21_C245_n857, 
      mult_21_C245_n856, mult_21_C245_n855, mult_21_C245_n854, 
      mult_21_C245_n853, mult_21_C245_n852, mult_21_C245_n851, 
      mult_21_C245_n850, mult_21_C245_n849, mult_21_C245_n848, 
      mult_21_C245_n847, mult_21_C245_n846, mult_21_C245_n845, 
      mult_21_C245_n844, mult_21_C245_n843, mult_21_C245_n842, 
      mult_21_C245_n841, mult_21_C245_n840, mult_21_C245_n839, 
      mult_21_C245_n838, mult_21_C245_n837, mult_21_C245_n836, 
      mult_21_C245_n835, mult_21_C245_n834, mult_21_C245_n833, 
      mult_21_C245_n832, mult_21_C245_n831, mult_21_C245_n830, 
      mult_21_C245_n829, mult_21_C245_n828, mult_21_C245_n827, 
      mult_21_C245_n826, mult_21_C245_n825, mult_21_C245_n824, 
      mult_21_C245_n823, mult_21_C245_n822, mult_21_C245_n821, 
      mult_21_C245_n820, mult_21_C245_n819, mult_21_C245_n818, 
      mult_21_C245_n817, mult_21_C245_n816, mult_21_C245_n815, 
      mult_21_C245_n814, mult_21_C245_n813, mult_21_C245_n812, 
      mult_21_C245_n811, mult_21_C245_n810, mult_21_C245_n809, 
      mult_21_C245_n808, mult_21_C245_n807, mult_21_C245_n806, 
      mult_21_C245_n805, mult_21_C245_n804, mult_21_C245_n803, 
      mult_21_C245_n802, mult_21_C245_n801, mult_21_C245_n800, 
      mult_21_C245_n799, mult_21_C245_n798, mult_21_C245_n797, 
      mult_21_C245_n796, mult_21_C245_n795, mult_21_C245_n794, 
      mult_21_C245_n793, mult_21_C245_n792, mult_21_C245_n791, 
      mult_21_C245_n790, mult_21_C245_n789, mult_21_C245_n788, 
      mult_21_C245_n787, mult_21_C245_n786, mult_21_C245_n785, 
      mult_21_C245_n784, mult_21_C245_n783, mult_21_C245_n782, 
      mult_21_C245_n781, mult_21_C245_n780, mult_21_C245_n779, 
      mult_21_C245_n778, mult_21_C245_n777, mult_21_C245_n776, 
      mult_21_C245_n775, mult_21_C245_n774, mult_21_C245_n773, 
      mult_21_C245_n772, mult_21_C245_n771, mult_21_C245_n770, 
      mult_21_C245_n769, mult_21_C245_n768, mult_21_C245_n767, 
      mult_21_C245_n766, mult_21_C245_n765, mult_21_C245_n764, 
      mult_21_C245_n763, mult_21_C245_n762, mult_21_C245_n761, 
      mult_21_C245_n760, mult_21_C245_n759, mult_21_C245_n758, 
      mult_21_C245_n757, mult_21_C245_n756, mult_21_C245_n755, 
      mult_21_C245_n754, mult_21_C245_n753, mult_21_C245_n752, 
      mult_21_C245_n751, mult_21_C245_n750, mult_21_C245_n749, 
      mult_21_C245_n748, mult_21_C245_n747, mult_21_C245_n746, 
      mult_21_C245_n745, mult_21_C245_n744, mult_21_C245_n743, 
      mult_21_C245_n742, mult_21_C245_n741, mult_21_C245_n740, 
      mult_21_C245_n739, mult_21_C245_n738, mult_21_C245_n737, 
      mult_21_C245_n736, mult_21_C245_n735, mult_21_C245_n734, 
      mult_21_C245_n733, mult_21_C245_n732, mult_21_C245_n731, 
      mult_21_C245_n730, mult_21_C245_n729, mult_21_C245_n728, 
      mult_21_C245_n727, mult_21_C245_n726, mult_21_C245_n725, 
      mult_21_C245_n724, mult_21_C245_n723, mult_21_C245_n722, 
      mult_21_C245_n721, mult_21_C245_n720, mult_21_C245_n719, 
      mult_21_C245_n718, mult_21_C245_n717, mult_21_C245_n716, 
      mult_21_C245_n715, mult_21_C245_n714, mult_21_C245_n713, 
      mult_21_C245_n712, mult_21_C245_n711, mult_21_C245_n710, 
      mult_21_C245_n709, mult_21_C245_n708, mult_21_C245_n707, 
      mult_21_C245_n706, mult_21_C245_n705, mult_21_C245_n704, 
      mult_21_C245_n703, mult_21_C245_n702, mult_21_C245_n701, 
      mult_21_C245_n700, mult_21_C245_n699, mult_21_C245_n698, 
      mult_21_C245_n697, mult_21_C245_n696, mult_21_C245_n695, 
      mult_21_C245_n694, mult_21_C245_n693, mult_21_C245_n692, 
      mult_21_C245_n691, mult_21_C245_n690, mult_21_C245_n689, 
      mult_21_C245_n688, mult_21_C245_n687, mult_21_C245_n686, 
      mult_21_C245_n685, mult_21_C245_n684, mult_21_C245_n683, 
      mult_21_C245_n682, mult_21_C245_n681, mult_21_C245_n680, 
      mult_21_C245_n679, mult_21_C245_n678, mult_21_C245_n677, 
      mult_21_C245_n676, mult_21_C245_n675, mult_21_C245_n674, 
      mult_21_C245_n673, mult_21_C245_n672, mult_21_C245_n671, 
      mult_21_C245_n670, mult_21_C245_n669, mult_21_C245_n668, 
      mult_21_C245_n667, mult_21_C245_n666, mult_21_C245_n665, 
      mult_21_C245_n664, mult_21_C245_n663, mult_21_C245_n662, 
      mult_21_C245_n661, mult_21_C245_n660, mult_21_C245_n659, 
      mult_21_C245_n658, mult_21_C245_n657, mult_21_C245_n656, 
      mult_21_C245_n655, mult_21_C245_n654, mult_21_C245_n653, 
      mult_21_C245_n652, mult_21_C245_n651, mult_21_C245_n650, 
      mult_21_C245_n649, mult_21_C245_n648, mult_21_C245_n647, 
      mult_21_C245_n646, mult_21_C245_n645, mult_21_C245_n644, 
      mult_21_C245_n643, mult_21_C245_n642, mult_21_C245_n641, 
      mult_21_C245_n640, mult_21_C245_n639, mult_21_C245_n638, 
      mult_21_C245_n637, mult_21_C245_n636, mult_21_C245_n635, 
      mult_21_C245_n634, mult_21_C245_n633, mult_21_C245_n632, 
      mult_21_C245_n631, mult_21_C245_n630, mult_21_C245_n629, 
      mult_21_C245_n628, mult_21_C245_n627, mult_21_C245_n626, 
      mult_21_C245_n625, mult_21_C245_n624, mult_21_C245_n623, 
      mult_21_C245_n622, mult_21_C245_n621, mult_21_C245_n620, 
      mult_21_C245_n619, mult_21_C245_n618, mult_21_C245_n617, 
      mult_21_C245_n616, mult_21_C245_n615, mult_21_C245_n614, 
      mult_21_C245_n613, mult_21_C245_n612, mult_21_C245_n611, 
      mult_21_C245_n610, mult_21_C245_n609, mult_21_C245_n608, 
      mult_21_C245_n607, mult_21_C245_n606, mult_21_C245_n605, 
      mult_21_C245_n604, mult_21_C245_n603, mult_21_C245_n602, 
      mult_21_C245_n601, mult_21_C245_n600, mult_21_C245_n599, 
      mult_21_C245_n598, mult_21_C245_n597, mult_21_C245_n596, 
      mult_21_C245_n595, mult_21_C245_n594, mult_21_C245_n593, 
      mult_21_C245_n592, mult_21_C245_n591, mult_21_C245_n590, 
      mult_21_C245_n589, mult_21_C245_n588, mult_21_C245_n587, 
      mult_21_C245_n586, mult_21_C245_n585, mult_21_C245_n584, 
      mult_21_C245_n583, mult_21_C245_n582, mult_21_C245_n581, 
      mult_21_C245_n580, mult_21_C245_n579, mult_21_C245_n578, 
      mult_21_C245_n577, mult_21_C245_n576, mult_21_C245_n575, 
      mult_21_C245_n574, mult_21_C245_n573, mult_21_C245_n572, 
      mult_21_C245_n571, mult_21_C245_n570, mult_21_C245_n569, 
      mult_21_C245_n568, mult_21_C245_n567, mult_21_C245_n566, 
      mult_21_C245_n565, mult_21_C245_n564, mult_21_C245_n563, 
      mult_21_C245_n562, mult_21_C245_n561, mult_21_C245_n560, 
      mult_21_C245_n559, mult_21_C245_n558, mult_21_C245_n557, 
      mult_21_C245_n556, mult_21_C245_n555, mult_21_C245_n554, 
      mult_21_C245_n553, mult_21_C245_n552, mult_21_C245_n551, 
      mult_21_C245_n550, mult_21_C245_n549, mult_21_C245_n548, 
      mult_21_C245_n547, mult_21_C245_n546, mult_21_C245_n545, 
      mult_21_C245_n544, mult_21_C245_n543, mult_21_C245_n542, 
      mult_21_C245_n541, mult_21_C245_n540, mult_21_C245_n539, 
      mult_21_C245_n538, mult_21_C245_n537, mult_21_C245_n536, 
      mult_21_C245_n535, mult_21_C245_n534, mult_21_C245_n533, 
      mult_21_C245_n532, mult_21_C245_n531, mult_21_C245_n530, 
      mult_21_C245_n529, mult_21_C245_n528, mult_21_C245_n527, 
      mult_21_C245_n526, mult_21_C245_n525, mult_21_C245_n524, 
      mult_21_C245_n523, mult_21_C245_n522, mult_21_C245_n521, 
      mult_21_C245_n520, mult_21_C245_n519, mult_21_C245_n518, 
      mult_21_C245_n517, mult_21_C245_n516, mult_21_C245_n515, 
      mult_21_C245_n514, mult_21_C245_n513, mult_21_C245_n512, 
      mult_21_C245_n511, mult_21_C245_n510, mult_21_C245_n509, 
      mult_21_C245_n508, mult_21_C245_n507, mult_21_C245_n506, 
      mult_21_C245_n505, mult_21_C245_n504, mult_21_C245_n503, 
      mult_21_C245_n502, mult_21_C245_n501, mult_21_C245_n500, 
      mult_21_C245_n499, mult_21_C245_n498, mult_21_C245_n497, 
      mult_21_C245_n496, mult_21_C245_n495, mult_21_C245_n494, 
      mult_21_C245_n493, mult_21_C245_n492, mult_21_C245_n491, 
      mult_21_C245_n490, mult_21_C245_n489, mult_21_C245_n488, 
      mult_21_C245_n487, mult_21_C245_n486, mult_21_C245_n485, 
      mult_21_C245_n484, mult_21_C245_n483, mult_21_C245_n482, 
      mult_21_C245_n481, mult_21_C245_n480, mult_21_C245_n479, 
      mult_21_C245_n478, mult_21_C245_n477, mult_21_C245_n476, 
      mult_21_C245_n475, mult_21_C245_n474, mult_21_C245_n473, 
      mult_21_C245_n472, mult_21_C245_n471, mult_21_C245_n470, 
      mult_21_C245_n469, mult_21_C245_n468, mult_21_C245_n467, 
      mult_21_C245_n466, mult_21_C245_n465, mult_21_C245_n464, 
      mult_21_C245_n463, mult_21_C245_n462, mult_21_C245_n461, 
      mult_21_C245_n460, mult_21_C245_n459, mult_21_C245_n458, 
      mult_21_C245_n457, mult_21_C245_n456, mult_21_C245_n455, 
      mult_21_C245_n454, mult_21_C245_n453, mult_21_C245_n452, 
      mult_21_C245_n451, mult_21_C245_n450, mult_21_C245_n449, 
      mult_21_C245_n448, mult_21_C245_n447, mult_21_C245_n446, 
      mult_21_C245_n445, mult_21_C245_n444, mult_21_C245_n443, 
      mult_21_C245_n442, mult_21_C245_n441, mult_21_C245_n440, 
      mult_21_C245_n439, mult_21_C245_n438, mult_21_C245_n437, 
      mult_21_C245_n436, mult_21_C245_n435, mult_21_C245_n434, 
      mult_21_C245_n433, mult_21_C245_n432, mult_21_C245_n431, 
      mult_21_C245_n430, mult_21_C245_n429, mult_21_C245_n428, 
      mult_21_C245_n427, mult_21_C245_n426, mult_21_C245_n425, 
      mult_21_C245_n424, mult_21_C245_n423, mult_21_C245_n422, 
      mult_21_C245_n421, mult_21_C245_n420, mult_21_C245_n419, 
      mult_21_C245_n418, mult_21_C245_n417, mult_21_C245_n416, 
      mult_21_C245_n415, mult_21_C245_n414, mult_21_C245_n413, 
      mult_21_C245_n412, mult_21_C245_n411, mult_21_C245_n410, 
      mult_21_C245_n409, mult_21_C245_n408, mult_21_C245_n407, 
      mult_21_C245_n406, mult_21_C245_n405, mult_21_C245_n404, 
      mult_21_C245_n403, mult_21_C245_n402, mult_21_C245_n401, 
      mult_21_C245_n400, mult_21_C245_n399, mult_21_C245_n398, 
      mult_21_C245_n397, mult_21_C245_n396, mult_21_C245_n395, 
      mult_21_C245_n394, mult_21_C245_n393, mult_21_C245_n392, 
      mult_21_C245_n391, mult_21_C245_n390, mult_21_C245_n389, 
      mult_21_C245_n388, mult_21_C245_n387, mult_21_C245_n386, 
      mult_21_C245_n385, mult_21_C245_n384, mult_21_C245_n383, 
      mult_21_C245_n382, mult_21_C245_n381, mult_21_C245_n380, 
      mult_21_C245_n379, mult_21_C245_n378, mult_21_C245_n377, 
      mult_21_C245_n376, mult_21_C245_n375, mult_21_C245_n374, 
      mult_21_C245_n373, mult_21_C245_n372, mult_21_C245_n371, 
      mult_21_C245_n370, mult_21_C245_n369, mult_21_C245_n368, 
      mult_21_C245_n367, mult_21_C245_n366, mult_21_C245_n365, 
      mult_21_C245_n364, mult_21_C245_n363, mult_21_C245_n362, 
      mult_21_C245_n361, mult_21_C245_n360, mult_21_C245_n359, 
      mult_21_C245_n358, mult_21_C245_n357, mult_21_C245_n356, 
      mult_21_C245_n355, mult_21_C245_n354, mult_21_C245_n353, 
      mult_21_C245_n352, mult_21_C245_n351, mult_21_C245_n350, 
      mult_21_C245_n349, mult_21_C245_n348, mult_21_C245_n347, 
      mult_21_C245_n346, mult_21_C245_n345, mult_21_C245_n344, 
      mult_21_C245_n343, mult_21_C245_n342, mult_21_C245_n341, 
      mult_21_C245_n340, mult_21_C245_n339, mult_21_C245_n338, 
      mult_21_C245_n337, mult_21_C245_n336, mult_21_C245_n335, 
      mult_21_C245_n334, mult_21_C245_n333, mult_21_C245_n332, 
      mult_21_C245_n331, mult_21_C245_n330, mult_21_C245_n329, 
      mult_21_C245_n326, mult_21_C245_n324, mult_21_C245_n323, 
      mult_21_C245_n322, mult_21_C245_n319, mult_21_C245_n318, 
      mult_21_C245_n315, mult_21_C245_n314, mult_21_C245_n313, 
      mult_21_C245_n312, mult_21_C245_n310, mult_21_C245_n305, 
      mult_21_C245_n303, mult_21_C245_n302, mult_21_C245_n301, 
      mult_21_C245_n297, mult_21_C245_n296, mult_21_C245_n295, 
      mult_21_C245_n294, mult_21_C245_n293, mult_21_C245_n289, 
      mult_21_C245_n288, mult_21_C245_n287, mult_21_C245_n286, 
      mult_21_C245_n285, mult_21_C245_n284, mult_21_C245_n283, 
      mult_21_C245_n282, mult_21_C245_n281, mult_21_C245_n280, 
      mult_21_C245_n279, mult_21_C245_n278, mult_21_C245_n277, 
      mult_21_C245_n276, mult_21_C245_n275, mult_21_C245_n273, 
      mult_21_C245_n271, mult_21_C245_n270, mult_21_C245_n268, 
      mult_21_C245_n266, mult_21_C245_n265, mult_21_C245_n264, 
      mult_21_C245_n263, mult_21_C245_n262, mult_21_C245_n261, 
      mult_21_C245_n260, mult_21_C245_n259, mult_21_C245_n258, 
      mult_21_C245_n257, mult_21_C245_n256, mult_21_C245_n255, 
      mult_21_C245_n254, mult_21_C245_n253, mult_21_C245_n251, 
      mult_21_C245_n249, mult_21_C245_n248, mult_21_C245_n246, 
      mult_21_C245_n244, mult_21_C245_n243, mult_21_C245_n242, 
      mult_21_C245_n241, mult_21_C245_n240, mult_21_C245_n239, 
      mult_21_C245_n238, mult_21_C245_n237, mult_21_C245_n236, 
      mult_21_C245_n235, mult_21_C245_n234, mult_21_C245_n233, 
      mult_21_C245_n232, mult_21_C245_n231, mult_21_C245_n230, 
      mult_21_C245_n229, mult_21_C245_n227, mult_21_C245_n226, 
      mult_21_C245_n225, mult_21_C245_n224, mult_21_C245_n223, 
      mult_21_C245_n222, mult_21_C245_n221, mult_21_C245_n219, 
      mult_21_C245_n217, mult_21_C245_n216, mult_21_C245_n215, 
      mult_21_C245_n214, mult_21_C245_n211, mult_21_C245_n209, 
      mult_21_C245_n208, mult_21_C245_n207, mult_21_C245_n206, 
      mult_21_C245_n204, mult_21_C245_n202, mult_21_C245_n201, 
      mult_21_C245_n200, mult_21_C245_n199, mult_21_C245_n197, 
      mult_21_C245_n195, mult_21_C245_n194, mult_21_C245_n190, 
      mult_21_C245_n189, mult_21_C245_n188, mult_21_C245_n187, 
      mult_21_C245_n185, mult_21_C245_n184, mult_21_C245_n183, 
      mult_21_C245_n182, mult_21_C245_n181, mult_21_C245_n180, 
      mult_21_C245_n179, mult_21_C245_n178, mult_21_C245_n176, 
      mult_21_C245_n175, mult_21_C245_n174, mult_21_C245_n173, 
      mult_21_C245_n172, mult_21_C245_n171, mult_21_C245_n170, 
      mult_21_C245_n169, mult_21_C245_n168, mult_21_C245_n167, 
      mult_21_C245_n166, mult_21_C245_n165, mult_21_C245_n164, 
      mult_21_C245_n163, mult_21_C245_n162, mult_21_C245_n161, 
      mult_21_C245_n160, mult_21_C245_n159, mult_21_C245_n158, 
      mult_21_C245_n157, mult_21_C245_n156, mult_21_C245_n155, 
      mult_21_C245_n106, mult_21_C245_n105, mult_21_C245_n104, 
      mult_21_C245_n103, mult_21_C245_n101, mult_21_C245_n99, mult_21_C245_n98,
      mult_21_C245_n96, mult_21_C245_n94, mult_21_C245_n93, mult_21_C245_n91, 
      mult_21_C245_n89, mult_21_C245_n88, mult_21_C245_n86, mult_21_C245_n84, 
      mult_21_C245_n83, mult_21_C245_n81, mult_21_C245_n79, mult_21_C245_n78, 
      mult_21_C245_n76, mult_21_C245_n73, mult_21_C245_n71, mult_21_C245_n69, 
      mult_21_C245_n66, mult_21_C245_n63, mult_21_C245_n61, mult_21_C245_n58, 
      mult_21_C245_n56, mult_21_C245_n53, mult_21_C245_n50, mult_21_C245_n48, 
      mult_21_C245_n45, mult_21_C245_n42, mult_21_C245_n38, mult_21_C245_n30, 
      mult_21_C245_n22, mult_21_C245_n14, mult_21_C245_n8, mult_21_C245_n6, 
      mult_21_C245_n3, mult_21_C247_n1557, mult_21_C247_n1556, 
      mult_21_C247_n1555, mult_21_C247_n1554, mult_21_C247_n1553, 
      mult_21_C247_n1552, mult_21_C247_n1551, mult_21_C247_n1550, 
      mult_21_C247_n1549, mult_21_C247_n1548, mult_21_C247_n1547, 
      mult_21_C247_n1546, mult_21_C247_n1545, mult_21_C247_n1544, 
      mult_21_C247_n1543, mult_21_C247_n1542, mult_21_C247_n1541, 
      mult_21_C247_n1540, mult_21_C247_n1539, mult_21_C247_n1538, 
      mult_21_C247_n1537, mult_21_C247_n1536, mult_21_C247_n1535, 
      mult_21_C247_n1534, mult_21_C247_n1533, mult_21_C247_n1532, 
      mult_21_C247_n1531, mult_21_C247_n1530, mult_21_C247_n1529, 
      mult_21_C247_n1528, mult_21_C247_n1527, mult_21_C247_n1526, 
      mult_21_C247_n1525, mult_21_C247_n1524, mult_21_C247_n1523, 
      mult_21_C247_n1522, mult_21_C247_n1521, mult_21_C247_n1519, 
      mult_21_C247_n1518, mult_21_C247_n1517, mult_21_C247_n1368, 
      mult_21_C247_n1367, mult_21_C247_n1366, mult_21_C247_n1365, 
      mult_21_C247_n1364, mult_21_C247_n1363, mult_21_C247_n1362, 
      mult_21_C247_n1361, mult_21_C247_n1360, mult_21_C247_n1359, 
      mult_21_C247_n1358, mult_21_C247_n1357, mult_21_C247_n1356, 
      mult_21_C247_n1355, mult_21_C247_n1354, mult_21_C247_n1353, 
      mult_21_C247_n1352, mult_21_C247_n1351, mult_21_C247_n1350, 
      mult_21_C247_n1349, mult_21_C247_n1348, mult_21_C247_n1347, 
      mult_21_C247_n1346, mult_21_C247_n1345, mult_21_C247_n1344, 
      mult_21_C247_n1343, mult_21_C247_n1342, mult_21_C247_n1341, 
      mult_21_C247_n1340, mult_21_C247_n1339, mult_21_C247_n1338, 
      mult_21_C247_n1337, mult_21_C247_n1336, mult_21_C247_n1335, 
      mult_21_C247_n1334, mult_21_C247_n1333, mult_21_C247_n1332, 
      mult_21_C247_n1331, mult_21_C247_n1330, mult_21_C247_n1329, 
      mult_21_C247_n1328, mult_21_C247_n1327, mult_21_C247_n1326, 
      mult_21_C247_n1325, mult_21_C247_n1324, mult_21_C247_n1323, 
      mult_21_C247_n1322, mult_21_C247_n1321, mult_21_C247_n1320, 
      mult_21_C247_n1319, mult_21_C247_n1318, mult_21_C247_n1317, 
      mult_21_C247_n1316, mult_21_C247_n1315, mult_21_C247_n1314, 
      mult_21_C247_n1313, mult_21_C247_n1312, mult_21_C247_n1311, 
      mult_21_C247_n1310, mult_21_C247_n1309, mult_21_C247_n1308, 
      mult_21_C247_n1307, mult_21_C247_n1306, mult_21_C247_n1305, 
      mult_21_C247_n1304, mult_21_C247_n1303, mult_21_C247_n1302, 
      mult_21_C247_n1301, mult_21_C247_n1300, mult_21_C247_n1299, 
      mult_21_C247_n1298, mult_21_C247_n1297, mult_21_C247_n1296, 
      mult_21_C247_n1295, mult_21_C247_n1294, mult_21_C247_n1293, 
      mult_21_C247_n1292, mult_21_C247_n1291, mult_21_C247_n1290, 
      mult_21_C247_n1289, mult_21_C247_n1288, mult_21_C247_n1287, 
      mult_21_C247_n1286, mult_21_C247_n1285, mult_21_C247_n1284, 
      mult_21_C247_n1283, mult_21_C247_n1282, mult_21_C247_n1281, 
      mult_21_C247_n1280, mult_21_C247_n1279, mult_21_C247_n1278, 
      mult_21_C247_n1277, mult_21_C247_n1276, mult_21_C247_n1275, 
      mult_21_C247_n1274, mult_21_C247_n1273, mult_21_C247_n1272, 
      mult_21_C247_n1271, mult_21_C247_n1270, mult_21_C247_n1269, 
      mult_21_C247_n1268, mult_21_C247_n1267, mult_21_C247_n1266, 
      mult_21_C247_n1265, mult_21_C247_n1264, mult_21_C247_n1263, 
      mult_21_C247_n1262, mult_21_C247_n1261, mult_21_C247_n1260, 
      mult_21_C247_n1259, mult_21_C247_n1258, mult_21_C247_n1257, 
      mult_21_C247_n1256, mult_21_C247_n1255, mult_21_C247_n1254, 
      mult_21_C247_n1253, mult_21_C247_n1252, mult_21_C247_n1251, 
      mult_21_C247_n1250, mult_21_C247_n1249, mult_21_C247_n1248, 
      mult_21_C247_n1247, mult_21_C247_n1246, mult_21_C247_n1245, 
      mult_21_C247_n1244, mult_21_C247_n1243, mult_21_C247_n1242, 
      mult_21_C247_n1241, mult_21_C247_n1240, mult_21_C247_n1239, 
      mult_21_C247_n1238, mult_21_C247_n1237, mult_21_C247_n1236, 
      mult_21_C247_n1235, mult_21_C247_n1234, mult_21_C247_n1233, 
      mult_21_C247_n1232, mult_21_C247_n1231, mult_21_C247_n1230, 
      mult_21_C247_n1229, mult_21_C247_n1228, mult_21_C247_n1227, 
      mult_21_C247_n1226, mult_21_C247_n1225, mult_21_C247_n1224, 
      mult_21_C247_n1223, mult_21_C247_n1222, mult_21_C247_n1221, 
      mult_21_C247_n1220, mult_21_C247_n1219, mult_21_C247_n1218, 
      mult_21_C247_n1217, mult_21_C247_n1216, mult_21_C247_n1215, 
      mult_21_C247_n1214, mult_21_C247_n1213, mult_21_C247_n1212, 
      mult_21_C247_n1211, mult_21_C247_n1210, mult_21_C247_n1209, 
      mult_21_C247_n1208, mult_21_C247_n1207, mult_21_C247_n1206, 
      mult_21_C247_n1205, mult_21_C247_n1204, mult_21_C247_n1203, 
      mult_21_C247_n1202, mult_21_C247_n1201, mult_21_C247_n1200, 
      mult_21_C247_n1199, mult_21_C247_n1198, mult_21_C247_n1197, 
      mult_21_C247_n1196, mult_21_C247_n1195, mult_21_C247_n1194, 
      mult_21_C247_n1193, mult_21_C247_n1192, mult_21_C247_n1191, 
      mult_21_C247_n1190, mult_21_C247_n1189, mult_21_C247_n1188, 
      mult_21_C247_n1187, mult_21_C247_n1186, mult_21_C247_n1185, 
      mult_21_C247_n1184, mult_21_C247_n1183, mult_21_C247_n1182, 
      mult_21_C247_n1181, mult_21_C247_n1180, mult_21_C247_n1179, 
      mult_21_C247_n1178, mult_21_C247_n1177, mult_21_C247_n1176, 
      mult_21_C247_n1175, mult_21_C247_n1174, mult_21_C247_n1173, 
      mult_21_C247_n1172, mult_21_C247_n1171, mult_21_C247_n1170, 
      mult_21_C247_n1169, mult_21_C247_n1168, mult_21_C247_n1167, 
      mult_21_C247_n1166, mult_21_C247_n1165, mult_21_C247_n1164, 
      mult_21_C247_n1163, mult_21_C247_n1162, mult_21_C247_n1161, 
      mult_21_C247_n1160, mult_21_C247_n1159, mult_21_C247_n1158, 
      mult_21_C247_n1157, mult_21_C247_n1156, mult_21_C247_n1155, 
      mult_21_C247_n1154, mult_21_C247_n1153, mult_21_C247_n1152, 
      mult_21_C247_n1151, mult_21_C247_n1150, mult_21_C247_n1149, 
      mult_21_C247_n1148, mult_21_C247_n1147, mult_21_C247_n1146, 
      mult_21_C247_n1145, mult_21_C247_n1144, mult_21_C247_n1143, 
      mult_21_C247_n1142, mult_21_C247_n1141, mult_21_C247_n1140, 
      mult_21_C247_n1139, mult_21_C247_n1138, mult_21_C247_n1137, 
      mult_21_C247_n1136, mult_21_C247_n1135, mult_21_C247_n1134, 
      mult_21_C247_n1133, mult_21_C247_n1132, mult_21_C247_n1131, 
      mult_21_C247_n1130, mult_21_C247_n1129, mult_21_C247_n1128, 
      mult_21_C247_n1127, mult_21_C247_n1126, mult_21_C247_n1125, 
      mult_21_C247_n1124, mult_21_C247_n1123, mult_21_C247_n1122, 
      mult_21_C247_n1121, mult_21_C247_n1120, mult_21_C247_n1119, 
      mult_21_C247_n1118, mult_21_C247_n1117, mult_21_C247_n1116, 
      mult_21_C247_n1115, mult_21_C247_n1114, mult_21_C247_n1113, 
      mult_21_C247_n1112, mult_21_C247_n1111, mult_21_C247_n1110, 
      mult_21_C247_n1109, mult_21_C247_n1108, mult_21_C247_n1107, 
      mult_21_C247_n1106, mult_21_C247_n1105, mult_21_C247_n1104, 
      mult_21_C247_n1103, mult_21_C247_n1102, mult_21_C247_n1101, 
      mult_21_C247_n1100, mult_21_C247_n1099, mult_21_C247_n1098, 
      mult_21_C247_n1097, mult_21_C247_n1096, mult_21_C247_n1095, 
      mult_21_C247_n1094, mult_21_C247_n1093, mult_21_C247_n1092, 
      mult_21_C247_n1091, mult_21_C247_n1090, mult_21_C247_n1089, 
      mult_21_C247_n1088, mult_21_C247_n1087, mult_21_C247_n1086, 
      mult_21_C247_n1085, mult_21_C247_n1084, mult_21_C247_n1083, 
      mult_21_C247_n1082, mult_21_C247_n1081, mult_21_C247_n1080, 
      mult_21_C247_n1079, mult_21_C247_n1078, mult_21_C247_n1077, 
      mult_21_C247_n1076, mult_21_C247_n1075, mult_21_C247_n1074, 
      mult_21_C247_n1073, mult_21_C247_n1072, mult_21_C247_n1071, 
      mult_21_C247_n1070, mult_21_C247_n1069, mult_21_C247_n1068, 
      mult_21_C247_n1067, mult_21_C247_n1066, mult_21_C247_n1065, 
      mult_21_C247_n1064, mult_21_C247_n1063, mult_21_C247_n1062, 
      mult_21_C247_n1061, mult_21_C247_n1060, mult_21_C247_n1059, 
      mult_21_C247_n1058, mult_21_C247_n1057, mult_21_C247_n1056, 
      mult_21_C247_n1055, mult_21_C247_n1054, mult_21_C247_n1053, 
      mult_21_C247_n1052, mult_21_C247_n1051, mult_21_C247_n1050, 
      mult_21_C247_n1049, mult_21_C247_n1048, mult_21_C247_n1047, 
      mult_21_C247_n1046, mult_21_C247_n1045, mult_21_C247_n1044, 
      mult_21_C247_n1043, mult_21_C247_n1042, mult_21_C247_n1041, 
      mult_21_C247_n1040, mult_21_C247_n1039, mult_21_C247_n1038, 
      mult_21_C247_n1037, mult_21_C247_n1036, mult_21_C247_n1035, 
      mult_21_C247_n1034, mult_21_C247_n1033, mult_21_C247_n1032, 
      mult_21_C247_n1031, mult_21_C247_n1030, mult_21_C247_n1029, 
      mult_21_C247_n1028, mult_21_C247_n1027, mult_21_C247_n1026, 
      mult_21_C247_n1025, mult_21_C247_n1024, mult_21_C247_n1023, 
      mult_21_C247_n1022, mult_21_C247_n1021, mult_21_C247_n1020, 
      mult_21_C247_n1019, mult_21_C247_n1018, mult_21_C247_n1017, 
      mult_21_C247_n1016, mult_21_C247_n1015, mult_21_C247_n1014, 
      mult_21_C247_n1013, mult_21_C247_n1012, mult_21_C247_n1011, 
      mult_21_C247_n1010, mult_21_C247_n1009, mult_21_C247_n1008, 
      mult_21_C247_n1007, mult_21_C247_n1006, mult_21_C247_n1005, 
      mult_21_C247_n1004, mult_21_C247_n1003, mult_21_C247_n1002, 
      mult_21_C247_n1001, mult_21_C247_n1000, mult_21_C247_n999, 
      mult_21_C247_n998, mult_21_C247_n997, mult_21_C247_n996, 
      mult_21_C247_n995, mult_21_C247_n994, mult_21_C247_n993, 
      mult_21_C247_n992, mult_21_C247_n991, mult_21_C247_n990, 
      mult_21_C247_n989, mult_21_C247_n988, mult_21_C247_n987, 
      mult_21_C247_n986, mult_21_C247_n985, mult_21_C247_n984, 
      mult_21_C247_n983, mult_21_C247_n982, mult_21_C247_n981, 
      mult_21_C247_n980, mult_21_C247_n979, mult_21_C247_n978, 
      mult_21_C247_n977, mult_21_C247_n976, mult_21_C247_n975, 
      mult_21_C247_n974, mult_21_C247_n973, mult_21_C247_n972, 
      mult_21_C247_n971, mult_21_C247_n970, mult_21_C247_n969, 
      mult_21_C247_n968, mult_21_C247_n967, mult_21_C247_n966, 
      mult_21_C247_n965, mult_21_C247_n964, mult_21_C247_n963, 
      mult_21_C247_n962, mult_21_C247_n961, mult_21_C247_n960, 
      mult_21_C247_n959, mult_21_C247_n958, mult_21_C247_n957, 
      mult_21_C247_n956, mult_21_C247_n955, mult_21_C247_n954, 
      mult_21_C247_n953, mult_21_C247_n952, mult_21_C247_n951, 
      mult_21_C247_n950, mult_21_C247_n949, mult_21_C247_n948, 
      mult_21_C247_n947, mult_21_C247_n946, mult_21_C247_n945, 
      mult_21_C247_n944, mult_21_C247_n943, mult_21_C247_n942, 
      mult_21_C247_n941, mult_21_C247_n940, mult_21_C247_n939, 
      mult_21_C247_n938, mult_21_C247_n937, mult_21_C247_n936, 
      mult_21_C247_n935, mult_21_C247_n934, mult_21_C247_n933, 
      mult_21_C247_n932, mult_21_C247_n931, mult_21_C247_n930, 
      mult_21_C247_n929, mult_21_C247_n928, mult_21_C247_n927, 
      mult_21_C247_n926, mult_21_C247_n925, mult_21_C247_n924, 
      mult_21_C247_n923, mult_21_C247_n922, mult_21_C247_n921, 
      mult_21_C247_n920, mult_21_C247_n919, mult_21_C247_n918, 
      mult_21_C247_n917, mult_21_C247_n916, mult_21_C247_n915, 
      mult_21_C247_n914, mult_21_C247_n913, mult_21_C247_n912, 
      mult_21_C247_n911, mult_21_C247_n910, mult_21_C247_n909, 
      mult_21_C247_n908, mult_21_C247_n907, mult_21_C247_n906, 
      mult_21_C247_n905, mult_21_C247_n904, mult_21_C247_n903, 
      mult_21_C247_n902, mult_21_C247_n901, mult_21_C247_n900, 
      mult_21_C247_n899, mult_21_C247_n898, mult_21_C247_n897, 
      mult_21_C247_n896, mult_21_C247_n895, mult_21_C247_n894, 
      mult_21_C247_n893, mult_21_C247_n892, mult_21_C247_n891, 
      mult_21_C247_n890, mult_21_C247_n889, mult_21_C247_n888, 
      mult_21_C247_n887, mult_21_C247_n886, mult_21_C247_n885, 
      mult_21_C247_n884, mult_21_C247_n883, mult_21_C247_n882, 
      mult_21_C247_n881, mult_21_C247_n880, mult_21_C247_n879, 
      mult_21_C247_n878, mult_21_C247_n877, mult_21_C247_n876, 
      mult_21_C247_n875, mult_21_C247_n874, mult_21_C247_n873, 
      mult_21_C247_n872, mult_21_C247_n871, mult_21_C247_n870, 
      mult_21_C247_n869, mult_21_C247_n868, mult_21_C247_n867, 
      mult_21_C247_n866, mult_21_C247_n865, mult_21_C247_n864, 
      mult_21_C247_n863, mult_21_C247_n862, mult_21_C247_n861, 
      mult_21_C247_n860, mult_21_C247_n859, mult_21_C247_n858, 
      mult_21_C247_n857, mult_21_C247_n856, mult_21_C247_n855, 
      mult_21_C247_n854, mult_21_C247_n853, mult_21_C247_n852, 
      mult_21_C247_n851, mult_21_C247_n850, mult_21_C247_n849, 
      mult_21_C247_n848, mult_21_C247_n847, mult_21_C247_n846, 
      mult_21_C247_n845, mult_21_C247_n844, mult_21_C247_n843, 
      mult_21_C247_n842, mult_21_C247_n841, mult_21_C247_n840, 
      mult_21_C247_n839, mult_21_C247_n838, mult_21_C247_n837, 
      mult_21_C247_n836, mult_21_C247_n835, mult_21_C247_n834, 
      mult_21_C247_n833, mult_21_C247_n832, mult_21_C247_n831, 
      mult_21_C247_n830, mult_21_C247_n829, mult_21_C247_n828, 
      mult_21_C247_n827, mult_21_C247_n826, mult_21_C247_n825, 
      mult_21_C247_n824, mult_21_C247_n823, mult_21_C247_n822, 
      mult_21_C247_n821, mult_21_C247_n820, mult_21_C247_n819, 
      mult_21_C247_n818, mult_21_C247_n817, mult_21_C247_n816, 
      mult_21_C247_n815, mult_21_C247_n814, mult_21_C247_n813, 
      mult_21_C247_n812, mult_21_C247_n811, mult_21_C247_n810, 
      mult_21_C247_n809, mult_21_C247_n808, mult_21_C247_n807, 
      mult_21_C247_n806, mult_21_C247_n805, mult_21_C247_n804, 
      mult_21_C247_n803, mult_21_C247_n802, mult_21_C247_n801, 
      mult_21_C247_n800, mult_21_C247_n799, mult_21_C247_n798, 
      mult_21_C247_n797, mult_21_C247_n796, mult_21_C247_n795, 
      mult_21_C247_n794, mult_21_C247_n793, mult_21_C247_n792, 
      mult_21_C247_n791, mult_21_C247_n790, mult_21_C247_n789, 
      mult_21_C247_n788, mult_21_C247_n787, mult_21_C247_n786, 
      mult_21_C247_n785, mult_21_C247_n784, mult_21_C247_n783, 
      mult_21_C247_n782, mult_21_C247_n781, mult_21_C247_n780, 
      mult_21_C247_n779, mult_21_C247_n778, mult_21_C247_n777, 
      mult_21_C247_n776, mult_21_C247_n775, mult_21_C247_n774, 
      mult_21_C247_n773, mult_21_C247_n772, mult_21_C247_n771, 
      mult_21_C247_n770, mult_21_C247_n769, mult_21_C247_n768, 
      mult_21_C247_n767, mult_21_C247_n766, mult_21_C247_n765, 
      mult_21_C247_n764, mult_21_C247_n763, mult_21_C247_n762, 
      mult_21_C247_n761, mult_21_C247_n760, mult_21_C247_n759, 
      mult_21_C247_n758, mult_21_C247_n757, mult_21_C247_n756, 
      mult_21_C247_n755, mult_21_C247_n754, mult_21_C247_n753, 
      mult_21_C247_n752, mult_21_C247_n751, mult_21_C247_n750, 
      mult_21_C247_n749, mult_21_C247_n748, mult_21_C247_n747, 
      mult_21_C247_n746, mult_21_C247_n745, mult_21_C247_n744, 
      mult_21_C247_n743, mult_21_C247_n742, mult_21_C247_n741, 
      mult_21_C247_n740, mult_21_C247_n739, mult_21_C247_n738, 
      mult_21_C247_n737, mult_21_C247_n736, mult_21_C247_n735, 
      mult_21_C247_n734, mult_21_C247_n733, mult_21_C247_n732, 
      mult_21_C247_n731, mult_21_C247_n730, mult_21_C247_n729, 
      mult_21_C247_n728, mult_21_C247_n727, mult_21_C247_n726, 
      mult_21_C247_n725, mult_21_C247_n724, mult_21_C247_n723, 
      mult_21_C247_n722, mult_21_C247_n721, mult_21_C247_n720, 
      mult_21_C247_n719, mult_21_C247_n718, mult_21_C247_n717, 
      mult_21_C247_n716, mult_21_C247_n715, mult_21_C247_n714, 
      mult_21_C247_n713, mult_21_C247_n712, mult_21_C247_n711, 
      mult_21_C247_n710, mult_21_C247_n709, mult_21_C247_n708, 
      mult_21_C247_n707, mult_21_C247_n706, mult_21_C247_n705, 
      mult_21_C247_n704, mult_21_C247_n703, mult_21_C247_n702, 
      mult_21_C247_n701, mult_21_C247_n700, mult_21_C247_n699, 
      mult_21_C247_n698, mult_21_C247_n697, mult_21_C247_n696, 
      mult_21_C247_n695, mult_21_C247_n694, mult_21_C247_n693, 
      mult_21_C247_n692, mult_21_C247_n691, mult_21_C247_n690, 
      mult_21_C247_n689, mult_21_C247_n688, mult_21_C247_n687, 
      mult_21_C247_n686, mult_21_C247_n685, mult_21_C247_n684, 
      mult_21_C247_n683, mult_21_C247_n682, mult_21_C247_n681, 
      mult_21_C247_n680, mult_21_C247_n679, mult_21_C247_n678, 
      mult_21_C247_n677, mult_21_C247_n676, mult_21_C247_n675, 
      mult_21_C247_n674, mult_21_C247_n673, mult_21_C247_n672, 
      mult_21_C247_n671, mult_21_C247_n670, mult_21_C247_n669, 
      mult_21_C247_n668, mult_21_C247_n667, mult_21_C247_n666, 
      mult_21_C247_n665, mult_21_C247_n664, mult_21_C247_n663, 
      mult_21_C247_n662, mult_21_C247_n661, mult_21_C247_n660, 
      mult_21_C247_n659, mult_21_C247_n658, mult_21_C247_n657, 
      mult_21_C247_n656, mult_21_C247_n655, mult_21_C247_n654, 
      mult_21_C247_n653, mult_21_C247_n652, mult_21_C247_n651, 
      mult_21_C247_n650, mult_21_C247_n649, mult_21_C247_n648, 
      mult_21_C247_n647, mult_21_C247_n646, mult_21_C247_n645, 
      mult_21_C247_n644, mult_21_C247_n643, mult_21_C247_n642, 
      mult_21_C247_n641, mult_21_C247_n640, mult_21_C247_n639, 
      mult_21_C247_n638, mult_21_C247_n637, mult_21_C247_n636, 
      mult_21_C247_n635, mult_21_C247_n634, mult_21_C247_n633, 
      mult_21_C247_n632, mult_21_C247_n631, mult_21_C247_n630, 
      mult_21_C247_n629, mult_21_C247_n628, mult_21_C247_n627, 
      mult_21_C247_n626, mult_21_C247_n625, mult_21_C247_n624, 
      mult_21_C247_n623, mult_21_C247_n622, mult_21_C247_n621, 
      mult_21_C247_n620, mult_21_C247_n619, mult_21_C247_n618, 
      mult_21_C247_n617, mult_21_C247_n616, mult_21_C247_n615, 
      mult_21_C247_n614, mult_21_C247_n613, mult_21_C247_n612, 
      mult_21_C247_n611, mult_21_C247_n610, mult_21_C247_n609, 
      mult_21_C247_n608, mult_21_C247_n607, mult_21_C247_n606, 
      mult_21_C247_n605, mult_21_C247_n604, mult_21_C247_n603, 
      mult_21_C247_n602, mult_21_C247_n601, mult_21_C247_n600, 
      mult_21_C247_n599, mult_21_C247_n598, mult_21_C247_n597, 
      mult_21_C247_n596, mult_21_C247_n595, mult_21_C247_n594, 
      mult_21_C247_n593, mult_21_C247_n592, mult_21_C247_n591, 
      mult_21_C247_n590, mult_21_C247_n589, mult_21_C247_n588, 
      mult_21_C247_n587, mult_21_C247_n586, mult_21_C247_n585, 
      mult_21_C247_n584, mult_21_C247_n583, mult_21_C247_n582, 
      mult_21_C247_n581, mult_21_C247_n580, mult_21_C247_n579, 
      mult_21_C247_n578, mult_21_C247_n577, mult_21_C247_n576, 
      mult_21_C247_n575, mult_21_C247_n574, mult_21_C247_n573, 
      mult_21_C247_n572, mult_21_C247_n571, mult_21_C247_n570, 
      mult_21_C247_n569, mult_21_C247_n568, mult_21_C247_n567, 
      mult_21_C247_n566, mult_21_C247_n565, mult_21_C247_n564, 
      mult_21_C247_n563, mult_21_C247_n562, mult_21_C247_n561, 
      mult_21_C247_n560, mult_21_C247_n559, mult_21_C247_n558, 
      mult_21_C247_n557, mult_21_C247_n556, mult_21_C247_n555, 
      mult_21_C247_n554, mult_21_C247_n553, mult_21_C247_n552, 
      mult_21_C247_n551, mult_21_C247_n550, mult_21_C247_n549, 
      mult_21_C247_n548, mult_21_C247_n547, mult_21_C247_n546, 
      mult_21_C247_n545, mult_21_C247_n544, mult_21_C247_n543, 
      mult_21_C247_n542, mult_21_C247_n541, mult_21_C247_n540, 
      mult_21_C247_n539, mult_21_C247_n538, mult_21_C247_n537, 
      mult_21_C247_n536, mult_21_C247_n535, mult_21_C247_n534, 
      mult_21_C247_n533, mult_21_C247_n532, mult_21_C247_n531, 
      mult_21_C247_n530, mult_21_C247_n529, mult_21_C247_n528, 
      mult_21_C247_n527, mult_21_C247_n526, mult_21_C247_n525, 
      mult_21_C247_n524, mult_21_C247_n523, mult_21_C247_n522, 
      mult_21_C247_n521, mult_21_C247_n520, mult_21_C247_n519, 
      mult_21_C247_n518, mult_21_C247_n517, mult_21_C247_n516, 
      mult_21_C247_n515, mult_21_C247_n514, mult_21_C247_n513, 
      mult_21_C247_n512, mult_21_C247_n511, mult_21_C247_n510, 
      mult_21_C247_n509, mult_21_C247_n508, mult_21_C247_n507, 
      mult_21_C247_n506, mult_21_C247_n505, mult_21_C247_n504, 
      mult_21_C247_n503, mult_21_C247_n502, mult_21_C247_n501, 
      mult_21_C247_n500, mult_21_C247_n499, mult_21_C247_n498, 
      mult_21_C247_n497, mult_21_C247_n496, mult_21_C247_n495, 
      mult_21_C247_n494, mult_21_C247_n493, mult_21_C247_n492, 
      mult_21_C247_n491, mult_21_C247_n490, mult_21_C247_n489, 
      mult_21_C247_n488, mult_21_C247_n487, mult_21_C247_n486, 
      mult_21_C247_n485, mult_21_C247_n484, mult_21_C247_n483, 
      mult_21_C247_n482, mult_21_C247_n481, mult_21_C247_n480, 
      mult_21_C247_n479, mult_21_C247_n478, mult_21_C247_n477, 
      mult_21_C247_n476, mult_21_C247_n475, mult_21_C247_n474, 
      mult_21_C247_n473, mult_21_C247_n472, mult_21_C247_n471, 
      mult_21_C247_n470, mult_21_C247_n469, mult_21_C247_n468, 
      mult_21_C247_n467, mult_21_C247_n466, mult_21_C247_n465, 
      mult_21_C247_n464, mult_21_C247_n463, mult_21_C247_n462, 
      mult_21_C247_n461, mult_21_C247_n460, mult_21_C247_n459, 
      mult_21_C247_n458, mult_21_C247_n457, mult_21_C247_n456, 
      mult_21_C247_n455, mult_21_C247_n454, mult_21_C247_n453, 
      mult_21_C247_n452, mult_21_C247_n451, mult_21_C247_n450, 
      mult_21_C247_n449, mult_21_C247_n448, mult_21_C247_n447, 
      mult_21_C247_n446, mult_21_C247_n445, mult_21_C247_n444, 
      mult_21_C247_n443, mult_21_C247_n442, mult_21_C247_n441, 
      mult_21_C247_n440, mult_21_C247_n439, mult_21_C247_n438, 
      mult_21_C247_n437, mult_21_C247_n436, mult_21_C247_n435, 
      mult_21_C247_n434, mult_21_C247_n433, mult_21_C247_n432, 
      mult_21_C247_n431, mult_21_C247_n430, mult_21_C247_n429, 
      mult_21_C247_n428, mult_21_C247_n427, mult_21_C247_n426, 
      mult_21_C247_n425, mult_21_C247_n424, mult_21_C247_n423, 
      mult_21_C247_n422, mult_21_C247_n421, mult_21_C247_n420, 
      mult_21_C247_n419, mult_21_C247_n418, mult_21_C247_n417, 
      mult_21_C247_n416, mult_21_C247_n415, mult_21_C247_n414, 
      mult_21_C247_n413, mult_21_C247_n412, mult_21_C247_n411, 
      mult_21_C247_n410, mult_21_C247_n409, mult_21_C247_n408, 
      mult_21_C247_n407, mult_21_C247_n406, mult_21_C247_n405, 
      mult_21_C247_n404, mult_21_C247_n403, mult_21_C247_n402, 
      mult_21_C247_n401, mult_21_C247_n400, mult_21_C247_n399, 
      mult_21_C247_n398, mult_21_C247_n397, mult_21_C247_n396, 
      mult_21_C247_n395, mult_21_C247_n394, mult_21_C247_n393, 
      mult_21_C247_n392, mult_21_C247_n391, mult_21_C247_n390, 
      mult_21_C247_n389, mult_21_C247_n388, mult_21_C247_n387, 
      mult_21_C247_n386, mult_21_C247_n385, mult_21_C247_n384, 
      mult_21_C247_n383, mult_21_C247_n382, mult_21_C247_n381, 
      mult_21_C247_n380, mult_21_C247_n379, mult_21_C247_n378, 
      mult_21_C247_n377, mult_21_C247_n376, mult_21_C247_n375, 
      mult_21_C247_n374, mult_21_C247_n373, mult_21_C247_n372, 
      mult_21_C247_n371, mult_21_C247_n370, mult_21_C247_n369, 
      mult_21_C247_n368, mult_21_C247_n367, mult_21_C247_n366, 
      mult_21_C247_n365, mult_21_C247_n364, mult_21_C247_n363, 
      mult_21_C247_n362, mult_21_C247_n361, mult_21_C247_n360, 
      mult_21_C247_n359, mult_21_C247_n358, mult_21_C247_n357, 
      mult_21_C247_n356, mult_21_C247_n355, mult_21_C247_n354, 
      mult_21_C247_n353, mult_21_C247_n352, mult_21_C247_n351, 
      mult_21_C247_n350, mult_21_C247_n349, mult_21_C247_n348, 
      mult_21_C247_n347, mult_21_C247_n346, mult_21_C247_n345, 
      mult_21_C247_n344, mult_21_C247_n343, mult_21_C247_n342, 
      mult_21_C247_n341, mult_21_C247_n340, mult_21_C247_n339, 
      mult_21_C247_n338, mult_21_C247_n337, mult_21_C247_n336, 
      mult_21_C247_n335, mult_21_C247_n334, mult_21_C247_n333, 
      mult_21_C247_n332, mult_21_C247_n331, mult_21_C247_n330, 
      mult_21_C247_n329, mult_21_C247_n326, mult_21_C247_n324, 
      mult_21_C247_n323, mult_21_C247_n322, mult_21_C247_n319, 
      mult_21_C247_n318, mult_21_C247_n315, mult_21_C247_n314, 
      mult_21_C247_n313, mult_21_C247_n312, mult_21_C247_n310, 
      mult_21_C247_n305, mult_21_C247_n303, mult_21_C247_n302, 
      mult_21_C247_n301, mult_21_C247_n297, mult_21_C247_n296, 
      mult_21_C247_n295, mult_21_C247_n294, mult_21_C247_n293, 
      mult_21_C247_n289, mult_21_C247_n288, mult_21_C247_n287, 
      mult_21_C247_n286, mult_21_C247_n285, mult_21_C247_n284, 
      mult_21_C247_n283, mult_21_C247_n282, mult_21_C247_n281, 
      mult_21_C247_n280, mult_21_C247_n279, mult_21_C247_n278, 
      mult_21_C247_n277, mult_21_C247_n276, mult_21_C247_n275, 
      mult_21_C247_n273, mult_21_C247_n271, mult_21_C247_n270, 
      mult_21_C247_n268, mult_21_C247_n266, mult_21_C247_n265, 
      mult_21_C247_n264, mult_21_C247_n263, mult_21_C247_n262, 
      mult_21_C247_n261, mult_21_C247_n260, mult_21_C247_n259, 
      mult_21_C247_n258, mult_21_C247_n257, mult_21_C247_n256, 
      mult_21_C247_n255, mult_21_C247_n254, mult_21_C247_n253, 
      mult_21_C247_n251, mult_21_C247_n249, mult_21_C247_n248, 
      mult_21_C247_n246, mult_21_C247_n244, mult_21_C247_n243, 
      mult_21_C247_n242, mult_21_C247_n241, mult_21_C247_n240, 
      mult_21_C247_n239, mult_21_C247_n238, mult_21_C247_n237, 
      mult_21_C247_n236, mult_21_C247_n235, mult_21_C247_n234, 
      mult_21_C247_n233, mult_21_C247_n232, mult_21_C247_n231, 
      mult_21_C247_n230, mult_21_C247_n229, mult_21_C247_n227, 
      mult_21_C247_n226, mult_21_C247_n225, mult_21_C247_n224, 
      mult_21_C247_n223, mult_21_C247_n222, mult_21_C247_n221, 
      mult_21_C247_n219, mult_21_C247_n217, mult_21_C247_n216, 
      mult_21_C247_n215, mult_21_C247_n214, mult_21_C247_n211, 
      mult_21_C247_n209, mult_21_C247_n208, mult_21_C247_n207, 
      mult_21_C247_n206, mult_21_C247_n204, mult_21_C247_n202, 
      mult_21_C247_n201, mult_21_C247_n200, mult_21_C247_n199, 
      mult_21_C247_n197, mult_21_C247_n195, mult_21_C247_n194, 
      mult_21_C247_n190, mult_21_C247_n189, mult_21_C247_n188, 
      mult_21_C247_n187, mult_21_C247_n185, mult_21_C247_n184, 
      mult_21_C247_n183, mult_21_C247_n182, mult_21_C247_n181, 
      mult_21_C247_n180, mult_21_C247_n179, mult_21_C247_n178, 
      mult_21_C247_n176, mult_21_C247_n175, mult_21_C247_n174, 
      mult_21_C247_n173, mult_21_C247_n172, mult_21_C247_n171, 
      mult_21_C247_n170, mult_21_C247_n169, mult_21_C247_n168, 
      mult_21_C247_n167, mult_21_C247_n166, mult_21_C247_n165, 
      mult_21_C247_n164, mult_21_C247_n163, mult_21_C247_n162, 
      mult_21_C247_n161, mult_21_C247_n160, mult_21_C247_n159, 
      mult_21_C247_n158, mult_21_C247_n157, mult_21_C247_n156, 
      mult_21_C247_n155, mult_21_C247_n106, mult_21_C247_n105, 
      mult_21_C247_n104, mult_21_C247_n103, mult_21_C247_n101, mult_21_C247_n99
      , mult_21_C247_n98, mult_21_C247_n96, mult_21_C247_n94, mult_21_C247_n93,
      mult_21_C247_n91, mult_21_C247_n89, mult_21_C247_n88, mult_21_C247_n86, 
      mult_21_C247_n84, mult_21_C247_n83, mult_21_C247_n81, mult_21_C247_n79, 
      mult_21_C247_n78, mult_21_C247_n76, mult_21_C247_n73, mult_21_C247_n71, 
      mult_21_C247_n69, mult_21_C247_n66, mult_21_C247_n63, mult_21_C247_n61, 
      mult_21_C247_n58, mult_21_C247_n56, mult_21_C247_n53, mult_21_C247_n50, 
      mult_21_C247_n48, mult_21_C247_n45, mult_21_C247_n42, mult_21_C247_n38, 
      mult_21_C247_n30, mult_21_C247_n22, mult_21_C247_n14, mult_21_C247_n8, 
      mult_21_C247_n6, mult_21_C247_n3, mult_21_C249_n1557, mult_21_C249_n1556,
      mult_21_C249_n1555, mult_21_C249_n1554, mult_21_C249_n1553, 
      mult_21_C249_n1552, mult_21_C249_n1551, mult_21_C249_n1550, 
      mult_21_C249_n1549, mult_21_C249_n1548, mult_21_C249_n1547, 
      mult_21_C249_n1546, mult_21_C249_n1545, mult_21_C249_n1544, 
      mult_21_C249_n1543, mult_21_C249_n1542, mult_21_C249_n1541, 
      mult_21_C249_n1540, mult_21_C249_n1539, mult_21_C249_n1538, 
      mult_21_C249_n1537, mult_21_C249_n1536, mult_21_C249_n1535, 
      mult_21_C249_n1534, mult_21_C249_n1533, mult_21_C249_n1532, 
      mult_21_C249_n1531, mult_21_C249_n1530, mult_21_C249_n1529, 
      mult_21_C249_n1528, mult_21_C249_n1527, mult_21_C249_n1526, 
      mult_21_C249_n1525, mult_21_C249_n1524, mult_21_C249_n1523, 
      mult_21_C249_n1521, mult_21_C249_n1520, mult_21_C249_n1519, 
      mult_21_C249_n1518, mult_21_C249_n1517, mult_21_C249_n1368, 
      mult_21_C249_n1367, mult_21_C249_n1366, mult_21_C249_n1365, 
      mult_21_C249_n1364, mult_21_C249_n1363, mult_21_C249_n1362, 
      mult_21_C249_n1361, mult_21_C249_n1360, mult_21_C249_n1359, 
      mult_21_C249_n1358, mult_21_C249_n1357, mult_21_C249_n1356, 
      mult_21_C249_n1355, mult_21_C249_n1354, mult_21_C249_n1353, 
      mult_21_C249_n1352, mult_21_C249_n1351, mult_21_C249_n1350, 
      mult_21_C249_n1349, mult_21_C249_n1348, mult_21_C249_n1347, 
      mult_21_C249_n1346, mult_21_C249_n1345, mult_21_C249_n1344, 
      mult_21_C249_n1343, mult_21_C249_n1342, mult_21_C249_n1341, 
      mult_21_C249_n1340, mult_21_C249_n1339, mult_21_C249_n1338, 
      mult_21_C249_n1337, mult_21_C249_n1336, mult_21_C249_n1335, 
      mult_21_C249_n1334, mult_21_C249_n1333, mult_21_C249_n1332, 
      mult_21_C249_n1331, mult_21_C249_n1330, mult_21_C249_n1329, 
      mult_21_C249_n1328, mult_21_C249_n1327, mult_21_C249_n1326, 
      mult_21_C249_n1325, mult_21_C249_n1324, mult_21_C249_n1323, 
      mult_21_C249_n1322, mult_21_C249_n1321, mult_21_C249_n1320, 
      mult_21_C249_n1319, mult_21_C249_n1318, mult_21_C249_n1317, 
      mult_21_C249_n1316, mult_21_C249_n1315, mult_21_C249_n1314, 
      mult_21_C249_n1313, mult_21_C249_n1312, mult_21_C249_n1311, 
      mult_21_C249_n1310, mult_21_C249_n1309, mult_21_C249_n1308, 
      mult_21_C249_n1307, mult_21_C249_n1306, mult_21_C249_n1305, 
      mult_21_C249_n1304, mult_21_C249_n1303, mult_21_C249_n1302, 
      mult_21_C249_n1301, mult_21_C249_n1300, mult_21_C249_n1299, 
      mult_21_C249_n1298, mult_21_C249_n1297, mult_21_C249_n1296, 
      mult_21_C249_n1295, mult_21_C249_n1294, mult_21_C249_n1293, 
      mult_21_C249_n1292, mult_21_C249_n1291, mult_21_C249_n1290, 
      mult_21_C249_n1289, mult_21_C249_n1288, mult_21_C249_n1287, 
      mult_21_C249_n1286, mult_21_C249_n1285, mult_21_C249_n1284, 
      mult_21_C249_n1283, mult_21_C249_n1282, mult_21_C249_n1281, 
      mult_21_C249_n1280, mult_21_C249_n1279, mult_21_C249_n1278, 
      mult_21_C249_n1277, mult_21_C249_n1276, mult_21_C249_n1275, 
      mult_21_C249_n1274, mult_21_C249_n1273, mult_21_C249_n1272, 
      mult_21_C249_n1271, mult_21_C249_n1270, mult_21_C249_n1269, 
      mult_21_C249_n1268, mult_21_C249_n1267, mult_21_C249_n1266, 
      mult_21_C249_n1265, mult_21_C249_n1264, mult_21_C249_n1263, 
      mult_21_C249_n1262, mult_21_C249_n1261, mult_21_C249_n1260, 
      mult_21_C249_n1259, mult_21_C249_n1258, mult_21_C249_n1257, 
      mult_21_C249_n1256, mult_21_C249_n1255, mult_21_C249_n1254, 
      mult_21_C249_n1253, mult_21_C249_n1252, mult_21_C249_n1251, 
      mult_21_C249_n1250, mult_21_C249_n1249, mult_21_C249_n1248, 
      mult_21_C249_n1247, mult_21_C249_n1246, mult_21_C249_n1245, 
      mult_21_C249_n1244, mult_21_C249_n1243, mult_21_C249_n1242, 
      mult_21_C249_n1241, mult_21_C249_n1240, mult_21_C249_n1239, 
      mult_21_C249_n1238, mult_21_C249_n1237, mult_21_C249_n1236, 
      mult_21_C249_n1235, mult_21_C249_n1234, mult_21_C249_n1233, 
      mult_21_C249_n1232, mult_21_C249_n1231, mult_21_C249_n1230, 
      mult_21_C249_n1229, mult_21_C249_n1228, mult_21_C249_n1227, 
      mult_21_C249_n1226, mult_21_C249_n1225, mult_21_C249_n1224, 
      mult_21_C249_n1223, mult_21_C249_n1222, mult_21_C249_n1221, 
      mult_21_C249_n1220, mult_21_C249_n1219, mult_21_C249_n1218, 
      mult_21_C249_n1217, mult_21_C249_n1216, mult_21_C249_n1215, 
      mult_21_C249_n1214, mult_21_C249_n1213, mult_21_C249_n1212, 
      mult_21_C249_n1211, mult_21_C249_n1210, mult_21_C249_n1209, 
      mult_21_C249_n1208, mult_21_C249_n1207, mult_21_C249_n1206, 
      mult_21_C249_n1205, mult_21_C249_n1204, mult_21_C249_n1203, 
      mult_21_C249_n1202, mult_21_C249_n1201, mult_21_C249_n1200, 
      mult_21_C249_n1199, mult_21_C249_n1198, mult_21_C249_n1197, 
      mult_21_C249_n1196, mult_21_C249_n1195, mult_21_C249_n1194, 
      mult_21_C249_n1193, mult_21_C249_n1192, mult_21_C249_n1191, 
      mult_21_C249_n1190, mult_21_C249_n1189, mult_21_C249_n1188, 
      mult_21_C249_n1187, mult_21_C249_n1186, mult_21_C249_n1185, 
      mult_21_C249_n1184, mult_21_C249_n1183, mult_21_C249_n1182, 
      mult_21_C249_n1181, mult_21_C249_n1180, mult_21_C249_n1179, 
      mult_21_C249_n1178, mult_21_C249_n1177, mult_21_C249_n1176, 
      mult_21_C249_n1175, mult_21_C249_n1174, mult_21_C249_n1173, 
      mult_21_C249_n1172, mult_21_C249_n1171, mult_21_C249_n1170, 
      mult_21_C249_n1169, mult_21_C249_n1168, mult_21_C249_n1167, 
      mult_21_C249_n1166, mult_21_C249_n1165, mult_21_C249_n1164, 
      mult_21_C249_n1163, mult_21_C249_n1162, mult_21_C249_n1161, 
      mult_21_C249_n1160, mult_21_C249_n1159, mult_21_C249_n1158, 
      mult_21_C249_n1157, mult_21_C249_n1156, mult_21_C249_n1155, 
      mult_21_C249_n1154, mult_21_C249_n1153, mult_21_C249_n1152, 
      mult_21_C249_n1151, mult_21_C249_n1150, mult_21_C249_n1149, 
      mult_21_C249_n1148, mult_21_C249_n1147, mult_21_C249_n1146, 
      mult_21_C249_n1145, mult_21_C249_n1144, mult_21_C249_n1143, 
      mult_21_C249_n1142, mult_21_C249_n1141, mult_21_C249_n1140, 
      mult_21_C249_n1139, mult_21_C249_n1138, mult_21_C249_n1137, 
      mult_21_C249_n1136, mult_21_C249_n1135, mult_21_C249_n1134, 
      mult_21_C249_n1133, mult_21_C249_n1132, mult_21_C249_n1131, 
      mult_21_C249_n1130, mult_21_C249_n1129, mult_21_C249_n1128, 
      mult_21_C249_n1127, mult_21_C249_n1126, mult_21_C249_n1125, 
      mult_21_C249_n1124, mult_21_C249_n1123, mult_21_C249_n1122, 
      mult_21_C249_n1121, mult_21_C249_n1120, mult_21_C249_n1119, 
      mult_21_C249_n1118, mult_21_C249_n1117, mult_21_C249_n1116, 
      mult_21_C249_n1115, mult_21_C249_n1114, mult_21_C249_n1113, 
      mult_21_C249_n1112, mult_21_C249_n1111, mult_21_C249_n1110, 
      mult_21_C249_n1109, mult_21_C249_n1108, mult_21_C249_n1107, 
      mult_21_C249_n1106, mult_21_C249_n1105, mult_21_C249_n1104, 
      mult_21_C249_n1103, mult_21_C249_n1102, mult_21_C249_n1101, 
      mult_21_C249_n1100, mult_21_C249_n1099, mult_21_C249_n1098, 
      mult_21_C249_n1097, mult_21_C249_n1096, mult_21_C249_n1095, 
      mult_21_C249_n1094, mult_21_C249_n1093, mult_21_C249_n1092, 
      mult_21_C249_n1091, mult_21_C249_n1090, mult_21_C249_n1089, 
      mult_21_C249_n1088, mult_21_C249_n1087, mult_21_C249_n1086, 
      mult_21_C249_n1085, mult_21_C249_n1084, mult_21_C249_n1083, 
      mult_21_C249_n1082, mult_21_C249_n1081, mult_21_C249_n1080, 
      mult_21_C249_n1079, mult_21_C249_n1078, mult_21_C249_n1077, 
      mult_21_C249_n1076, mult_21_C249_n1075, mult_21_C249_n1074, 
      mult_21_C249_n1073, mult_21_C249_n1072, mult_21_C249_n1071, 
      mult_21_C249_n1070, mult_21_C249_n1069, mult_21_C249_n1068, 
      mult_21_C249_n1067, mult_21_C249_n1066, mult_21_C249_n1065, 
      mult_21_C249_n1064, mult_21_C249_n1063, mult_21_C249_n1062, 
      mult_21_C249_n1061, mult_21_C249_n1060, mult_21_C249_n1059, 
      mult_21_C249_n1058, mult_21_C249_n1057, mult_21_C249_n1056, 
      mult_21_C249_n1055, mult_21_C249_n1054, mult_21_C249_n1053, 
      mult_21_C249_n1052, mult_21_C249_n1051, mult_21_C249_n1050, 
      mult_21_C249_n1049, mult_21_C249_n1048, mult_21_C249_n1047, 
      mult_21_C249_n1046, mult_21_C249_n1045, mult_21_C249_n1044, 
      mult_21_C249_n1043, mult_21_C249_n1042, mult_21_C249_n1041, 
      mult_21_C249_n1040, mult_21_C249_n1039, mult_21_C249_n1038, 
      mult_21_C249_n1037, mult_21_C249_n1036, mult_21_C249_n1035, 
      mult_21_C249_n1034, mult_21_C249_n1033, mult_21_C249_n1032, 
      mult_21_C249_n1031, mult_21_C249_n1030, mult_21_C249_n1029, 
      mult_21_C249_n1028, mult_21_C249_n1027, mult_21_C249_n1026, 
      mult_21_C249_n1025, mult_21_C249_n1024, mult_21_C249_n1023, 
      mult_21_C249_n1022, mult_21_C249_n1021, mult_21_C249_n1020, 
      mult_21_C249_n1019, mult_21_C249_n1018, mult_21_C249_n1017, 
      mult_21_C249_n1016, mult_21_C249_n1015, mult_21_C249_n1014, 
      mult_21_C249_n1013, mult_21_C249_n1012, mult_21_C249_n1011, 
      mult_21_C249_n1010, mult_21_C249_n1009, mult_21_C249_n1008, 
      mult_21_C249_n1007, mult_21_C249_n1006, mult_21_C249_n1005, 
      mult_21_C249_n1004, mult_21_C249_n1003, mult_21_C249_n1002, 
      mult_21_C249_n1001, mult_21_C249_n1000, mult_21_C249_n999, 
      mult_21_C249_n998, mult_21_C249_n997, mult_21_C249_n996, 
      mult_21_C249_n995, mult_21_C249_n994, mult_21_C249_n993, 
      mult_21_C249_n992, mult_21_C249_n991, mult_21_C249_n990, 
      mult_21_C249_n989, mult_21_C249_n988, mult_21_C249_n987, 
      mult_21_C249_n986, mult_21_C249_n985, mult_21_C249_n984, 
      mult_21_C249_n983, mult_21_C249_n982, mult_21_C249_n981, 
      mult_21_C249_n980, mult_21_C249_n979, mult_21_C249_n978, 
      mult_21_C249_n977, mult_21_C249_n976, mult_21_C249_n975, 
      mult_21_C249_n974, mult_21_C249_n973, mult_21_C249_n972, 
      mult_21_C249_n971, mult_21_C249_n970, mult_21_C249_n969, 
      mult_21_C249_n968, mult_21_C249_n967, mult_21_C249_n966, 
      mult_21_C249_n965, mult_21_C249_n964, mult_21_C249_n963, 
      mult_21_C249_n962, mult_21_C249_n961, mult_21_C249_n960, 
      mult_21_C249_n959, mult_21_C249_n958, mult_21_C249_n957, 
      mult_21_C249_n956, mult_21_C249_n955, mult_21_C249_n954, 
      mult_21_C249_n953, mult_21_C249_n952, mult_21_C249_n951, 
      mult_21_C249_n950, mult_21_C249_n949, mult_21_C249_n948, 
      mult_21_C249_n947, mult_21_C249_n946, mult_21_C249_n945, 
      mult_21_C249_n944, mult_21_C249_n943, mult_21_C249_n942, 
      mult_21_C249_n941, mult_21_C249_n940, mult_21_C249_n939, 
      mult_21_C249_n938, mult_21_C249_n937, mult_21_C249_n936, 
      mult_21_C249_n935, mult_21_C249_n934, mult_21_C249_n933, 
      mult_21_C249_n932, mult_21_C249_n931, mult_21_C249_n930, 
      mult_21_C249_n929, mult_21_C249_n928, mult_21_C249_n927, 
      mult_21_C249_n926, mult_21_C249_n925, mult_21_C249_n924, 
      mult_21_C249_n923, mult_21_C249_n922, mult_21_C249_n921, 
      mult_21_C249_n920, mult_21_C249_n919, mult_21_C249_n918, 
      mult_21_C249_n917, mult_21_C249_n916, mult_21_C249_n915, 
      mult_21_C249_n914, mult_21_C249_n913, mult_21_C249_n912, 
      mult_21_C249_n911, mult_21_C249_n910, mult_21_C249_n909, 
      mult_21_C249_n908, mult_21_C249_n907, mult_21_C249_n906, 
      mult_21_C249_n905, mult_21_C249_n904, mult_21_C249_n903, 
      mult_21_C249_n902, mult_21_C249_n901, mult_21_C249_n900, 
      mult_21_C249_n899, mult_21_C249_n898, mult_21_C249_n897, 
      mult_21_C249_n896, mult_21_C249_n895, mult_21_C249_n894, 
      mult_21_C249_n893, mult_21_C249_n892, mult_21_C249_n891, 
      mult_21_C249_n890, mult_21_C249_n889, mult_21_C249_n888, 
      mult_21_C249_n887, mult_21_C249_n886, mult_21_C249_n885, 
      mult_21_C249_n884, mult_21_C249_n883, mult_21_C249_n882, 
      mult_21_C249_n881, mult_21_C249_n880, mult_21_C249_n879, 
      mult_21_C249_n878, mult_21_C249_n877, mult_21_C249_n876, 
      mult_21_C249_n875, mult_21_C249_n874, mult_21_C249_n873, 
      mult_21_C249_n872, mult_21_C249_n871, mult_21_C249_n870, 
      mult_21_C249_n869, mult_21_C249_n868, mult_21_C249_n867, 
      mult_21_C249_n866, mult_21_C249_n865, mult_21_C249_n864, 
      mult_21_C249_n863, mult_21_C249_n862, mult_21_C249_n861, 
      mult_21_C249_n860, mult_21_C249_n859, mult_21_C249_n858, 
      mult_21_C249_n857, mult_21_C249_n856, mult_21_C249_n855, 
      mult_21_C249_n854, mult_21_C249_n853, mult_21_C249_n852, 
      mult_21_C249_n851, mult_21_C249_n850, mult_21_C249_n849, 
      mult_21_C249_n848, mult_21_C249_n847, mult_21_C249_n846, 
      mult_21_C249_n845, mult_21_C249_n844, mult_21_C249_n843, 
      mult_21_C249_n842, mult_21_C249_n841, mult_21_C249_n840, 
      mult_21_C249_n839, mult_21_C249_n838, mult_21_C249_n837, 
      mult_21_C249_n836, mult_21_C249_n835, mult_21_C249_n834, 
      mult_21_C249_n833, mult_21_C249_n832, mult_21_C249_n831, 
      mult_21_C249_n830, mult_21_C249_n829, mult_21_C249_n828, 
      mult_21_C249_n827, mult_21_C249_n826, mult_21_C249_n825, 
      mult_21_C249_n824, mult_21_C249_n823, mult_21_C249_n822, 
      mult_21_C249_n821, mult_21_C249_n820, mult_21_C249_n819, 
      mult_21_C249_n818, mult_21_C249_n817, mult_21_C249_n816, 
      mult_21_C249_n815, mult_21_C249_n814, mult_21_C249_n813, 
      mult_21_C249_n812, mult_21_C249_n811, mult_21_C249_n810, 
      mult_21_C249_n809, mult_21_C249_n808, mult_21_C249_n807, 
      mult_21_C249_n806, mult_21_C249_n805, mult_21_C249_n804, 
      mult_21_C249_n803, mult_21_C249_n802, mult_21_C249_n801, 
      mult_21_C249_n800, mult_21_C249_n799, mult_21_C249_n798, 
      mult_21_C249_n797, mult_21_C249_n796, mult_21_C249_n795, 
      mult_21_C249_n794, mult_21_C249_n793, mult_21_C249_n792, 
      mult_21_C249_n791, mult_21_C249_n790, mult_21_C249_n789, 
      mult_21_C249_n788, mult_21_C249_n787, mult_21_C249_n786, 
      mult_21_C249_n785, mult_21_C249_n784, mult_21_C249_n783, 
      mult_21_C249_n782, mult_21_C249_n781, mult_21_C249_n780, 
      mult_21_C249_n779, mult_21_C249_n778, mult_21_C249_n777, 
      mult_21_C249_n776, mult_21_C249_n775, mult_21_C249_n774, 
      mult_21_C249_n773, mult_21_C249_n772, mult_21_C249_n771, 
      mult_21_C249_n770, mult_21_C249_n769, mult_21_C249_n768, 
      mult_21_C249_n767, mult_21_C249_n766, mult_21_C249_n765, 
      mult_21_C249_n764, mult_21_C249_n763, mult_21_C249_n762, 
      mult_21_C249_n761, mult_21_C249_n760, mult_21_C249_n759, 
      mult_21_C249_n758, mult_21_C249_n757, mult_21_C249_n756, 
      mult_21_C249_n755, mult_21_C249_n754, mult_21_C249_n753, 
      mult_21_C249_n752, mult_21_C249_n751, mult_21_C249_n750, 
      mult_21_C249_n749, mult_21_C249_n748, mult_21_C249_n747, 
      mult_21_C249_n746, mult_21_C249_n745, mult_21_C249_n744, 
      mult_21_C249_n743, mult_21_C249_n742, mult_21_C249_n741, 
      mult_21_C249_n740, mult_21_C249_n739, mult_21_C249_n738, 
      mult_21_C249_n737, mult_21_C249_n736, mult_21_C249_n735, 
      mult_21_C249_n734, mult_21_C249_n733, mult_21_C249_n732, 
      mult_21_C249_n731, mult_21_C249_n730, mult_21_C249_n729, 
      mult_21_C249_n728, mult_21_C249_n727, mult_21_C249_n726, 
      mult_21_C249_n725, mult_21_C249_n724, mult_21_C249_n723, 
      mult_21_C249_n722, mult_21_C249_n721, mult_21_C249_n720, 
      mult_21_C249_n719, mult_21_C249_n718, mult_21_C249_n717, 
      mult_21_C249_n716, mult_21_C249_n715, mult_21_C249_n714, 
      mult_21_C249_n713, mult_21_C249_n712, mult_21_C249_n711, 
      mult_21_C249_n710, mult_21_C249_n709, mult_21_C249_n708, 
      mult_21_C249_n707, mult_21_C249_n706, mult_21_C249_n705, 
      mult_21_C249_n704, mult_21_C249_n703, mult_21_C249_n702, 
      mult_21_C249_n701, mult_21_C249_n700, mult_21_C249_n699, 
      mult_21_C249_n698, mult_21_C249_n697, mult_21_C249_n696, 
      mult_21_C249_n695, mult_21_C249_n694, mult_21_C249_n693, 
      mult_21_C249_n692, mult_21_C249_n691, mult_21_C249_n690, 
      mult_21_C249_n689, mult_21_C249_n688, mult_21_C249_n687, 
      mult_21_C249_n686, mult_21_C249_n685, mult_21_C249_n684, 
      mult_21_C249_n683, mult_21_C249_n682, mult_21_C249_n681, 
      mult_21_C249_n680, mult_21_C249_n679, mult_21_C249_n678, 
      mult_21_C249_n677, mult_21_C249_n676, mult_21_C249_n675, 
      mult_21_C249_n674, mult_21_C249_n673, mult_21_C249_n672, 
      mult_21_C249_n671, mult_21_C249_n670, mult_21_C249_n669, 
      mult_21_C249_n668, mult_21_C249_n667, mult_21_C249_n666, 
      mult_21_C249_n665, mult_21_C249_n664, mult_21_C249_n663, 
      mult_21_C249_n662, mult_21_C249_n661, mult_21_C249_n660, 
      mult_21_C249_n659, mult_21_C249_n658, mult_21_C249_n657, 
      mult_21_C249_n656, mult_21_C249_n655, mult_21_C249_n654, 
      mult_21_C249_n653, mult_21_C249_n652, mult_21_C249_n651, 
      mult_21_C249_n650, mult_21_C249_n649, mult_21_C249_n648, 
      mult_21_C249_n647, mult_21_C249_n646, mult_21_C249_n645, 
      mult_21_C249_n644, mult_21_C249_n643, mult_21_C249_n642, 
      mult_21_C249_n641, mult_21_C249_n640, mult_21_C249_n639, 
      mult_21_C249_n638, mult_21_C249_n637, mult_21_C249_n636, 
      mult_21_C249_n635, mult_21_C249_n634, mult_21_C249_n633, 
      mult_21_C249_n632, mult_21_C249_n631, mult_21_C249_n630, 
      mult_21_C249_n629, mult_21_C249_n628, mult_21_C249_n627, 
      mult_21_C249_n626, mult_21_C249_n625, mult_21_C249_n624, 
      mult_21_C249_n623, mult_21_C249_n622, mult_21_C249_n621, 
      mult_21_C249_n620, mult_21_C249_n619, mult_21_C249_n618, 
      mult_21_C249_n617, mult_21_C249_n616, mult_21_C249_n615, 
      mult_21_C249_n614, mult_21_C249_n613, mult_21_C249_n612, 
      mult_21_C249_n611, mult_21_C249_n610, mult_21_C249_n609, 
      mult_21_C249_n608, mult_21_C249_n607, mult_21_C249_n606, 
      mult_21_C249_n605, mult_21_C249_n604, mult_21_C249_n603, 
      mult_21_C249_n602, mult_21_C249_n601, mult_21_C249_n600, 
      mult_21_C249_n599, mult_21_C249_n598, mult_21_C249_n597, 
      mult_21_C249_n596, mult_21_C249_n595, mult_21_C249_n594, 
      mult_21_C249_n593, mult_21_C249_n592, mult_21_C249_n591, 
      mult_21_C249_n590, mult_21_C249_n589, mult_21_C249_n588, 
      mult_21_C249_n587, mult_21_C249_n586, mult_21_C249_n585, 
      mult_21_C249_n584, mult_21_C249_n583, mult_21_C249_n582, 
      mult_21_C249_n581, mult_21_C249_n580, mult_21_C249_n579, 
      mult_21_C249_n578, mult_21_C249_n577, mult_21_C249_n576, 
      mult_21_C249_n575, mult_21_C249_n574, mult_21_C249_n573, 
      mult_21_C249_n572, mult_21_C249_n571, mult_21_C249_n570, 
      mult_21_C249_n569, mult_21_C249_n568, mult_21_C249_n567, 
      mult_21_C249_n566, mult_21_C249_n565, mult_21_C249_n564, 
      mult_21_C249_n563, mult_21_C249_n562, mult_21_C249_n561, 
      mult_21_C249_n560, mult_21_C249_n559, mult_21_C249_n558, 
      mult_21_C249_n557, mult_21_C249_n556, mult_21_C249_n555, 
      mult_21_C249_n554, mult_21_C249_n553, mult_21_C249_n552, 
      mult_21_C249_n551, mult_21_C249_n550, mult_21_C249_n549, 
      mult_21_C249_n548, mult_21_C249_n547, mult_21_C249_n546, 
      mult_21_C249_n545, mult_21_C249_n544, mult_21_C249_n543, 
      mult_21_C249_n542, mult_21_C249_n541, mult_21_C249_n540, 
      mult_21_C249_n539, mult_21_C249_n538, mult_21_C249_n537, 
      mult_21_C249_n536, mult_21_C249_n535, mult_21_C249_n534, 
      mult_21_C249_n533, mult_21_C249_n532, mult_21_C249_n531, 
      mult_21_C249_n530, mult_21_C249_n529, mult_21_C249_n528, 
      mult_21_C249_n527, mult_21_C249_n526, mult_21_C249_n525, 
      mult_21_C249_n524, mult_21_C249_n523, mult_21_C249_n522, 
      mult_21_C249_n521, mult_21_C249_n520, mult_21_C249_n519, 
      mult_21_C249_n518, mult_21_C249_n517, mult_21_C249_n516, 
      mult_21_C249_n515, mult_21_C249_n514, mult_21_C249_n513, 
      mult_21_C249_n512, mult_21_C249_n511, mult_21_C249_n510, 
      mult_21_C249_n509, mult_21_C249_n508, mult_21_C249_n507, 
      mult_21_C249_n506, mult_21_C249_n505, mult_21_C249_n504, 
      mult_21_C249_n503, mult_21_C249_n502, mult_21_C249_n501, 
      mult_21_C249_n500, mult_21_C249_n499, mult_21_C249_n498, 
      mult_21_C249_n497, mult_21_C249_n496, mult_21_C249_n495, 
      mult_21_C249_n494, mult_21_C249_n493, mult_21_C249_n492, 
      mult_21_C249_n491, mult_21_C249_n490, mult_21_C249_n489, 
      mult_21_C249_n488, mult_21_C249_n487, mult_21_C249_n486, 
      mult_21_C249_n485, mult_21_C249_n484, mult_21_C249_n483, 
      mult_21_C249_n482, mult_21_C249_n481, mult_21_C249_n480, 
      mult_21_C249_n479, mult_21_C249_n478, mult_21_C249_n477, 
      mult_21_C249_n476, mult_21_C249_n475, mult_21_C249_n474, 
      mult_21_C249_n473, mult_21_C249_n472, mult_21_C249_n471, 
      mult_21_C249_n470, mult_21_C249_n469, mult_21_C249_n468, 
      mult_21_C249_n467, mult_21_C249_n466, mult_21_C249_n465, 
      mult_21_C249_n464, mult_21_C249_n463, mult_21_C249_n462, 
      mult_21_C249_n461, mult_21_C249_n460, mult_21_C249_n459, 
      mult_21_C249_n458, mult_21_C249_n457, mult_21_C249_n456, 
      mult_21_C249_n455, mult_21_C249_n454, mult_21_C249_n453, 
      mult_21_C249_n452, mult_21_C249_n451, mult_21_C249_n450, 
      mult_21_C249_n449, mult_21_C249_n448, mult_21_C249_n447, 
      mult_21_C249_n446, mult_21_C249_n445, mult_21_C249_n444, 
      mult_21_C249_n443, mult_21_C249_n442, mult_21_C249_n441, 
      mult_21_C249_n440, mult_21_C249_n439, mult_21_C249_n438, 
      mult_21_C249_n437, mult_21_C249_n436, mult_21_C249_n435, 
      mult_21_C249_n434, mult_21_C249_n433, mult_21_C249_n432, 
      mult_21_C249_n431, mult_21_C249_n430, mult_21_C249_n429, 
      mult_21_C249_n428, mult_21_C249_n427, mult_21_C249_n426, 
      mult_21_C249_n425, mult_21_C249_n424, mult_21_C249_n423, 
      mult_21_C249_n422, mult_21_C249_n421, mult_21_C249_n420, 
      mult_21_C249_n419, mult_21_C249_n418, mult_21_C249_n417, 
      mult_21_C249_n416, mult_21_C249_n415, mult_21_C249_n414, 
      mult_21_C249_n413, mult_21_C249_n412, mult_21_C249_n411, 
      mult_21_C249_n410, mult_21_C249_n409, mult_21_C249_n408, 
      mult_21_C249_n407, mult_21_C249_n406, mult_21_C249_n405, 
      mult_21_C249_n404, mult_21_C249_n403, mult_21_C249_n402, 
      mult_21_C249_n401, mult_21_C249_n400, mult_21_C249_n399, 
      mult_21_C249_n398, mult_21_C249_n397, mult_21_C249_n396, 
      mult_21_C249_n395, mult_21_C249_n394, mult_21_C249_n393, 
      mult_21_C249_n392, mult_21_C249_n391, mult_21_C249_n390, 
      mult_21_C249_n389, mult_21_C249_n388, mult_21_C249_n387, 
      mult_21_C249_n386, mult_21_C249_n385, mult_21_C249_n384, 
      mult_21_C249_n383, mult_21_C249_n382, mult_21_C249_n381, 
      mult_21_C249_n380, mult_21_C249_n379, mult_21_C249_n378, 
      mult_21_C249_n377, mult_21_C249_n376, mult_21_C249_n375, 
      mult_21_C249_n374, mult_21_C249_n373, mult_21_C249_n372, 
      mult_21_C249_n371, mult_21_C249_n370, mult_21_C249_n369, 
      mult_21_C249_n368, mult_21_C249_n367, mult_21_C249_n366, 
      mult_21_C249_n365, mult_21_C249_n364, mult_21_C249_n363, 
      mult_21_C249_n362, mult_21_C249_n361, mult_21_C249_n360, 
      mult_21_C249_n359, mult_21_C249_n358, mult_21_C249_n357, 
      mult_21_C249_n356, mult_21_C249_n355, mult_21_C249_n354, 
      mult_21_C249_n353, mult_21_C249_n352, mult_21_C249_n351, 
      mult_21_C249_n350, mult_21_C249_n349, mult_21_C249_n348, 
      mult_21_C249_n347, mult_21_C249_n346, mult_21_C249_n345, 
      mult_21_C249_n344, mult_21_C249_n343, mult_21_C249_n342, 
      mult_21_C249_n341, mult_21_C249_n340, mult_21_C249_n339, 
      mult_21_C249_n338, mult_21_C249_n337, mult_21_C249_n336, 
      mult_21_C249_n335, mult_21_C249_n334, mult_21_C249_n333, 
      mult_21_C249_n332, mult_21_C249_n331, mult_21_C249_n330, 
      mult_21_C249_n329, mult_21_C249_n326, mult_21_C249_n324, 
      mult_21_C249_n323, mult_21_C249_n322, mult_21_C249_n319, 
      mult_21_C249_n318, mult_21_C249_n315, mult_21_C249_n314, 
      mult_21_C249_n313, mult_21_C249_n312, mult_21_C249_n310, 
      mult_21_C249_n305, mult_21_C249_n303, mult_21_C249_n302, 
      mult_21_C249_n301, mult_21_C249_n297, mult_21_C249_n296, 
      mult_21_C249_n295, mult_21_C249_n294, mult_21_C249_n293, 
      mult_21_C249_n289, mult_21_C249_n288, mult_21_C249_n287, 
      mult_21_C249_n286, mult_21_C249_n285, mult_21_C249_n284, 
      mult_21_C249_n283, mult_21_C249_n282, mult_21_C249_n281, 
      mult_21_C249_n280, mult_21_C249_n279, mult_21_C249_n278, 
      mult_21_C249_n277, mult_21_C249_n276, mult_21_C249_n275, 
      mult_21_C249_n273, mult_21_C249_n271, mult_21_C249_n270, 
      mult_21_C249_n268, mult_21_C249_n266, mult_21_C249_n265, 
      mult_21_C249_n264, mult_21_C249_n263, mult_21_C249_n262, 
      mult_21_C249_n261, mult_21_C249_n260, mult_21_C249_n259, 
      mult_21_C249_n258, mult_21_C249_n257, mult_21_C249_n256, 
      mult_21_C249_n255, mult_21_C249_n254, mult_21_C249_n253, 
      mult_21_C249_n251, mult_21_C249_n249, mult_21_C249_n248, 
      mult_21_C249_n246, mult_21_C249_n244, mult_21_C249_n243, 
      mult_21_C249_n242, mult_21_C249_n241, mult_21_C249_n240, 
      mult_21_C249_n239, mult_21_C249_n238, mult_21_C249_n237, 
      mult_21_C249_n236, mult_21_C249_n235, mult_21_C249_n234, 
      mult_21_C249_n233, mult_21_C249_n232, mult_21_C249_n231, 
      mult_21_C249_n230, mult_21_C249_n229, mult_21_C249_n227, 
      mult_21_C249_n226, mult_21_C249_n225, mult_21_C249_n224, 
      mult_21_C249_n223, mult_21_C249_n222, mult_21_C249_n221, 
      mult_21_C249_n219, mult_21_C249_n217, mult_21_C249_n216, 
      mult_21_C249_n215, mult_21_C249_n214, mult_21_C249_n211, 
      mult_21_C249_n209, mult_21_C249_n208, mult_21_C249_n207, 
      mult_21_C249_n206, mult_21_C249_n204, mult_21_C249_n202, 
      mult_21_C249_n201, mult_21_C249_n200, mult_21_C249_n199, 
      mult_21_C249_n197, mult_21_C249_n195, mult_21_C249_n194, 
      mult_21_C249_n190, mult_21_C249_n189, mult_21_C249_n188, 
      mult_21_C249_n187, mult_21_C249_n185, mult_21_C249_n184, 
      mult_21_C249_n183, mult_21_C249_n182, mult_21_C249_n181, 
      mult_21_C249_n180, mult_21_C249_n179, mult_21_C249_n178, 
      mult_21_C249_n176, mult_21_C249_n175, mult_21_C249_n174, 
      mult_21_C249_n173, mult_21_C249_n172, mult_21_C249_n171, 
      mult_21_C249_n170, mult_21_C249_n169, mult_21_C249_n168, 
      mult_21_C249_n167, mult_21_C249_n166, mult_21_C249_n165, 
      mult_21_C249_n164, mult_21_C249_n163, mult_21_C249_n162, 
      mult_21_C249_n161, mult_21_C249_n160, mult_21_C249_n159, 
      mult_21_C249_n158, mult_21_C249_n157, mult_21_C249_n156, 
      mult_21_C249_n155, mult_21_C249_n106, mult_21_C249_n105, 
      mult_21_C249_n104, mult_21_C249_n103, mult_21_C249_n101, mult_21_C249_n99
      , mult_21_C249_n98, mult_21_C249_n96, mult_21_C249_n94, mult_21_C249_n93,
      mult_21_C249_n91, mult_21_C249_n89, mult_21_C249_n88, mult_21_C249_n86, 
      mult_21_C249_n84, mult_21_C249_n83, mult_21_C249_n81, mult_21_C249_n79, 
      mult_21_C249_n78, mult_21_C249_n76, mult_21_C249_n73, mult_21_C249_n71, 
      mult_21_C249_n69, mult_21_C249_n66, mult_21_C249_n63, mult_21_C249_n61, 
      mult_21_C249_n58, mult_21_C249_n56, mult_21_C249_n53, mult_21_C249_n50, 
      mult_21_C249_n48, mult_21_C249_n45, mult_21_C249_n42, mult_21_C249_n38, 
      mult_21_C249_n30, mult_21_C249_n22, mult_21_C249_n14, mult_21_C249_n8, 
      mult_21_C249_n6, mult_21_C249_n3 : std_logic;

begin
   avs_readdata <= ( avs_readdata_31_port, avs_readdata_30_port, 
      avs_readdata_29_port, avs_readdata_28_port, avs_readdata_27_port, 
      avs_readdata_26_port, avs_readdata_25_port, avs_readdata_24_port, 
      avs_readdata_23_port, avs_readdata_22_port, avs_readdata_21_port, 
      avs_readdata_20_port, avs_readdata_19_port, avs_readdata_18_port, 
      avs_readdata_17_port, avs_readdata_16_port, avs_readdata_15_port, 
      avs_readdata_14_port, avs_readdata_13_port, avs_readdata_12_port, 
      avs_readdata_11_port, avs_readdata_10_port, avs_readdata_9_port, 
      avs_readdata_8_port, avs_readdata_7_port, avs_readdata_6_port, 
      avs_readdata_5_port, avs_readdata_4_port, avs_readdata_3_port, 
      avs_readdata_2_port, avs_readdata_1_port, avs_readdata_0_port );
   clk_out <= clk;
   stop_sim <= stop_sim_port;
   
   U3 : OAI22D1 port map( A1 => N63, A2 => n4, B1 => n5, B2 => n813, Z => n201)
                           ;
   U4 : AOI21D1 port map( A1 => out_busy, A2 => n810, B => n801, Z => n5);
   U7 : AOI22D1 port map( A1 => N1978, A2 => n268, B1 => N2010, B2 => n698, Z 
                           => n10);
   U9 : AOI22D1 port map( A1 => N2011, A2 => n12, B1 => avs_readdata_30_port, 
                           B2 => n700, Z => n15);
   U12 : AOI22D1 port map( A1 => N1980, A2 => n268, B1 => N2012, B2 => n698, Z 
                           => n16);
   U14 : AOI22D1 port map( A1 => N2013, A2 => n698, B1 => avs_readdata_28_port,
                           B2 => n700, Z => n18);
   U17 : AOI22D1 port map( A1 => N1982, A2 => n268, B1 => N2014, B2 => n698, Z 
                           => n19);
   U19 : AOI22D1 port map( A1 => N2015, A2 => n698, B1 => avs_readdata_26_port,
                           B2 => n700, Z => n21);
   U22 : AOI22D1 port map( A1 => N1984, A2 => n268, B1 => N2016, B2 => n698, Z 
                           => n22);
   U24 : AOI22D1 port map( A1 => N2017, A2 => n698, B1 => avs_readdata_24_port,
                           B2 => n700, Z => n24);
   U27 : AOI22D1 port map( A1 => N1986, A2 => n268, B1 => N2018, B2 => n698, Z 
                           => n25);
   U29 : AOI22D1 port map( A1 => N2019, A2 => n12, B1 => avs_readdata_22_port, 
                           B2 => n700, Z => n27);
   U32 : AOI22D1 port map( A1 => N1988, A2 => n268, B1 => N2020, B2 => n698, Z 
                           => n28);
   U34 : AOI22D1 port map( A1 => N2021, A2 => n12, B1 => avs_readdata_20_port, 
                           B2 => n700, Z => n30);
   U37 : AOI22D1 port map( A1 => N1990, A2 => n268, B1 => N2022, B2 => n698, Z 
                           => n31);
   U39 : AOI22D1 port map( A1 => N2023, A2 => n12, B1 => avs_readdata_18_port, 
                           B2 => n700, Z => n33);
   U42 : AOI22D1 port map( A1 => N1992, A2 => n268, B1 => N2024, B2 => n698, Z 
                           => n34);
   U44 : AOI22D1 port map( A1 => N2025, A2 => n12, B1 => avs_readdata_16_port, 
                           B2 => n700, Z => n36);
   U47 : AOI22D1 port map( A1 => N1994, A2 => n268, B1 => N2026, B2 => n698, Z 
                           => n37);
   U49 : AOI22D1 port map( A1 => N2027, A2 => n12, B1 => avs_readdata_14_port, 
                           B2 => n700, Z => n39);
   U52 : AOI22D1 port map( A1 => N1996, A2 => n268, B1 => N2028, B2 => n12, Z 
                           => n40);
   U54 : AOI22D1 port map( A1 => N2029, A2 => n12, B1 => avs_readdata_12_port, 
                           B2 => n700, Z => n42);
   U57 : AOI22D1 port map( A1 => N1998, A2 => n268, B1 => N2030, B2 => n12, Z 
                           => n43);
   U59 : AOI22D1 port map( A1 => N2031, A2 => n12, B1 => avs_readdata_10_port, 
                           B2 => n700, Z => n45);
   U62 : AOI22D1 port map( A1 => N2000, A2 => n268, B1 => N2032, B2 => n12, Z 
                           => n46);
   U64 : AOI22D1 port map( A1 => N2033, A2 => n12, B1 => avs_readdata_8_port, 
                           B2 => n700, Z => n48);
   U67 : AOI22D1 port map( A1 => N2002, A2 => n268, B1 => N2034, B2 => n698, Z 
                           => n49);
   U69 : AOI22D1 port map( A1 => N2035, A2 => n12, B1 => avs_readdata_6_port, 
                           B2 => n700, Z => n51);
   U72 : AOI22D1 port map( A1 => N2004, A2 => n268, B1 => N2036, B2 => n698, Z 
                           => n52);
   U74 : AOI22D1 port map( A1 => N2037, A2 => n12, B1 => avs_readdata_4_port, 
                           B2 => n700, Z => n54);
   U77 : AOI22D1 port map( A1 => N2006, A2 => n268, B1 => N2038, B2 => n698, Z 
                           => n55);
   U79 : AOI22D1 port map( A1 => N2039, A2 => n12, B1 => avs_readdata_2_port, 
                           B2 => n700, Z => n57);
   U82 : AOI22D1 port map( A1 => N2008, A2 => n268, B1 => N2040, B2 => n698, Z 
                           => n58);
   U84 : AOI22D1 port map( A1 => N2041, A2 => n698, B1 => avs_readdata_0_port, 
                           B2 => n700, Z => n6100);
   U94 : AOI21D1 port map( A1 => n798, A2 => in_trigger, B => n72, Z => n70);
   U95 : OAI22D1 port map( A1 => n6400, A2 => n73, B1 => n74, B2 => n802, Z => 
                           n72);
   U96 : AOI22D1 port map( A1 => in_busy, A2 => n307, B1 => out_busy, B2 => 
                           n306, Z => n73);
   U97 : EXNOR2D1 port map( A1 => n811, A2 => n76, Z => n234);
   U98 : AOI22D1 port map( A1 => n77, A2 => out_busy, B1 => n811, B2 => n802, Z
                           => n76);
   U100 : OAI22D1 port map( A1 => n813, A2 => n4, B1 => n79, B2 => n696, Z => 
                           n235);
   U103 : OAI32D1 port map( A1 => n801, A2 => N62, A3 => n811, B1 => n810, B2 
                           => n81, Z => n236);
   U105 : OAI32D1 port map( A1 => n812, A2 => n811, A3 => n78, B1 => out_busy, 
                           B2 => n802, Z => n81);
   U111 : OAI211D1 port map( A1 => n808, A2 => n84, B => n85, C => n86, Z => 
                           n237);
   U113 : OAI22D1 port map( A1 => n800, A2 => n88, B1 => n89, B2 => n809, Z => 
                           n238);
   U115 : EXNOR2D1 port map( A1 => in_busy, A2 => n161, Z => n239);
   U117 : AOI22D1 port map( A1 => avs_writedata(0), A2 => n797, B1 => 
                           out_trigger, B2 => n74, Z => n92);
   U122 : AOI22D1 port map( A1 => avs_writedata(0), A2 => n798, B1 => 
                           in_trigger, B2 => n96, Z => n95);
   U125 : EXNOR2D1 port map( A1 => n811, A2 => n697, Z => n154);
   U126 : EXNOR2D1 port map( A1 => n803, A2 => in_busy, Z => n156);
   U130 : AOI22D1 port map( A1 => odd, A2 => n91, B1 => n101, B2 => in_busy, Z 
                           => n100);
   U131 : OAI21D1 port map( A1 => in_counter_1_port, A2 => n806, B => n804, Z 
                           => n91);
   U200 : OA21M20D1 port map( A1 => n806, A2 => in_trigger, B => n176, Z => 
                           n161);
   comp_res_reg_4_30 : DFFRPQ1 port map( D => N3391, CK => clk, RB => resetn, Q
                           => comp_res_30_port);
   comp_res_reg_4_28 : DFFRPQ1 port map( D => N3389, CK => clk, RB => resetn, Q
                           => comp_res_28_port);
   comp_res_reg_4_26 : DFFRPQ1 port map( D => N3387, CK => clk, RB => resetn, Q
                           => comp_res_26_port);
   comp_res_reg_4_24 : DFFRPQ1 port map( D => N3385, CK => clk, RB => resetn, Q
                           => comp_res_24_port);
   comp_res_reg_4_22 : DFFRPQ1 port map( D => N3383, CK => clk, RB => resetn, Q
                           => comp_res_22_port);
   comp_res_reg_4_20 : DFFRPQ1 port map( D => N3381, CK => clk, RB => resetn, Q
                           => comp_res_20_port);
   comp_res_reg_4_18 : DFFRPQ1 port map( D => N3379, CK => clk, RB => resetn, Q
                           => comp_res_18_port);
   comp_res_reg_4_16 : DFFRPQ1 port map( D => N3377, CK => clk, RB => resetn, Q
                           => comp_res_16_port);
   comp_res_reg_4_14 : DFFRPQ1 port map( D => N3375, CK => clk, RB => resetn, Q
                           => comp_res_14_port);
   comp_res_reg_4_12 : DFFRPQ1 port map( D => N3373, CK => clk, RB => resetn, Q
                           => comp_res_12_port);
   comp_res_reg_4_10 : DFFRPQ1 port map( D => N3371, CK => clk, RB => resetn, Q
                           => comp_res_10_port);
   comp_res_reg_4_8 : DFFRPQ1 port map( D => N3369, CK => clk, RB => resetn, Q 
                           => comp_res_8_port);
   comp_res_reg_4_6 : DFFRPQ1 port map( D => N3367, CK => clk, RB => resetn, Q 
                           => comp_res_6_port);
   comp_res_reg_4_4 : DFFRPQ1 port map( D => N3365, CK => clk, RB => resetn, Q 
                           => comp_res_4_port);
   comp_res_reg_4_2 : DFFRPQ1 port map( D => N3363, CK => clk, RB => resetn, Q 
                           => comp_res_2_port);
   comp_res_reg_4_0 : DFFRPQ1 port map( D => N3361, CK => clk, RB => resetn, Q 
                           => comp_res_0_port);
   comp_res_reg_4_31 : DFFRPQ1 port map( D => N3392, CK => clk, RB => resetn, Q
                           => comp_res_31_port);
   comp_res_reg_4_29 : DFFRPQ1 port map( D => N3390, CK => clk, RB => resetn, Q
                           => comp_res_29_port);
   comp_res_reg_4_27 : DFFRPQ1 port map( D => N3388, CK => clk, RB => resetn, Q
                           => comp_res_27_port);
   comp_res_reg_4_25 : DFFRPQ1 port map( D => N3386, CK => clk, RB => resetn, Q
                           => comp_res_25_port);
   comp_res_reg_4_23 : DFFRPQ1 port map( D => N3384, CK => clk, RB => resetn, Q
                           => comp_res_23_port);
   comp_res_reg_4_21 : DFFRPQ1 port map( D => N3382, CK => clk, RB => resetn, Q
                           => comp_res_21_port);
   comp_res_reg_4_19 : DFFRPQ1 port map( D => N3380, CK => clk, RB => resetn, Q
                           => comp_res_19_port);
   comp_res_reg_4_17 : DFFRPQ1 port map( D => N3378, CK => clk, RB => resetn, Q
                           => comp_res_17_port);
   comp_res_reg_4_15 : DFFRPQ1 port map( D => N3376, CK => clk, RB => resetn, Q
                           => comp_res_15_port);
   comp_res_reg_4_13 : DFFRPQ1 port map( D => N3374, CK => clk, RB => resetn, Q
                           => comp_res_13_port);
   comp_res_reg_4_11 : DFFRPQ1 port map( D => N3372, CK => clk, RB => resetn, Q
                           => comp_res_11_port);
   comp_res_reg_4_9 : DFFRPQ1 port map( D => N3370, CK => clk, RB => resetn, Q 
                           => comp_res_9_port);
   comp_res_reg_4_7 : DFFRPQ1 port map( D => N3368, CK => clk, RB => resetn, Q 
                           => comp_res_7_port);
   comp_res_reg_4_5 : DFFRPQ1 port map( D => N3366, CK => clk, RB => resetn, Q 
                           => comp_res_5_port);
   comp_res_reg_4_3 : DFFRPQ1 port map( D => N3364, CK => clk, RB => resetn, Q 
                           => comp_res_3_port);
   comp_res_reg_4_1 : DFFRPQ1 port map( D => N3362, CK => clk, RB => resetn, Q 
                           => comp_res_1_port);
   comp_res_reg_3_30 : DFFRPQ1 port map( D => N3359, CK => clk, RB => resetn, Q
                           => comp_res_62_port);
   comp_res_reg_3_28 : DFFRPQ1 port map( D => N3357, CK => clk, RB => resetn, Q
                           => comp_res_60_port);
   comp_res_reg_3_26 : DFFRPQ1 port map( D => N3355, CK => clk, RB => resetn, Q
                           => comp_res_58_port);
   comp_res_reg_3_24 : DFFRPQ1 port map( D => N3353, CK => clk, RB => resetn, Q
                           => comp_res_56_port);
   comp_res_reg_3_22 : DFFRPQ1 port map( D => N3351, CK => clk, RB => resetn, Q
                           => comp_res_54_port);
   comp_res_reg_3_20 : DFFRPQ1 port map( D => N3349, CK => clk, RB => resetn, Q
                           => comp_res_52_port);
   comp_res_reg_3_18 : DFFRPQ1 port map( D => N3347, CK => clk, RB => resetn, Q
                           => comp_res_50_port);
   comp_res_reg_3_16 : DFFRPQ1 port map( D => N3345, CK => clk, RB => resetn, Q
                           => comp_res_48_port);
   comp_res_reg_3_14 : DFFRPQ1 port map( D => N3343, CK => clk, RB => resetn, Q
                           => comp_res_46_port);
   comp_res_reg_3_12 : DFFRPQ1 port map( D => N3341, CK => clk, RB => resetn, Q
                           => comp_res_44_port);
   comp_res_reg_3_10 : DFFRPQ1 port map( D => N3339, CK => clk, RB => resetn, Q
                           => comp_res_42_port);
   comp_res_reg_3_8 : DFFRPQ1 port map( D => N3337, CK => clk, RB => resetn, Q 
                           => comp_res_40_port);
   comp_res_reg_3_6 : DFFRPQ1 port map( D => N3335, CK => clk, RB => resetn, Q 
                           => comp_res_38_port);
   comp_res_reg_3_4 : DFFRPQ1 port map( D => N3333, CK => clk, RB => resetn, Q 
                           => comp_res_36_port);
   comp_res_reg_3_2 : DFFRPQ1 port map( D => N3331, CK => clk, RB => resetn, Q 
                           => comp_res_34_port);
   comp_res_reg_2_30 : DFFRPQ1 port map( D => N3327, CK => clk, RB => resetn, Q
                           => comp_res_94_port);
   comp_res_reg_2_28 : DFFRPQ1 port map( D => N3325, CK => clk, RB => resetn, Q
                           => comp_res_92_port);
   comp_res_reg_2_26 : DFFRPQ1 port map( D => N3323, CK => clk, RB => resetn, Q
                           => comp_res_90_port);
   comp_res_reg_2_24 : DFFRPQ1 port map( D => N3321, CK => clk, RB => resetn, Q
                           => comp_res_88_port);
   comp_res_reg_2_22 : DFFRPQ1 port map( D => N3319, CK => clk, RB => resetn, Q
                           => comp_res_86_port);
   comp_res_reg_2_20 : DFFRPQ1 port map( D => N3317, CK => clk, RB => resetn, Q
                           => comp_res_84_port);
   comp_res_reg_2_18 : DFFRPQ1 port map( D => N3315, CK => clk, RB => resetn, Q
                           => comp_res_82_port);
   comp_res_reg_2_16 : DFFRPQ1 port map( D => N3313, CK => clk, RB => resetn, Q
                           => comp_res_80_port);
   comp_res_reg_2_14 : DFFRPQ1 port map( D => N3311, CK => clk, RB => resetn, Q
                           => comp_res_78_port);
   comp_res_reg_2_12 : DFFRPQ1 port map( D => N3309, CK => clk, RB => resetn, Q
                           => comp_res_76_port);
   comp_res_reg_2_10 : DFFRPQ1 port map( D => N3307, CK => clk, RB => resetn, Q
                           => comp_res_74_port);
   comp_res_reg_2_8 : DFFRPQ1 port map( D => N3305, CK => clk, RB => resetn, Q 
                           => comp_res_72_port);
   comp_res_reg_2_6 : DFFRPQ1 port map( D => N3303, CK => clk, RB => resetn, Q 
                           => comp_res_70_port);
   comp_res_reg_2_4 : DFFRPQ1 port map( D => N3301, CK => clk, RB => resetn, Q 
                           => comp_res_68_port);
   comp_res_reg_2_2 : DFFRPQ1 port map( D => N3299, CK => clk, RB => resetn, Q 
                           => comp_res_66_port);
   comp_res_reg_1_30 : DFFRPQ1 port map( D => N3295, CK => clk, RB => resetn, Q
                           => comp_res_126_port);
   comp_res_reg_1_28 : DFFRPQ1 port map( D => N3293, CK => clk, RB => resetn, Q
                           => comp_res_124_port);
   comp_res_reg_1_26 : DFFRPQ1 port map( D => N3291, CK => clk, RB => resetn, Q
                           => comp_res_122_port);
   comp_res_reg_1_24 : DFFRPQ1 port map( D => N3289, CK => clk, RB => resetn, Q
                           => comp_res_120_port);
   comp_res_reg_1_22 : DFFRPQ1 port map( D => N3287, CK => clk, RB => resetn, Q
                           => comp_res_118_port);
   comp_res_reg_1_20 : DFFRPQ1 port map( D => N3285, CK => clk, RB => resetn, Q
                           => comp_res_116_port);
   comp_res_reg_1_18 : DFFRPQ1 port map( D => N3283, CK => clk, RB => resetn, Q
                           => comp_res_114_port);
   comp_res_reg_1_16 : DFFRPQ1 port map( D => N3281, CK => clk, RB => resetn, Q
                           => comp_res_112_port);
   comp_res_reg_1_14 : DFFRPQ1 port map( D => N3279, CK => clk, RB => resetn, Q
                           => comp_res_110_port);
   comp_res_reg_1_12 : DFFRPQ1 port map( D => N3277, CK => clk, RB => resetn, Q
                           => comp_res_108_port);
   comp_res_reg_1_10 : DFFRPQ1 port map( D => N3275, CK => clk, RB => resetn, Q
                           => comp_res_106_port);
   comp_res_reg_1_8 : DFFRPQ1 port map( D => N3273, CK => clk, RB => resetn, Q 
                           => comp_res_104_port);
   comp_res_reg_1_6 : DFFRPQ1 port map( D => N3271, CK => clk, RB => resetn, Q 
                           => comp_res_102_port);
   comp_res_reg_1_4 : DFFRPQ1 port map( D => N3269, CK => clk, RB => resetn, Q 
                           => comp_res_100_port);
   comp_res_reg_1_2 : DFFRPQ1 port map( D => N3267, CK => clk, RB => resetn, Q 
                           => comp_res_98_port);
   comp_res_reg_0_30 : DFFRPQ1 port map( D => N3263, CK => clk, RB => resetn, Q
                           => comp_res_158_port);
   comp_res_reg_0_28 : DFFRPQ1 port map( D => N3261, CK => clk, RB => resetn, Q
                           => comp_res_156_port);
   comp_res_reg_0_26 : DFFRPQ1 port map( D => N3259, CK => clk, RB => resetn, Q
                           => comp_res_154_port);
   comp_res_reg_0_24 : DFFRPQ1 port map( D => N3257, CK => clk, RB => resetn, Q
                           => comp_res_152_port);
   comp_res_reg_0_22 : DFFRPQ1 port map( D => N3255, CK => clk, RB => resetn, Q
                           => comp_res_150_port);
   comp_res_reg_0_20 : DFFRPQ1 port map( D => N3253, CK => clk, RB => resetn, Q
                           => comp_res_148_port);
   comp_res_reg_0_18 : DFFRPQ1 port map( D => N3251, CK => clk, RB => resetn, Q
                           => comp_res_146_port);
   comp_res_reg_0_16 : DFFRPQ1 port map( D => N3249, CK => clk, RB => resetn, Q
                           => comp_res_144_port);
   comp_res_reg_0_14 : DFFRPQ1 port map( D => N3247, CK => clk, RB => resetn, Q
                           => comp_res_142_port);
   comp_res_reg_0_12 : DFFRPQ1 port map( D => N3245, CK => clk, RB => resetn, Q
                           => comp_res_140_port);
   comp_res_reg_0_10 : DFFRPQ1 port map( D => N3243, CK => clk, RB => resetn, Q
                           => comp_res_138_port);
   comp_res_reg_0_8 : DFFRPQ1 port map( D => N3241, CK => clk, RB => resetn, Q 
                           => comp_res_136_port);
   comp_res_reg_0_6 : DFFRPQ1 port map( D => N3239, CK => clk, RB => resetn, Q 
                           => comp_res_134_port);
   comp_res_reg_0_4 : DFFRPQ1 port map( D => N3237, CK => clk, RB => resetn, Q 
                           => comp_res_132_port);
   comp_res_reg_0_2 : DFFRPQ1 port map( D => N3235, CK => clk, RB => resetn, Q 
                           => comp_res_130_port);
   comp_res_reg_3_0 : DFFRPQ1 port map( D => N3329, CK => clk, RB => resetn, Q 
                           => comp_res_32_port);
   comp_res_reg_2_0 : DFFRPQ1 port map( D => N3297, CK => clk, RB => resetn, Q 
                           => comp_res_64_port);
   comp_res_reg_1_0 : DFFRPQ1 port map( D => N3265, CK => clk, RB => resetn, Q 
                           => comp_res_96_port);
   comp_res_reg_0_0 : DFFRPQ1 port map( D => N3233, CK => clk, RB => resetn, Q 
                           => comp_res_128_port);
   in_buf_reg_7_31 : DFERPQ1 port map( D => siso_data_in(15), CEB => n176, CK 
                           => clk, RB => resetn, Q => in_buf_31_port);
   in_buf_reg_7_29 : DFERPQ1 port map( D => siso_data_in(13), CEB => n176, CK 
                           => clk, RB => resetn, Q => in_buf_29_port);
   in_buf_reg_7_27 : DFERPQ1 port map( D => siso_data_in(11), CEB => n176, CK 
                           => clk, RB => resetn, Q => in_buf_27_port);
   in_buf_reg_7_25 : DFERPQ1 port map( D => siso_data_in(9), CEB => n176, CK =>
                           clk, RB => resetn, Q => in_buf_25_port);
   in_buf_reg_7_23 : DFERPQ1 port map( D => siso_data_in(7), CEB => n176, CK =>
                           clk, RB => resetn, Q => in_buf_23_port);
   in_buf_reg_7_21 : DFERPQ1 port map( D => siso_data_in(5), CEB => n176, CK =>
                           clk, RB => resetn, Q => in_buf_21_port);
   in_buf_reg_7_19 : DFERPQ1 port map( D => siso_data_in(3), CEB => n176, CK =>
                           clk, RB => resetn, Q => in_buf_19_port);
   in_buf_reg_7_17 : DFERPQ1 port map( D => siso_data_in(1), CEB => n176, CK =>
                           clk, RB => resetn, Q => in_buf_17_port);
   in_buf_reg_7_15 : DFERPQ1 port map( D => siso_data_in(15), CEB => n177, CK 
                           => clk, RB => resetn, Q => in_buf_15_port);
   in_buf_reg_7_13 : DFERPQ1 port map( D => siso_data_in(13), CEB => n177, CK 
                           => clk, RB => resetn, Q => in_buf_13_port);
   in_buf_reg_7_11 : DFERPQ1 port map( D => siso_data_in(11), CEB => n177, CK 
                           => clk, RB => resetn, Q => in_buf_11_port);
   in_buf_reg_7_9 : DFERPQ1 port map( D => siso_data_in(9), CEB => n177, CK => 
                           clk, RB => resetn, Q => in_buf_9_port);
   in_buf_reg_7_7 : DFERPQ1 port map( D => siso_data_in(7), CEB => n177, CK => 
                           clk, RB => resetn, Q => in_buf_7_port);
   in_buf_reg_7_5 : DFERPQ1 port map( D => siso_data_in(5), CEB => n177, CK => 
                           clk, RB => resetn, Q => in_buf_5_port);
   in_buf_reg_7_3 : DFERPQ1 port map( D => siso_data_in(3), CEB => n177, CK => 
                           clk, RB => resetn, Q => in_buf_3_port);
   in_buf_reg_7_1 : DFERPQ1 port map( D => siso_data_in(1), CEB => n177, CK => 
                           clk, RB => resetn, Q => in_buf_1_port);
   comp_res_reg_3_31 : DFFRPQ1 port map( D => N3360, CK => clk, RB => resetn, Q
                           => comp_res_63_port);
   comp_res_reg_3_29 : DFFRPQ1 port map( D => N3358, CK => clk, RB => resetn, Q
                           => comp_res_61_port);
   comp_res_reg_3_27 : DFFRPQ1 port map( D => N3356, CK => clk, RB => resetn, Q
                           => comp_res_59_port);
   comp_res_reg_3_25 : DFFRPQ1 port map( D => N3354, CK => clk, RB => resetn, Q
                           => comp_res_57_port);
   comp_res_reg_3_23 : DFFRPQ1 port map( D => N3352, CK => clk, RB => resetn, Q
                           => comp_res_55_port);
   comp_res_reg_3_21 : DFFRPQ1 port map( D => N3350, CK => clk, RB => resetn, Q
                           => comp_res_53_port);
   comp_res_reg_3_19 : DFFRPQ1 port map( D => N3348, CK => clk, RB => resetn, Q
                           => comp_res_51_port);
   comp_res_reg_3_17 : DFFRPQ1 port map( D => N3346, CK => clk, RB => resetn, Q
                           => comp_res_49_port);
   comp_res_reg_3_15 : DFFRPQ1 port map( D => N3344, CK => clk, RB => resetn, Q
                           => comp_res_47_port);
   comp_res_reg_3_13 : DFFRPQ1 port map( D => N3342, CK => clk, RB => resetn, Q
                           => comp_res_45_port);
   comp_res_reg_3_11 : DFFRPQ1 port map( D => N3340, CK => clk, RB => resetn, Q
                           => comp_res_43_port);
   comp_res_reg_3_9 : DFFRPQ1 port map( D => N3338, CK => clk, RB => resetn, Q 
                           => comp_res_41_port);
   comp_res_reg_3_7 : DFFRPQ1 port map( D => N3336, CK => clk, RB => resetn, Q 
                           => comp_res_39_port);
   comp_res_reg_3_5 : DFFRPQ1 port map( D => N3334, CK => clk, RB => resetn, Q 
                           => comp_res_37_port);
   comp_res_reg_3_3 : DFFRPQ1 port map( D => N3332, CK => clk, RB => resetn, Q 
                           => comp_res_35_port);
   comp_res_reg_3_1 : DFFRPQ1 port map( D => N3330, CK => clk, RB => resetn, Q 
                           => comp_res_33_port);
   comp_res_reg_2_31 : DFFRPQ1 port map( D => N3328, CK => clk, RB => resetn, Q
                           => comp_res_95_port);
   comp_res_reg_2_29 : DFFRPQ1 port map( D => N3326, CK => clk, RB => resetn, Q
                           => comp_res_93_port);
   comp_res_reg_2_27 : DFFRPQ1 port map( D => N3324, CK => clk, RB => resetn, Q
                           => comp_res_91_port);
   comp_res_reg_2_25 : DFFRPQ1 port map( D => N3322, CK => clk, RB => resetn, Q
                           => comp_res_89_port);
   comp_res_reg_2_23 : DFFRPQ1 port map( D => N3320, CK => clk, RB => resetn, Q
                           => comp_res_87_port);
   comp_res_reg_2_21 : DFFRPQ1 port map( D => N3318, CK => clk, RB => resetn, Q
                           => comp_res_85_port);
   comp_res_reg_2_19 : DFFRPQ1 port map( D => N3316, CK => clk, RB => resetn, Q
                           => comp_res_83_port);
   comp_res_reg_2_17 : DFFRPQ1 port map( D => N3314, CK => clk, RB => resetn, Q
                           => comp_res_81_port);
   comp_res_reg_2_15 : DFFRPQ1 port map( D => N3312, CK => clk, RB => resetn, Q
                           => comp_res_79_port);
   comp_res_reg_2_13 : DFFRPQ1 port map( D => N3310, CK => clk, RB => resetn, Q
                           => comp_res_77_port);
   comp_res_reg_2_11 : DFFRPQ1 port map( D => N3308, CK => clk, RB => resetn, Q
                           => comp_res_75_port);
   comp_res_reg_2_9 : DFFRPQ1 port map( D => N3306, CK => clk, RB => resetn, Q 
                           => comp_res_73_port);
   comp_res_reg_2_7 : DFFRPQ1 port map( D => N3304, CK => clk, RB => resetn, Q 
                           => comp_res_71_port);
   comp_res_reg_2_5 : DFFRPQ1 port map( D => N3302, CK => clk, RB => resetn, Q 
                           => comp_res_69_port);
   comp_res_reg_2_3 : DFFRPQ1 port map( D => N3300, CK => clk, RB => resetn, Q 
                           => comp_res_67_port);
   comp_res_reg_2_1 : DFFRPQ1 port map( D => N3298, CK => clk, RB => resetn, Q 
                           => comp_res_65_port);
   in_buf_reg_3_31 : DFERPQ1 port map( D => siso_data_in(15), CEB => n168, CK 
                           => clk, RB => resetn, Q => in_buf_159_port);
   in_buf_reg_3_29 : DFERPQ1 port map( D => siso_data_in(13), CEB => n168, CK 
                           => clk, RB => resetn, Q => in_buf_157_port);
   in_buf_reg_3_27 : DFERPQ1 port map( D => siso_data_in(11), CEB => n168, CK 
                           => clk, RB => resetn, Q => in_buf_155_port);
   in_buf_reg_3_25 : DFERPQ1 port map( D => siso_data_in(9), CEB => n168, CK =>
                           clk, RB => resetn, Q => in_buf_153_port);
   in_buf_reg_3_23 : DFERPQ1 port map( D => siso_data_in(7), CEB => n168, CK =>
                           clk, RB => resetn, Q => in_buf_151_port);
   in_buf_reg_3_21 : DFERPQ1 port map( D => siso_data_in(5), CEB => n168, CK =>
                           clk, RB => resetn, Q => in_buf_149_port);
   in_buf_reg_3_19 : DFERPQ1 port map( D => siso_data_in(3), CEB => n168, CK =>
                           clk, RB => resetn, Q => in_buf_147_port);
   in_buf_reg_3_17 : DFERPQ1 port map( D => siso_data_in(1), CEB => n168, CK =>
                           clk, RB => resetn, Q => in_buf_145_port);
   in_buf_reg_3_15 : DFERPQ1 port map( D => siso_data_in(15), CEB => n169, CK 
                           => clk, RB => resetn, Q => in_buf_143_port);
   in_buf_reg_3_13 : DFERPQ1 port map( D => siso_data_in(13), CEB => n169, CK 
                           => clk, RB => resetn, Q => in_buf_141_port);
   in_buf_reg_3_11 : DFERPQ1 port map( D => siso_data_in(11), CEB => n169, CK 
                           => clk, RB => resetn, Q => in_buf_139_port);
   in_buf_reg_3_9 : DFERPQ1 port map( D => siso_data_in(9), CEB => n169, CK => 
                           clk, RB => resetn, Q => in_buf_137_port);
   in_buf_reg_3_7 : DFERPQ1 port map( D => siso_data_in(7), CEB => n169, CK => 
                           clk, RB => resetn, Q => in_buf_135_port);
   in_buf_reg_3_5 : DFERPQ1 port map( D => siso_data_in(5), CEB => n169, CK => 
                           clk, RB => resetn, Q => in_buf_133_port);
   in_buf_reg_3_3 : DFERPQ1 port map( D => siso_data_in(3), CEB => n169, CK => 
                           clk, RB => resetn, Q => in_buf_131_port);
   in_buf_reg_3_1 : DFERPQ1 port map( D => siso_data_in(1), CEB => n169, CK => 
                           clk, RB => resetn, Q => in_buf_129_port);
   in_buf_reg_2_31 : DFERPQ1 port map( D => siso_data_in(15), CEB => n166, CK 
                           => clk, RB => resetn, Q => in_buf_191_port);
   in_buf_reg_2_29 : DFERPQ1 port map( D => siso_data_in(13), CEB => n166, CK 
                           => clk, RB => resetn, Q => in_buf_189_port);
   in_buf_reg_2_27 : DFERPQ1 port map( D => siso_data_in(11), CEB => n166, CK 
                           => clk, RB => resetn, Q => in_buf_187_port);
   in_buf_reg_2_25 : DFERPQ1 port map( D => siso_data_in(9), CEB => n166, CK =>
                           clk, RB => resetn, Q => in_buf_185_port);
   in_buf_reg_2_23 : DFERPQ1 port map( D => siso_data_in(7), CEB => n166, CK =>
                           clk, RB => resetn, Q => in_buf_183_port);
   in_buf_reg_2_21 : DFERPQ1 port map( D => siso_data_in(5), CEB => n166, CK =>
                           clk, RB => resetn, Q => in_buf_181_port);
   in_buf_reg_2_19 : DFERPQ1 port map( D => siso_data_in(3), CEB => n166, CK =>
                           clk, RB => resetn, Q => in_buf_179_port);
   in_buf_reg_2_17 : DFERPQ1 port map( D => siso_data_in(1), CEB => n166, CK =>
                           clk, RB => resetn, Q => in_buf_177_port);
   in_buf_reg_6_31 : DFERPQ1 port map( D => siso_data_in(15), CEB => n174, CK 
                           => clk, RB => resetn, Q => in_buf_63_port);
   in_buf_reg_6_29 : DFERPQ1 port map( D => siso_data_in(13), CEB => n174, CK 
                           => clk, RB => resetn, Q => in_buf_61_port);
   in_buf_reg_6_27 : DFERPQ1 port map( D => siso_data_in(11), CEB => n174, CK 
                           => clk, RB => resetn, Q => in_buf_59_port);
   in_buf_reg_6_25 : DFERPQ1 port map( D => siso_data_in(9), CEB => n174, CK =>
                           clk, RB => resetn, Q => in_buf_57_port);
   in_buf_reg_6_23 : DFERPQ1 port map( D => siso_data_in(7), CEB => n174, CK =>
                           clk, RB => resetn, Q => in_buf_55_port);
   in_buf_reg_6_21 : DFERPQ1 port map( D => siso_data_in(5), CEB => n174, CK =>
                           clk, RB => resetn, Q => in_buf_53_port);
   in_buf_reg_6_19 : DFERPQ1 port map( D => siso_data_in(3), CEB => n174, CK =>
                           clk, RB => resetn, Q => in_buf_51_port);
   in_buf_reg_6_17 : DFERPQ1 port map( D => siso_data_in(1), CEB => n174, CK =>
                           clk, RB => resetn, Q => in_buf_49_port);
   in_buf_reg_2_15 : DFERPQ1 port map( D => siso_data_in(15), CEB => n167, CK 
                           => clk, RB => resetn, Q => in_buf_175_port);
   in_buf_reg_2_13 : DFERPQ1 port map( D => siso_data_in(13), CEB => n167, CK 
                           => clk, RB => resetn, Q => in_buf_173_port);
   in_buf_reg_2_11 : DFERPQ1 port map( D => siso_data_in(11), CEB => n167, CK 
                           => clk, RB => resetn, Q => in_buf_171_port);
   in_buf_reg_2_9 : DFERPQ1 port map( D => siso_data_in(9), CEB => n167, CK => 
                           clk, RB => resetn, Q => in_buf_169_port);
   in_buf_reg_2_7 : DFERPQ1 port map( D => siso_data_in(7), CEB => n167, CK => 
                           clk, RB => resetn, Q => in_buf_167_port);
   in_buf_reg_2_5 : DFERPQ1 port map( D => siso_data_in(5), CEB => n167, CK => 
                           clk, RB => resetn, Q => in_buf_165_port);
   in_buf_reg_2_3 : DFERPQ1 port map( D => siso_data_in(3), CEB => n167, CK => 
                           clk, RB => resetn, Q => in_buf_163_port);
   in_buf_reg_2_1 : DFERPQ1 port map( D => siso_data_in(1), CEB => n167, CK => 
                           clk, RB => resetn, Q => in_buf_161_port);
   in_buf_reg_6_15 : DFERPQ1 port map( D => siso_data_in(15), CEB => n175, CK 
                           => clk, RB => resetn, Q => in_buf_47_port);
   in_buf_reg_6_13 : DFERPQ1 port map( D => siso_data_in(13), CEB => n175, CK 
                           => clk, RB => resetn, Q => in_buf_45_port);
   in_buf_reg_6_11 : DFERPQ1 port map( D => siso_data_in(11), CEB => n175, CK 
                           => clk, RB => resetn, Q => in_buf_43_port);
   in_buf_reg_6_9 : DFERPQ1 port map( D => siso_data_in(9), CEB => n175, CK => 
                           clk, RB => resetn, Q => in_buf_41_port);
   in_buf_reg_6_7 : DFERPQ1 port map( D => siso_data_in(7), CEB => n175, CK => 
                           clk, RB => resetn, Q => in_buf_39_port);
   in_buf_reg_6_5 : DFERPQ1 port map( D => siso_data_in(5), CEB => n175, CK => 
                           clk, RB => resetn, Q => in_buf_37_port);
   in_buf_reg_6_3 : DFERPQ1 port map( D => siso_data_in(3), CEB => n175, CK => 
                           clk, RB => resetn, Q => in_buf_35_port);
   in_buf_reg_6_1 : DFERPQ1 port map( D => siso_data_in(1), CEB => n175, CK => 
                           clk, RB => resetn, Q => in_buf_33_port);
   in_buf_reg_5_31 : DFERPQ1 port map( D => siso_data_in(15), CEB => n172, CK 
                           => clk, RB => resetn, Q => in_buf_95_port);
   in_buf_reg_5_29 : DFERPQ1 port map( D => siso_data_in(13), CEB => n172, CK 
                           => clk, RB => resetn, Q => in_buf_93_port);
   in_buf_reg_5_27 : DFERPQ1 port map( D => siso_data_in(11), CEB => n172, CK 
                           => clk, RB => resetn, Q => in_buf_91_port);
   in_buf_reg_5_25 : DFERPQ1 port map( D => siso_data_in(9), CEB => n172, CK =>
                           clk, RB => resetn, Q => in_buf_89_port);
   in_buf_reg_5_23 : DFERPQ1 port map( D => siso_data_in(7), CEB => n172, CK =>
                           clk, RB => resetn, Q => in_buf_87_port);
   in_buf_reg_5_21 : DFERPQ1 port map( D => siso_data_in(5), CEB => n172, CK =>
                           clk, RB => resetn, Q => in_buf_85_port);
   in_buf_reg_5_19 : DFERPQ1 port map( D => siso_data_in(3), CEB => n172, CK =>
                           clk, RB => resetn, Q => in_buf_83_port);
   in_buf_reg_5_17 : DFERPQ1 port map( D => siso_data_in(1), CEB => n172, CK =>
                           clk, RB => resetn, Q => in_buf_81_port);
   in_buf_reg_5_15 : DFERPQ1 port map( D => siso_data_in(15), CEB => n173, CK 
                           => clk, RB => resetn, Q => in_buf_79_port);
   in_buf_reg_5_13 : DFERPQ1 port map( D => siso_data_in(13), CEB => n173, CK 
                           => clk, RB => resetn, Q => in_buf_77_port);
   in_buf_reg_5_11 : DFERPQ1 port map( D => siso_data_in(11), CEB => n173, CK 
                           => clk, RB => resetn, Q => in_buf_75_port);
   in_buf_reg_5_9 : DFERPQ1 port map( D => siso_data_in(9), CEB => n173, CK => 
                           clk, RB => resetn, Q => in_buf_73_port);
   in_buf_reg_5_7 : DFERPQ1 port map( D => siso_data_in(7), CEB => n173, CK => 
                           clk, RB => resetn, Q => in_buf_71_port);
   in_buf_reg_5_5 : DFERPQ1 port map( D => siso_data_in(5), CEB => n173, CK => 
                           clk, RB => resetn, Q => in_buf_69_port);
   in_buf_reg_5_3 : DFERPQ1 port map( D => siso_data_in(3), CEB => n173, CK => 
                           clk, RB => resetn, Q => in_buf_67_port);
   in_buf_reg_5_1 : DFERPQ1 port map( D => siso_data_in(1), CEB => n173, CK => 
                           clk, RB => resetn, Q => in_buf_65_port);
   comp_res_reg_1_31 : DFFRPQ1 port map( D => N3296, CK => clk, RB => resetn, Q
                           => comp_res_127_port);
   comp_res_reg_1_29 : DFFRPQ1 port map( D => N3294, CK => clk, RB => resetn, Q
                           => comp_res_125_port);
   comp_res_reg_1_27 : DFFRPQ1 port map( D => N3292, CK => clk, RB => resetn, Q
                           => comp_res_123_port);
   comp_res_reg_1_25 : DFFRPQ1 port map( D => N3290, CK => clk, RB => resetn, Q
                           => comp_res_121_port);
   comp_res_reg_1_23 : DFFRPQ1 port map( D => N3288, CK => clk, RB => resetn, Q
                           => comp_res_119_port);
   comp_res_reg_1_21 : DFFRPQ1 port map( D => N3286, CK => clk, RB => resetn, Q
                           => comp_res_117_port);
   comp_res_reg_1_19 : DFFRPQ1 port map( D => N3284, CK => clk, RB => resetn, Q
                           => comp_res_115_port);
   comp_res_reg_1_17 : DFFRPQ1 port map( D => N3282, CK => clk, RB => resetn, Q
                           => comp_res_113_port);
   comp_res_reg_1_15 : DFFRPQ1 port map( D => N3280, CK => clk, RB => resetn, Q
                           => comp_res_111_port);
   comp_res_reg_1_13 : DFFRPQ1 port map( D => N3278, CK => clk, RB => resetn, Q
                           => comp_res_109_port);
   comp_res_reg_1_11 : DFFRPQ1 port map( D => N3276, CK => clk, RB => resetn, Q
                           => comp_res_107_port);
   comp_res_reg_1_9 : DFFRPQ1 port map( D => N3274, CK => clk, RB => resetn, Q 
                           => comp_res_105_port);
   comp_res_reg_1_7 : DFFRPQ1 port map( D => N3272, CK => clk, RB => resetn, Q 
                           => comp_res_103_port);
   comp_res_reg_1_5 : DFFRPQ1 port map( D => N3270, CK => clk, RB => resetn, Q 
                           => comp_res_101_port);
   comp_res_reg_1_3 : DFFRPQ1 port map( D => N3268, CK => clk, RB => resetn, Q 
                           => comp_res_99_port);
   comp_res_reg_1_1 : DFFRPQ1 port map( D => N3266, CK => clk, RB => resetn, Q 
                           => comp_res_97_port);
   comp_res_reg_0_31 : DFFRPQ1 port map( D => N3264, CK => clk, RB => resetn, Q
                           => comp_res_159_port);
   comp_res_reg_0_29 : DFFRPQ1 port map( D => N3262, CK => clk, RB => resetn, Q
                           => comp_res_157_port);
   comp_res_reg_0_27 : DFFRPQ1 port map( D => N3260, CK => clk, RB => resetn, Q
                           => comp_res_155_port);
   comp_res_reg_0_25 : DFFRPQ1 port map( D => N3258, CK => clk, RB => resetn, Q
                           => comp_res_153_port);
   comp_res_reg_0_23 : DFFRPQ1 port map( D => N3256, CK => clk, RB => resetn, Q
                           => comp_res_151_port);
   comp_res_reg_0_21 : DFFRPQ1 port map( D => N3254, CK => clk, RB => resetn, Q
                           => comp_res_149_port);
   comp_res_reg_0_19 : DFFRPQ1 port map( D => N3252, CK => clk, RB => resetn, Q
                           => comp_res_147_port);
   comp_res_reg_0_17 : DFFRPQ1 port map( D => N3250, CK => clk, RB => resetn, Q
                           => comp_res_145_port);
   comp_res_reg_0_15 : DFFRPQ1 port map( D => N3248, CK => clk, RB => resetn, Q
                           => comp_res_143_port);
   comp_res_reg_0_13 : DFFRPQ1 port map( D => N3246, CK => clk, RB => resetn, Q
                           => comp_res_141_port);
   comp_res_reg_0_11 : DFFRPQ1 port map( D => N3244, CK => clk, RB => resetn, Q
                           => comp_res_139_port);
   comp_res_reg_0_9 : DFFRPQ1 port map( D => N3242, CK => clk, RB => resetn, Q 
                           => comp_res_137_port);
   comp_res_reg_0_7 : DFFRPQ1 port map( D => N3240, CK => clk, RB => resetn, Q 
                           => comp_res_135_port);
   comp_res_reg_0_5 : DFFRPQ1 port map( D => N3238, CK => clk, RB => resetn, Q 
                           => comp_res_133_port);
   comp_res_reg_0_3 : DFFRPQ1 port map( D => N3236, CK => clk, RB => resetn, Q 
                           => comp_res_131_port);
   comp_res_reg_0_1 : DFFRPQ1 port map( D => N3234, CK => clk, RB => resetn, Q 
                           => comp_res_129_port);
   in_buf_reg_1_31 : DFERPQ1 port map( D => siso_data_in(15), CEB => n164, CK 
                           => clk, RB => resetn, Q => in_buf_223_port);
   in_buf_reg_1_29 : DFERPQ1 port map( D => siso_data_in(13), CEB => n164, CK 
                           => clk, RB => resetn, Q => in_buf_221_port);
   in_buf_reg_1_27 : DFERPQ1 port map( D => siso_data_in(11), CEB => n164, CK 
                           => clk, RB => resetn, Q => in_buf_219_port);
   in_buf_reg_1_25 : DFERPQ1 port map( D => siso_data_in(9), CEB => n164, CK =>
                           clk, RB => resetn, Q => in_buf_217_port);
   in_buf_reg_1_23 : DFERPQ1 port map( D => siso_data_in(7), CEB => n164, CK =>
                           clk, RB => resetn, Q => in_buf_215_port);
   in_buf_reg_1_21 : DFERPQ1 port map( D => siso_data_in(5), CEB => n164, CK =>
                           clk, RB => resetn, Q => in_buf_213_port);
   in_buf_reg_1_19 : DFERPQ1 port map( D => siso_data_in(3), CEB => n164, CK =>
                           clk, RB => resetn, Q => in_buf_211_port);
   in_buf_reg_1_17 : DFERPQ1 port map( D => siso_data_in(1), CEB => n164, CK =>
                           clk, RB => resetn, Q => in_buf_209_port);
   in_buf_reg_1_15 : DFERPQ1 port map( D => siso_data_in(15), CEB => n165, CK 
                           => clk, RB => resetn, Q => in_buf_207_port);
   in_buf_reg_1_13 : DFERPQ1 port map( D => siso_data_in(13), CEB => n165, CK 
                           => clk, RB => resetn, Q => in_buf_205_port);
   in_buf_reg_1_11 : DFERPQ1 port map( D => siso_data_in(11), CEB => n165, CK 
                           => clk, RB => resetn, Q => in_buf_203_port);
   in_buf_reg_1_9 : DFERPQ1 port map( D => siso_data_in(9), CEB => n165, CK => 
                           clk, RB => resetn, Q => in_buf_201_port);
   in_buf_reg_1_7 : DFERPQ1 port map( D => siso_data_in(7), CEB => n165, CK => 
                           clk, RB => resetn, Q => in_buf_199_port);
   in_buf_reg_1_5 : DFERPQ1 port map( D => siso_data_in(5), CEB => n165, CK => 
                           clk, RB => resetn, Q => in_buf_197_port);
   in_buf_reg_1_3 : DFERPQ1 port map( D => siso_data_in(3), CEB => n165, CK => 
                           clk, RB => resetn, Q => in_buf_195_port);
   in_buf_reg_1_1 : DFERPQ1 port map( D => siso_data_in(1), CEB => n165, CK => 
                           clk, RB => resetn, Q => in_buf_193_port);
   in_buf_reg_4_31 : DFERPQ1 port map( D => siso_data_in(15), CEB => n170, CK 
                           => clk, RB => resetn, Q => in_buf_127_port);
   in_buf_reg_4_29 : DFERPQ1 port map( D => siso_data_in(13), CEB => n170, CK 
                           => clk, RB => resetn, Q => in_buf_125_port);
   in_buf_reg_4_27 : DFERPQ1 port map( D => siso_data_in(11), CEB => n170, CK 
                           => clk, RB => resetn, Q => in_buf_123_port);
   in_buf_reg_4_25 : DFERPQ1 port map( D => siso_data_in(9), CEB => n170, CK =>
                           clk, RB => resetn, Q => in_buf_121_port);
   in_buf_reg_4_23 : DFERPQ1 port map( D => siso_data_in(7), CEB => n170, CK =>
                           clk, RB => resetn, Q => in_buf_119_port);
   in_buf_reg_4_21 : DFERPQ1 port map( D => siso_data_in(5), CEB => n170, CK =>
                           clk, RB => resetn, Q => in_buf_117_port);
   in_buf_reg_4_19 : DFERPQ1 port map( D => siso_data_in(3), CEB => n170, CK =>
                           clk, RB => resetn, Q => in_buf_115_port);
   in_buf_reg_4_17 : DFERPQ1 port map( D => siso_data_in(1), CEB => n170, CK =>
                           clk, RB => resetn, Q => in_buf_113_port);
   in_buf_reg_0_31 : DFERPQ1 port map( D => siso_data_in(15), CEB => n162, CK 
                           => clk, RB => resetn, Q => in_buf_255_port);
   in_buf_reg_0_29 : DFERPQ1 port map( D => siso_data_in(13), CEB => n162, CK 
                           => clk, RB => resetn, Q => in_buf_253_port);
   in_buf_reg_0_27 : DFERPQ1 port map( D => siso_data_in(11), CEB => n162, CK 
                           => clk, RB => resetn, Q => in_buf_251_port);
   in_buf_reg_0_25 : DFERPQ1 port map( D => siso_data_in(9), CEB => n162, CK =>
                           clk, RB => resetn, Q => in_buf_249_port);
   in_buf_reg_0_23 : DFERPQ1 port map( D => siso_data_in(7), CEB => n162, CK =>
                           clk, RB => resetn, Q => in_buf_247_port);
   in_buf_reg_0_21 : DFERPQ1 port map( D => siso_data_in(5), CEB => n162, CK =>
                           clk, RB => resetn, Q => in_buf_245_port);
   in_buf_reg_0_19 : DFERPQ1 port map( D => siso_data_in(3), CEB => n162, CK =>
                           clk, RB => resetn, Q => in_buf_243_port);
   in_buf_reg_0_17 : DFERPQ1 port map( D => siso_data_in(1), CEB => n162, CK =>
                           clk, RB => resetn, Q => in_buf_241_port);
   in_buf_reg_0_15 : DFERPQ1 port map( D => siso_data_in(15), CEB => n163, CK 
                           => clk, RB => resetn, Q => in_buf_239_port);
   in_buf_reg_0_13 : DFERPQ1 port map( D => siso_data_in(13), CEB => n163, CK 
                           => clk, RB => resetn, Q => in_buf_237_port);
   in_buf_reg_0_11 : DFERPQ1 port map( D => siso_data_in(11), CEB => n163, CK 
                           => clk, RB => resetn, Q => in_buf_235_port);
   in_buf_reg_0_9 : DFERPQ1 port map( D => siso_data_in(9), CEB => n163, CK => 
                           clk, RB => resetn, Q => in_buf_233_port);
   in_buf_reg_0_7 : DFERPQ1 port map( D => siso_data_in(7), CEB => n163, CK => 
                           clk, RB => resetn, Q => in_buf_231_port);
   in_buf_reg_0_5 : DFERPQ1 port map( D => siso_data_in(5), CEB => n163, CK => 
                           clk, RB => resetn, Q => in_buf_229_port);
   in_buf_reg_0_3 : DFERPQ1 port map( D => siso_data_in(3), CEB => n163, CK => 
                           clk, RB => resetn, Q => in_buf_227_port);
   in_buf_reg_0_1 : DFERPQ1 port map( D => siso_data_in(1), CEB => n163, CK => 
                           clk, RB => resetn, Q => in_buf_225_port);
   in_buf_reg_4_15 : DFERPQ1 port map( D => siso_data_in(15), CEB => n171, CK 
                           => clk, RB => resetn, Q => in_buf_111_port);
   in_buf_reg_4_13 : DFERPQ1 port map( D => siso_data_in(13), CEB => n171, CK 
                           => clk, RB => resetn, Q => in_buf_109_port);
   in_buf_reg_4_11 : DFERPQ1 port map( D => siso_data_in(11), CEB => n171, CK 
                           => clk, RB => resetn, Q => in_buf_107_port);
   in_buf_reg_4_9 : DFERPQ1 port map( D => siso_data_in(9), CEB => n171, CK => 
                           clk, RB => resetn, Q => in_buf_105_port);
   in_buf_reg_4_7 : DFERPQ1 port map( D => siso_data_in(7), CEB => n171, CK => 
                           clk, RB => resetn, Q => in_buf_103_port);
   in_buf_reg_4_5 : DFERPQ1 port map( D => siso_data_in(5), CEB => n171, CK => 
                           clk, RB => resetn, Q => in_buf_101_port);
   in_buf_reg_4_3 : DFERPQ1 port map( D => siso_data_in(3), CEB => n171, CK => 
                           clk, RB => resetn, Q => in_buf_99_port);
   in_buf_reg_4_1 : DFERPQ1 port map( D => siso_data_in(1), CEB => n171, CK => 
                           clk, RB => resetn, Q => in_buf_97_port);
   in_buf_reg_7_30 : DFERPQ1 port map( D => siso_data_in(14), CEB => n176, CK 
                           => clk, RB => resetn, Q => in_buf_30_port);
   in_buf_reg_7_28 : DFERPQ1 port map( D => siso_data_in(12), CEB => n176, CK 
                           => clk, RB => resetn, Q => in_buf_28_port);
   in_buf_reg_7_26 : DFERPQ1 port map( D => siso_data_in(10), CEB => n176, CK 
                           => clk, RB => resetn, Q => in_buf_26_port);
   in_buf_reg_7_24 : DFERPQ1 port map( D => siso_data_in(8), CEB => n176, CK =>
                           clk, RB => resetn, Q => in_buf_24_port);
   in_buf_reg_7_22 : DFERPQ1 port map( D => siso_data_in(6), CEB => n176, CK =>
                           clk, RB => resetn, Q => in_buf_22_port);
   in_buf_reg_7_20 : DFERPQ1 port map( D => siso_data_in(4), CEB => n176, CK =>
                           clk, RB => resetn, Q => in_buf_20_port);
   in_buf_reg_7_18 : DFERPQ1 port map( D => siso_data_in(2), CEB => n176, CK =>
                           clk, RB => resetn, Q => in_buf_18_port);
   in_buf_reg_7_16 : DFERPQ1 port map( D => siso_data_in(0), CEB => n176, CK =>
                           clk, RB => resetn, Q => in_buf_16_port);
   in_buf_reg_7_14 : DFERPQ1 port map( D => siso_data_in(14), CEB => n177, CK 
                           => clk, RB => resetn, Q => in_buf_14_port);
   in_buf_reg_7_12 : DFERPQ1 port map( D => siso_data_in(12), CEB => n177, CK 
                           => clk, RB => resetn, Q => in_buf_12_port);
   in_buf_reg_7_10 : DFERPQ1 port map( D => siso_data_in(10), CEB => n177, CK 
                           => clk, RB => resetn, Q => in_buf_10_port);
   in_buf_reg_7_8 : DFERPQ1 port map( D => siso_data_in(8), CEB => n177, CK => 
                           clk, RB => resetn, Q => in_buf_8_port);
   in_buf_reg_7_6 : DFERPQ1 port map( D => siso_data_in(6), CEB => n177, CK => 
                           clk, RB => resetn, Q => in_buf_6_port);
   in_buf_reg_7_4 : DFERPQ1 port map( D => siso_data_in(4), CEB => n177, CK => 
                           clk, RB => resetn, Q => in_buf_4_port);
   in_buf_reg_7_2 : DFERPQ1 port map( D => siso_data_in(2), CEB => n177, CK => 
                           clk, RB => resetn, Q => in_buf_2_port);
   in_trigger_reg : DFFRPQ1 port map( D => n241, CK => clk, RB => resetn, Q => 
                           in_trigger);
   in_buf_reg_3_30 : DFERPQ1 port map( D => siso_data_in(14), CEB => n168, CK 
                           => clk, RB => resetn, Q => in_buf_158_port);
   in_buf_reg_3_28 : DFERPQ1 port map( D => siso_data_in(12), CEB => n168, CK 
                           => clk, RB => resetn, Q => in_buf_156_port);
   in_buf_reg_3_26 : DFERPQ1 port map( D => siso_data_in(10), CEB => n168, CK 
                           => clk, RB => resetn, Q => in_buf_154_port);
   in_buf_reg_3_24 : DFERPQ1 port map( D => siso_data_in(8), CEB => n168, CK =>
                           clk, RB => resetn, Q => in_buf_152_port);
   in_buf_reg_3_22 : DFERPQ1 port map( D => siso_data_in(6), CEB => n168, CK =>
                           clk, RB => resetn, Q => in_buf_150_port);
   in_buf_reg_3_20 : DFERPQ1 port map( D => siso_data_in(4), CEB => n168, CK =>
                           clk, RB => resetn, Q => in_buf_148_port);
   in_buf_reg_3_18 : DFERPQ1 port map( D => siso_data_in(2), CEB => n168, CK =>
                           clk, RB => resetn, Q => in_buf_146_port);
   in_buf_reg_3_16 : DFERPQ1 port map( D => siso_data_in(0), CEB => n168, CK =>
                           clk, RB => resetn, Q => in_buf_144_port);
   in_buf_reg_3_14 : DFERPQ1 port map( D => siso_data_in(14), CEB => n169, CK 
                           => clk, RB => resetn, Q => in_buf_142_port);
   in_buf_reg_3_12 : DFERPQ1 port map( D => siso_data_in(12), CEB => n169, CK 
                           => clk, RB => resetn, Q => in_buf_140_port);
   in_buf_reg_3_10 : DFERPQ1 port map( D => siso_data_in(10), CEB => n169, CK 
                           => clk, RB => resetn, Q => in_buf_138_port);
   in_buf_reg_3_8 : DFERPQ1 port map( D => siso_data_in(8), CEB => n169, CK => 
                           clk, RB => resetn, Q => in_buf_136_port);
   in_buf_reg_3_6 : DFERPQ1 port map( D => siso_data_in(6), CEB => n169, CK => 
                           clk, RB => resetn, Q => in_buf_134_port);
   in_buf_reg_3_4 : DFERPQ1 port map( D => siso_data_in(4), CEB => n169, CK => 
                           clk, RB => resetn, Q => in_buf_132_port);
   in_buf_reg_3_2 : DFERPQ1 port map( D => siso_data_in(2), CEB => n169, CK => 
                           clk, RB => resetn, Q => in_buf_130_port);
   in_buf_reg_2_30 : DFERPQ1 port map( D => siso_data_in(14), CEB => n166, CK 
                           => clk, RB => resetn, Q => in_buf_190_port);
   in_buf_reg_2_28 : DFERPQ1 port map( D => siso_data_in(12), CEB => n166, CK 
                           => clk, RB => resetn, Q => in_buf_188_port);
   in_buf_reg_2_26 : DFERPQ1 port map( D => siso_data_in(10), CEB => n166, CK 
                           => clk, RB => resetn, Q => in_buf_186_port);
   in_buf_reg_2_24 : DFERPQ1 port map( D => siso_data_in(8), CEB => n166, CK =>
                           clk, RB => resetn, Q => in_buf_184_port);
   in_buf_reg_2_22 : DFERPQ1 port map( D => siso_data_in(6), CEB => n166, CK =>
                           clk, RB => resetn, Q => in_buf_182_port);
   in_buf_reg_2_20 : DFERPQ1 port map( D => siso_data_in(4), CEB => n166, CK =>
                           clk, RB => resetn, Q => in_buf_180_port);
   in_buf_reg_2_18 : DFERPQ1 port map( D => siso_data_in(2), CEB => n166, CK =>
                           clk, RB => resetn, Q => in_buf_178_port);
   in_buf_reg_2_16 : DFERPQ1 port map( D => siso_data_in(0), CEB => n166, CK =>
                           clk, RB => resetn, Q => in_buf_176_port);
   in_buf_reg_6_30 : DFERPQ1 port map( D => siso_data_in(14), CEB => n174, CK 
                           => clk, RB => resetn, Q => in_buf_62_port);
   in_buf_reg_6_28 : DFERPQ1 port map( D => siso_data_in(12), CEB => n174, CK 
                           => clk, RB => resetn, Q => in_buf_60_port);
   in_buf_reg_6_26 : DFERPQ1 port map( D => siso_data_in(10), CEB => n174, CK 
                           => clk, RB => resetn, Q => in_buf_58_port);
   in_buf_reg_6_24 : DFERPQ1 port map( D => siso_data_in(8), CEB => n174, CK =>
                           clk, RB => resetn, Q => in_buf_56_port);
   in_buf_reg_6_22 : DFERPQ1 port map( D => siso_data_in(6), CEB => n174, CK =>
                           clk, RB => resetn, Q => in_buf_54_port);
   in_buf_reg_6_20 : DFERPQ1 port map( D => siso_data_in(4), CEB => n174, CK =>
                           clk, RB => resetn, Q => in_buf_52_port);
   in_buf_reg_6_18 : DFERPQ1 port map( D => siso_data_in(2), CEB => n174, CK =>
                           clk, RB => resetn, Q => in_buf_50_port);
   in_buf_reg_6_16 : DFERPQ1 port map( D => siso_data_in(0), CEB => n174, CK =>
                           clk, RB => resetn, Q => in_buf_48_port);
   in_buf_reg_2_14 : DFERPQ1 port map( D => siso_data_in(14), CEB => n167, CK 
                           => clk, RB => resetn, Q => in_buf_174_port);
   in_buf_reg_2_12 : DFERPQ1 port map( D => siso_data_in(12), CEB => n167, CK 
                           => clk, RB => resetn, Q => in_buf_172_port);
   in_buf_reg_2_10 : DFERPQ1 port map( D => siso_data_in(10), CEB => n167, CK 
                           => clk, RB => resetn, Q => in_buf_170_port);
   in_buf_reg_2_8 : DFERPQ1 port map( D => siso_data_in(8), CEB => n167, CK => 
                           clk, RB => resetn, Q => in_buf_168_port);
   in_buf_reg_2_6 : DFERPQ1 port map( D => siso_data_in(6), CEB => n167, CK => 
                           clk, RB => resetn, Q => in_buf_166_port);
   in_buf_reg_2_4 : DFERPQ1 port map( D => siso_data_in(4), CEB => n167, CK => 
                           clk, RB => resetn, Q => in_buf_164_port);
   in_buf_reg_2_2 : DFERPQ1 port map( D => siso_data_in(2), CEB => n167, CK => 
                           clk, RB => resetn, Q => in_buf_162_port);
   in_buf_reg_6_14 : DFERPQ1 port map( D => siso_data_in(14), CEB => n175, CK 
                           => clk, RB => resetn, Q => in_buf_46_port);
   in_buf_reg_6_12 : DFERPQ1 port map( D => siso_data_in(12), CEB => n175, CK 
                           => clk, RB => resetn, Q => in_buf_44_port);
   in_buf_reg_6_10 : DFERPQ1 port map( D => siso_data_in(10), CEB => n175, CK 
                           => clk, RB => resetn, Q => in_buf_42_port);
   in_buf_reg_6_8 : DFERPQ1 port map( D => siso_data_in(8), CEB => n175, CK => 
                           clk, RB => resetn, Q => in_buf_40_port);
   in_buf_reg_6_6 : DFERPQ1 port map( D => siso_data_in(6), CEB => n175, CK => 
                           clk, RB => resetn, Q => in_buf_38_port);
   in_buf_reg_6_4 : DFERPQ1 port map( D => siso_data_in(4), CEB => n175, CK => 
                           clk, RB => resetn, Q => in_buf_36_port);
   in_buf_reg_6_2 : DFERPQ1 port map( D => siso_data_in(2), CEB => n175, CK => 
                           clk, RB => resetn, Q => in_buf_34_port);
   in_buf_reg_5_30 : DFERPQ1 port map( D => siso_data_in(14), CEB => n172, CK 
                           => clk, RB => resetn, Q => in_buf_94_port);
   in_buf_reg_5_28 : DFERPQ1 port map( D => siso_data_in(12), CEB => n172, CK 
                           => clk, RB => resetn, Q => in_buf_92_port);
   in_buf_reg_5_26 : DFERPQ1 port map( D => siso_data_in(10), CEB => n172, CK 
                           => clk, RB => resetn, Q => in_buf_90_port);
   in_buf_reg_5_24 : DFERPQ1 port map( D => siso_data_in(8), CEB => n172, CK =>
                           clk, RB => resetn, Q => in_buf_88_port);
   in_buf_reg_5_22 : DFERPQ1 port map( D => siso_data_in(6), CEB => n172, CK =>
                           clk, RB => resetn, Q => in_buf_86_port);
   in_buf_reg_5_20 : DFERPQ1 port map( D => siso_data_in(4), CEB => n172, CK =>
                           clk, RB => resetn, Q => in_buf_84_port);
   in_buf_reg_5_18 : DFERPQ1 port map( D => siso_data_in(2), CEB => n172, CK =>
                           clk, RB => resetn, Q => in_buf_82_port);
   in_buf_reg_5_16 : DFERPQ1 port map( D => siso_data_in(0), CEB => n172, CK =>
                           clk, RB => resetn, Q => in_buf_80_port);
   in_buf_reg_5_14 : DFERPQ1 port map( D => siso_data_in(14), CEB => n173, CK 
                           => clk, RB => resetn, Q => in_buf_78_port);
   in_buf_reg_5_12 : DFERPQ1 port map( D => siso_data_in(12), CEB => n173, CK 
                           => clk, RB => resetn, Q => in_buf_76_port);
   in_buf_reg_5_10 : DFERPQ1 port map( D => siso_data_in(10), CEB => n173, CK 
                           => clk, RB => resetn, Q => in_buf_74_port);
   in_buf_reg_5_8 : DFERPQ1 port map( D => siso_data_in(8), CEB => n173, CK => 
                           clk, RB => resetn, Q => in_buf_72_port);
   in_buf_reg_5_6 : DFERPQ1 port map( D => siso_data_in(6), CEB => n173, CK => 
                           clk, RB => resetn, Q => in_buf_70_port);
   in_buf_reg_5_4 : DFERPQ1 port map( D => siso_data_in(4), CEB => n173, CK => 
                           clk, RB => resetn, Q => in_buf_68_port);
   in_buf_reg_5_2 : DFERPQ1 port map( D => siso_data_in(2), CEB => n173, CK => 
                           clk, RB => resetn, Q => in_buf_66_port);
   in_buf_reg_7_0 : DFERPQ1 port map( D => siso_data_in(0), CEB => n177, CK => 
                           clk, RB => resetn, Q => in_buf_0_port);
   in_buf_reg_1_30 : DFERPQ1 port map( D => siso_data_in(14), CEB => n164, CK 
                           => clk, RB => resetn, Q => in_buf_222_port);
   in_buf_reg_1_28 : DFERPQ1 port map( D => siso_data_in(12), CEB => n164, CK 
                           => clk, RB => resetn, Q => in_buf_220_port);
   in_buf_reg_1_26 : DFERPQ1 port map( D => siso_data_in(10), CEB => n164, CK 
                           => clk, RB => resetn, Q => in_buf_218_port);
   in_buf_reg_1_24 : DFERPQ1 port map( D => siso_data_in(8), CEB => n164, CK =>
                           clk, RB => resetn, Q => in_buf_216_port);
   in_buf_reg_1_22 : DFERPQ1 port map( D => siso_data_in(6), CEB => n164, CK =>
                           clk, RB => resetn, Q => in_buf_214_port);
   in_buf_reg_1_20 : DFERPQ1 port map( D => siso_data_in(4), CEB => n164, CK =>
                           clk, RB => resetn, Q => in_buf_212_port);
   in_buf_reg_1_18 : DFERPQ1 port map( D => siso_data_in(2), CEB => n164, CK =>
                           clk, RB => resetn, Q => in_buf_210_port);
   in_buf_reg_1_16 : DFERPQ1 port map( D => siso_data_in(0), CEB => n164, CK =>
                           clk, RB => resetn, Q => in_buf_208_port);
   in_buf_reg_1_14 : DFERPQ1 port map( D => siso_data_in(14), CEB => n165, CK 
                           => clk, RB => resetn, Q => in_buf_206_port);
   in_buf_reg_1_12 : DFERPQ1 port map( D => siso_data_in(12), CEB => n165, CK 
                           => clk, RB => resetn, Q => in_buf_204_port);
   in_buf_reg_1_10 : DFERPQ1 port map( D => siso_data_in(10), CEB => n165, CK 
                           => clk, RB => resetn, Q => in_buf_202_port);
   in_buf_reg_1_8 : DFERPQ1 port map( D => siso_data_in(8), CEB => n165, CK => 
                           clk, RB => resetn, Q => in_buf_200_port);
   in_buf_reg_1_6 : DFERPQ1 port map( D => siso_data_in(6), CEB => n165, CK => 
                           clk, RB => resetn, Q => in_buf_198_port);
   in_buf_reg_1_4 : DFERPQ1 port map( D => siso_data_in(4), CEB => n165, CK => 
                           clk, RB => resetn, Q => in_buf_196_port);
   in_buf_reg_1_2 : DFERPQ1 port map( D => siso_data_in(2), CEB => n165, CK => 
                           clk, RB => resetn, Q => in_buf_194_port);
   in_buf_reg_4_30 : DFERPQ1 port map( D => siso_data_in(14), CEB => n170, CK 
                           => clk, RB => resetn, Q => in_buf_126_port);
   in_buf_reg_4_28 : DFERPQ1 port map( D => siso_data_in(12), CEB => n170, CK 
                           => clk, RB => resetn, Q => in_buf_124_port);
   in_buf_reg_4_26 : DFERPQ1 port map( D => siso_data_in(10), CEB => n170, CK 
                           => clk, RB => resetn, Q => in_buf_122_port);
   in_buf_reg_4_24 : DFERPQ1 port map( D => siso_data_in(8), CEB => n170, CK =>
                           clk, RB => resetn, Q => in_buf_120_port);
   in_buf_reg_4_22 : DFERPQ1 port map( D => siso_data_in(6), CEB => n170, CK =>
                           clk, RB => resetn, Q => in_buf_118_port);
   in_buf_reg_4_20 : DFERPQ1 port map( D => siso_data_in(4), CEB => n170, CK =>
                           clk, RB => resetn, Q => in_buf_116_port);
   in_buf_reg_4_18 : DFERPQ1 port map( D => siso_data_in(2), CEB => n170, CK =>
                           clk, RB => resetn, Q => in_buf_114_port);
   in_buf_reg_4_16 : DFERPQ1 port map( D => siso_data_in(0), CEB => n170, CK =>
                           clk, RB => resetn, Q => in_buf_112_port);
   in_buf_reg_0_30 : DFERPQ1 port map( D => siso_data_in(14), CEB => n162, CK 
                           => clk, RB => resetn, Q => in_buf_254_port);
   in_buf_reg_0_28 : DFERPQ1 port map( D => siso_data_in(12), CEB => n162, CK 
                           => clk, RB => resetn, Q => in_buf_252_port);
   in_buf_reg_0_26 : DFERPQ1 port map( D => siso_data_in(10), CEB => n162, CK 
                           => clk, RB => resetn, Q => in_buf_250_port);
   in_buf_reg_0_24 : DFERPQ1 port map( D => siso_data_in(8), CEB => n162, CK =>
                           clk, RB => resetn, Q => in_buf_248_port);
   in_buf_reg_0_22 : DFERPQ1 port map( D => siso_data_in(6), CEB => n162, CK =>
                           clk, RB => resetn, Q => in_buf_246_port);
   in_buf_reg_0_20 : DFERPQ1 port map( D => siso_data_in(4), CEB => n162, CK =>
                           clk, RB => resetn, Q => in_buf_244_port);
   in_buf_reg_0_18 : DFERPQ1 port map( D => siso_data_in(2), CEB => n162, CK =>
                           clk, RB => resetn, Q => in_buf_242_port);
   in_buf_reg_0_16 : DFERPQ1 port map( D => siso_data_in(0), CEB => n162, CK =>
                           clk, RB => resetn, Q => in_buf_240_port);
   in_buf_reg_0_14 : DFERPQ1 port map( D => siso_data_in(14), CEB => n163, CK 
                           => clk, RB => resetn, Q => in_buf_238_port);
   in_buf_reg_0_12 : DFERPQ1 port map( D => siso_data_in(12), CEB => n163, CK 
                           => clk, RB => resetn, Q => in_buf_236_port);
   in_buf_reg_0_10 : DFERPQ1 port map( D => siso_data_in(10), CEB => n163, CK 
                           => clk, RB => resetn, Q => in_buf_234_port);
   in_buf_reg_0_8 : DFERPQ1 port map( D => siso_data_in(8), CEB => n163, CK => 
                           clk, RB => resetn, Q => in_buf_232_port);
   in_buf_reg_0_6 : DFERPQ1 port map( D => siso_data_in(6), CEB => n163, CK => 
                           clk, RB => resetn, Q => in_buf_230_port);
   in_buf_reg_0_4 : DFERPQ1 port map( D => siso_data_in(4), CEB => n163, CK => 
                           clk, RB => resetn, Q => in_buf_228_port);
   in_buf_reg_0_2 : DFERPQ1 port map( D => siso_data_in(2), CEB => n163, CK => 
                           clk, RB => resetn, Q => in_buf_226_port);
   in_buf_reg_4_14 : DFERPQ1 port map( D => siso_data_in(14), CEB => n171, CK 
                           => clk, RB => resetn, Q => in_buf_110_port);
   in_buf_reg_4_12 : DFERPQ1 port map( D => siso_data_in(12), CEB => n171, CK 
                           => clk, RB => resetn, Q => in_buf_108_port);
   in_buf_reg_4_10 : DFERPQ1 port map( D => siso_data_in(10), CEB => n171, CK 
                           => clk, RB => resetn, Q => in_buf_106_port);
   in_buf_reg_4_8 : DFERPQ1 port map( D => siso_data_in(8), CEB => n171, CK => 
                           clk, RB => resetn, Q => in_buf_104_port);
   in_buf_reg_4_6 : DFERPQ1 port map( D => siso_data_in(6), CEB => n171, CK => 
                           clk, RB => resetn, Q => in_buf_102_port);
   in_buf_reg_4_4 : DFERPQ1 port map( D => siso_data_in(4), CEB => n171, CK => 
                           clk, RB => resetn, Q => in_buf_100_port);
   in_buf_reg_4_2 : DFERPQ1 port map( D => siso_data_in(2), CEB => n171, CK => 
                           clk, RB => resetn, Q => in_buf_98_port);
   in_buf_reg_3_0 : DFERPQ1 port map( D => siso_data_in(0), CEB => n169, CK => 
                           clk, RB => resetn, Q => in_buf_128_port);
   in_buf_reg_2_0 : DFERPQ1 port map( D => siso_data_in(0), CEB => n167, CK => 
                           clk, RB => resetn, Q => in_buf_160_port);
   in_buf_reg_6_0 : DFERPQ1 port map( D => siso_data_in(0), CEB => n175, CK => 
                           clk, RB => resetn, Q => in_buf_32_port);
   in_buf_reg_5_0 : DFERPQ1 port map( D => siso_data_in(0), CEB => n173, CK => 
                           clk, RB => resetn, Q => in_buf_64_port);
   out_buf_reg_7_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_15_port);
   out_buf_reg_7_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_14_port);
   out_buf_reg_7_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_13_port);
   out_buf_reg_7_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_12_port);
   out_buf_reg_7_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_11_port);
   out_buf_reg_7_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_10_port);
   out_buf_reg_7_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n246, CK 
                           => clk, RB => resetn, Q => out_buf_9_port);
   out_buf_reg_7_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n246, CK 
                           => clk, RB => resetn, Q => out_buf_8_port);
   out_buf_reg_7_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n246, CK 
                           => clk, RB => resetn, Q => out_buf_7_port);
   out_buf_reg_7_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n246, CK 
                           => clk, RB => resetn, Q => out_buf_6_port);
   out_buf_reg_7_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n246, CK 
                           => clk, RB => resetn, Q => out_buf_5_port);
   out_buf_reg_7_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n246, CK 
                           => clk, RB => resetn, Q => out_buf_4_port);
   out_buf_reg_7_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n246, CK 
                           => clk, RB => resetn, Q => out_buf_3_port);
   out_buf_reg_7_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n246, CK 
                           => clk, RB => resetn, Q => out_buf_2_port);
   out_buf_reg_7_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n246, CK 
                           => clk, RB => resetn, Q => out_buf_1_port);
   out_buf_reg_7_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n246, CK 
                           => clk, RB => resetn, Q => out_buf_0_port);
   in_buf_reg_1_0 : DFERPQ1 port map( D => siso_data_in(0), CEB => n165, CK => 
                           clk, RB => resetn, Q => in_buf_192_port);
   out_buf_reg_3_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => n253, CK
                           => clk, RB => resetn, Q => out_buf_143_port);
   out_buf_reg_3_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => n253, CK
                           => clk, RB => resetn, Q => out_buf_142_port);
   out_buf_reg_3_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => n253, CK
                           => clk, RB => resetn, Q => out_buf_141_port);
   out_buf_reg_3_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => n253, CK
                           => clk, RB => resetn, Q => out_buf_140_port);
   out_buf_reg_3_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => n253, CK
                           => clk, RB => resetn, Q => out_buf_139_port);
   out_buf_reg_3_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => n253, CK
                           => clk, RB => resetn, Q => out_buf_138_port);
   out_buf_reg_3_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n253, CK 
                           => clk, RB => resetn, Q => out_buf_137_port);
   out_buf_reg_3_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n253, CK 
                           => clk, RB => resetn, Q => out_buf_136_port);
   out_buf_reg_3_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n253, CK 
                           => clk, RB => resetn, Q => out_buf_135_port);
   out_buf_reg_3_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n253, CK 
                           => clk, RB => resetn, Q => out_buf_134_port);
   out_buf_reg_3_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n253, CK 
                           => clk, RB => resetn, Q => out_buf_133_port);
   out_buf_reg_3_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n253, CK 
                           => clk, RB => resetn, Q => out_buf_132_port);
   out_buf_reg_3_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n253, CK 
                           => clk, RB => resetn, Q => out_buf_131_port);
   out_buf_reg_3_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n253, CK 
                           => clk, RB => resetn, Q => out_buf_130_port);
   out_buf_reg_3_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n253, CK 
                           => clk, RB => resetn, Q => out_buf_129_port);
   out_buf_reg_3_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n253, CK 
                           => clk, RB => resetn, Q => out_buf_128_port);
   in_buf_reg_0_0 : DFERPQ1 port map( D => siso_data_in(0), CEB => n163, CK => 
                           clk, RB => resetn, Q => in_buf_224_port);
   in_buf_reg_4_0 : DFERPQ1 port map( D => siso_data_in(0), CEB => n171, CK => 
                           clk, RB => resetn, Q => in_buf_96_port);
   out_buf_reg_2_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_175_port);
   out_buf_reg_2_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_174_port);
   out_buf_reg_2_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_173_port);
   out_buf_reg_2_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_172_port);
   out_buf_reg_2_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_171_port);
   out_buf_reg_2_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_170_port);
   out_buf_reg_2_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n252, CK 
                           => clk, RB => resetn, Q => out_buf_169_port);
   out_buf_reg_2_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n252, CK 
                           => clk, RB => resetn, Q => out_buf_168_port);
   out_buf_reg_2_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n252, CK 
                           => clk, RB => resetn, Q => out_buf_167_port);
   out_buf_reg_2_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n252, CK 
                           => clk, RB => resetn, Q => out_buf_166_port);
   out_buf_reg_2_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n252, CK 
                           => clk, RB => resetn, Q => out_buf_165_port);
   out_buf_reg_2_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n252, CK 
                           => clk, RB => resetn, Q => out_buf_164_port);
   out_buf_reg_2_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n252, CK 
                           => clk, RB => resetn, Q => out_buf_163_port);
   out_buf_reg_2_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n252, CK 
                           => clk, RB => resetn, Q => out_buf_162_port);
   out_buf_reg_2_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n252, CK 
                           => clk, RB => resetn, Q => out_buf_161_port);
   out_buf_reg_2_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n252, CK 
                           => clk, RB => resetn, Q => out_buf_160_port);
   out_buf_reg_6_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_47_port);
   out_buf_reg_6_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_46_port);
   out_buf_reg_6_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_45_port);
   out_buf_reg_6_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_44_port);
   out_buf_reg_6_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_43_port);
   out_buf_reg_6_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_42_port);
   out_buf_reg_6_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n251, CK 
                           => clk, RB => resetn, Q => out_buf_41_port);
   out_buf_reg_6_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n251, CK 
                           => clk, RB => resetn, Q => out_buf_40_port);
   out_buf_reg_6_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n251, CK 
                           => clk, RB => resetn, Q => out_buf_39_port);
   out_buf_reg_6_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n251, CK 
                           => clk, RB => resetn, Q => out_buf_38_port);
   out_buf_reg_6_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n251, CK 
                           => clk, RB => resetn, Q => out_buf_37_port);
   out_buf_reg_6_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n251, CK 
                           => clk, RB => resetn, Q => out_buf_36_port);
   out_buf_reg_6_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n251, CK 
                           => clk, RB => resetn, Q => out_buf_35_port);
   out_buf_reg_6_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n251, CK 
                           => clk, RB => resetn, Q => out_buf_34_port);
   out_buf_reg_6_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n251, CK 
                           => clk, RB => resetn, Q => out_buf_33_port);
   out_buf_reg_6_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n251, CK 
                           => clk, RB => resetn, Q => out_buf_32_port);
   out_buf_reg_7_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_31_port);
   out_buf_reg_7_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_30_port);
   out_buf_reg_7_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_29_port);
   out_buf_reg_7_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_28_port);
   out_buf_reg_7_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_27_port);
   out_buf_reg_7_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_26_port);
   out_buf_reg_7_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_25_port);
   out_buf_reg_7_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_24_port);
   out_buf_reg_7_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_23_port);
   out_buf_reg_7_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_22_port);
   out_buf_reg_7_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_21_port);
   out_buf_reg_7_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_20_port);
   out_buf_reg_7_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_19_port);
   out_buf_reg_7_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_18_port);
   out_buf_reg_7_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_17_port);
   out_buf_reg_7_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_16_port);
   out_buf_reg_5_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_79_port);
   out_buf_reg_5_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_78_port);
   out_buf_reg_5_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_77_port);
   out_buf_reg_5_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_76_port);
   out_buf_reg_5_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_75_port);
   out_buf_reg_5_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_74_port);
   out_buf_reg_5_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n250, CK 
                           => clk, RB => resetn, Q => out_buf_73_port);
   out_buf_reg_5_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n250, CK 
                           => clk, RB => resetn, Q => out_buf_72_port);
   out_buf_reg_5_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n250, CK 
                           => clk, RB => resetn, Q => out_buf_71_port);
   out_buf_reg_5_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n250, CK 
                           => clk, RB => resetn, Q => out_buf_70_port);
   out_buf_reg_5_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n250, CK 
                           => clk, RB => resetn, Q => out_buf_69_port);
   out_buf_reg_5_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n250, CK 
                           => clk, RB => resetn, Q => out_buf_68_port);
   out_buf_reg_5_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n250, CK 
                           => clk, RB => resetn, Q => out_buf_67_port);
   out_buf_reg_5_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n250, CK 
                           => clk, RB => resetn, Q => out_buf_66_port);
   out_buf_reg_5_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n250, CK 
                           => clk, RB => resetn, Q => out_buf_65_port);
   out_buf_reg_5_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n250, CK 
                           => clk, RB => resetn, Q => out_buf_64_port);
   out_buf_reg_3_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => n253, CK
                           => clk, RB => resetn, Q => out_buf_159_port);
   out_buf_reg_3_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => n253, CK
                           => clk, RB => resetn, Q => out_buf_158_port);
   out_buf_reg_3_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => n253, CK
                           => clk, RB => resetn, Q => out_buf_157_port);
   out_buf_reg_3_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => n253, CK
                           => clk, RB => resetn, Q => out_buf_156_port);
   out_buf_reg_3_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => n253, CK
                           => clk, RB => resetn, Q => out_buf_155_port);
   out_buf_reg_3_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => n253, CK
                           => clk, RB => resetn, Q => out_buf_154_port);
   out_buf_reg_3_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => n253, CK
                           => clk, RB => resetn, Q => out_buf_153_port);
   out_buf_reg_3_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => n253, CK
                           => clk, RB => resetn, Q => out_buf_152_port);
   out_buf_reg_3_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => n253, CK
                           => clk, RB => resetn, Q => out_buf_151_port);
   out_buf_reg_3_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => n253, CK
                           => clk, RB => resetn, Q => out_buf_150_port);
   out_buf_reg_3_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => n253, CK
                           => clk, RB => resetn, Q => out_buf_149_port);
   out_buf_reg_3_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => n253, CK
                           => clk, RB => resetn, Q => out_buf_148_port);
   out_buf_reg_3_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => n253, CK
                           => clk, RB => resetn, Q => out_buf_147_port);
   out_buf_reg_3_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => n253, CK
                           => clk, RB => resetn, Q => out_buf_146_port);
   out_buf_reg_3_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => n253, CK
                           => clk, RB => resetn, Q => out_buf_145_port);
   out_buf_reg_3_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => n253, CK
                           => clk, RB => resetn, Q => out_buf_144_port);
   out_buf_reg_1_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_207_port);
   out_buf_reg_1_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_206_port);
   out_buf_reg_1_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_205_port);
   out_buf_reg_1_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_204_port);
   out_buf_reg_1_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_203_port);
   out_buf_reg_1_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_202_port);
   out_buf_reg_1_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n249, CK 
                           => clk, RB => resetn, Q => out_buf_201_port);
   out_buf_reg_1_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n249, CK 
                           => clk, RB => resetn, Q => out_buf_200_port);
   out_buf_reg_1_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n249, CK 
                           => clk, RB => resetn, Q => out_buf_199_port);
   out_buf_reg_1_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n249, CK 
                           => clk, RB => resetn, Q => out_buf_198_port);
   out_buf_reg_1_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n249, CK 
                           => clk, RB => resetn, Q => out_buf_197_port);
   out_buf_reg_1_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n249, CK 
                           => clk, RB => resetn, Q => out_buf_196_port);
   out_buf_reg_1_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n249, CK 
                           => clk, RB => resetn, Q => out_buf_195_port);
   out_buf_reg_1_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n249, CK 
                           => clk, RB => resetn, Q => out_buf_194_port);
   out_buf_reg_1_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n249, CK 
                           => clk, RB => resetn, Q => out_buf_193_port);
   out_buf_reg_1_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n249, CK 
                           => clk, RB => resetn, Q => out_buf_192_port);
   out_buf_reg_2_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_191_port);
   out_buf_reg_2_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_190_port);
   out_buf_reg_2_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_189_port);
   out_buf_reg_2_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_188_port);
   out_buf_reg_2_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_187_port);
   out_buf_reg_2_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_186_port);
   out_buf_reg_2_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_185_port);
   out_buf_reg_2_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_184_port);
   out_buf_reg_2_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_183_port);
   out_buf_reg_2_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_182_port);
   out_buf_reg_2_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_181_port);
   out_buf_reg_2_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_180_port);
   out_buf_reg_2_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_179_port);
   out_buf_reg_2_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_178_port);
   out_buf_reg_2_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_177_port);
   out_buf_reg_2_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_176_port);
   out_buf_reg_6_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_63_port);
   out_buf_reg_6_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_62_port);
   out_buf_reg_6_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_61_port);
   out_buf_reg_6_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_60_port);
   out_buf_reg_6_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_59_port);
   out_buf_reg_6_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_58_port);
   out_buf_reg_6_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_57_port);
   out_buf_reg_6_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_56_port);
   out_buf_reg_6_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_55_port);
   out_buf_reg_6_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_54_port);
   out_buf_reg_6_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_53_port);
   out_buf_reg_6_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_52_port);
   out_buf_reg_6_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_51_port);
   out_buf_reg_6_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_50_port);
   out_buf_reg_6_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_49_port);
   out_buf_reg_6_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_48_port);
   out_buf_reg_0_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_239_port);
   out_buf_reg_0_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_238_port);
   out_buf_reg_0_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_237_port);
   out_buf_reg_0_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_236_port);
   out_buf_reg_0_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_235_port);
   out_buf_reg_0_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_234_port);
   out_buf_reg_0_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n248, CK 
                           => clk, RB => resetn, Q => out_buf_233_port);
   out_buf_reg_0_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n248, CK 
                           => clk, RB => resetn, Q => out_buf_232_port);
   out_buf_reg_0_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n248, CK 
                           => clk, RB => resetn, Q => out_buf_231_port);
   out_buf_reg_0_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n248, CK 
                           => clk, RB => resetn, Q => out_buf_230_port);
   out_buf_reg_0_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n248, CK 
                           => clk, RB => resetn, Q => out_buf_229_port);
   out_buf_reg_0_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n248, CK 
                           => clk, RB => resetn, Q => out_buf_228_port);
   out_buf_reg_0_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n248, CK 
                           => clk, RB => resetn, Q => out_buf_227_port);
   out_buf_reg_0_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n248, CK 
                           => clk, RB => resetn, Q => out_buf_226_port);
   out_buf_reg_0_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n248, CK 
                           => clk, RB => resetn, Q => out_buf_225_port);
   out_buf_reg_0_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n248, CK 
                           => clk, RB => resetn, Q => out_buf_224_port);
   out_buf_reg_4_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_111_port);
   out_buf_reg_4_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_110_port);
   out_buf_reg_4_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_109_port);
   out_buf_reg_4_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_108_port);
   out_buf_reg_4_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_107_port);
   out_buf_reg_4_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_106_port);
   out_buf_reg_4_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n247, CK 
                           => clk, RB => resetn, Q => out_buf_105_port);
   out_buf_reg_4_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n247, CK 
                           => clk, RB => resetn, Q => out_buf_104_port);
   out_buf_reg_4_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n247, CK 
                           => clk, RB => resetn, Q => out_buf_103_port);
   out_buf_reg_4_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n247, CK 
                           => clk, RB => resetn, Q => out_buf_102_port);
   out_buf_reg_4_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n247, CK 
                           => clk, RB => resetn, Q => out_buf_101_port);
   out_buf_reg_4_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n247, CK 
                           => clk, RB => resetn, Q => out_buf_100_port);
   out_buf_reg_4_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n247, CK 
                           => clk, RB => resetn, Q => out_buf_99_port);
   out_buf_reg_4_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n247, CK 
                           => clk, RB => resetn, Q => out_buf_98_port);
   out_buf_reg_4_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n247, CK 
                           => clk, RB => resetn, Q => out_buf_97_port);
   out_buf_reg_4_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n247, CK 
                           => clk, RB => resetn, Q => out_buf_96_port);
   out_buf_reg_5_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_95_port);
   out_buf_reg_5_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_94_port);
   out_buf_reg_5_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_93_port);
   out_buf_reg_5_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_92_port);
   out_buf_reg_5_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_91_port);
   out_buf_reg_5_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_90_port);
   out_buf_reg_5_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_89_port);
   out_buf_reg_5_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_88_port);
   out_buf_reg_5_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_87_port);
   out_buf_reg_5_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_86_port);
   out_buf_reg_5_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_85_port);
   out_buf_reg_5_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_84_port);
   out_buf_reg_5_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_83_port);
   out_buf_reg_5_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_82_port);
   out_buf_reg_5_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_81_port);
   out_buf_reg_5_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_80_port);
   out_buf_reg_1_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_223_port);
   out_buf_reg_1_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_222_port);
   out_buf_reg_1_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_221_port);
   out_buf_reg_1_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_220_port);
   out_buf_reg_1_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_219_port);
   out_buf_reg_1_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_218_port);
   out_buf_reg_1_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_217_port);
   out_buf_reg_1_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_216_port);
   out_buf_reg_1_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_215_port);
   out_buf_reg_1_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_214_port);
   out_buf_reg_1_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_213_port);
   out_buf_reg_1_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_212_port);
   out_buf_reg_1_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_211_port);
   out_buf_reg_1_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_210_port);
   out_buf_reg_1_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_209_port);
   out_buf_reg_1_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_208_port);
   out_buf_reg_0_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_255_port);
   out_buf_reg_0_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_254_port);
   out_buf_reg_0_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_253_port);
   out_buf_reg_0_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_252_port);
   out_buf_reg_0_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_251_port);
   out_buf_reg_0_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_250_port);
   out_buf_reg_0_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_249_port);
   out_buf_reg_0_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_248_port);
   out_buf_reg_0_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_247_port);
   out_buf_reg_0_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_246_port);
   out_buf_reg_0_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_245_port);
   out_buf_reg_0_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_244_port);
   out_buf_reg_0_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_243_port);
   out_buf_reg_0_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_242_port);
   out_buf_reg_0_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_241_port);
   out_buf_reg_0_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_240_port);
   out_buf_reg_4_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_127_port);
   out_buf_reg_4_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_126_port);
   out_buf_reg_4_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_125_port);
   out_buf_reg_4_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_124_port);
   out_buf_reg_4_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_123_port);
   out_buf_reg_4_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_122_port);
   out_buf_reg_4_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_121_port);
   out_buf_reg_4_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_120_port);
   out_buf_reg_4_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_119_port);
   out_buf_reg_4_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_118_port);
   out_buf_reg_4_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_117_port);
   out_buf_reg_4_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_116_port);
   out_buf_reg_4_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_115_port);
   out_buf_reg_4_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_114_port);
   out_buf_reg_4_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_113_port);
   out_buf_reg_4_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_112_port);
   out_trigger_reg : DFFRPQ1 port map( D => n240, CK => clk, RB => resetn, Q =>
                           out_trigger);
   read_comp_res_reg : DFERPQ1 port map( D => avs_writedata(2), CEB => n179, CK
                           => clk, RB => resetn, Q => read_comp_res);
   in_counter_reg_0 : DFERPQ1 port map( D => n155, CEB => n800, CK => clk, RB 
                           => resetn, Q => in_counter_0_port);
   in_counter_reg_2 : DFFRPQ1 port map( D => n238, CK => clk, RB => resetn, Q 
                           => in_counter_2_port);
   in_counter_reg_1 : DFFRPQ1 port map( D => n237, CK => clk, RB => resetn, Q 
                           => in_counter_1_port);
   in_busy_reg : DFFRPQ1 port map( D => n239, CK => clk, RB => resetn, Q => 
                           in_busy);
   odd_reg : DFFRPQ1 port map( D => n156, CK => clk, RB => resetn, Q => odd);
   out_busy_reg : DFFRPQ1 port map( D => n234, CK => clk, RB => resetn, Q => 
                           out_busy);
   odd_reg2 : DFFRPQ1 port map( D => n154, CK => clk, RB => resetn, Q => odd1);
   operand_load_reg : DFERPQ1 port map( D => avs_writedata(1), CEB => n179, CK 
                           => clk, RB => resetn, Q => operand_load);
   coeff_load_reg : DFERPQ1 port map( D => avs_writedata(0), CEB => n179, CK =>
                           clk, RB => resetn, Q => coeff_load);
   out_counter_reg_0 : DFFRPQ1 port map( D => n236, CK => clk, RB => resetn, Q 
                           => N62);
   out_counter_reg_2 : DFFRPQ1 port map( D => n235, CK => clk, RB => resetn, Q 
                           => N64);
   out_counter_reg_1 : DFFRPQ1 port map( D => n201, CK => clk, RB => resetn, Q 
                           => N63);
   operand_regs_reg_3_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_159_port);
   operand_regs_reg_5_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_95_port);
   operand_regs_reg_1_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_223_port);
   coeff_memory_reg_0_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_31);
   coeff_memory_reg_1_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_31);
   coeff_memory_reg_2_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_31);
   coeff_memory_reg_3_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_31);
   coeff_memory_reg_4_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_31);
   operand_regs_reg_2_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_191_port);
   operand_regs_reg_4_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_127_port);
   operand_regs_reg_6_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_63_port);
   operand_regs_reg_7_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_31_port);
   operand_regs_reg_0_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_255_port);
   operand_regs_reg_3_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_158_port);
   operand_regs_reg_5_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_94_port);
   operand_regs_reg_3_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_157_port);
   operand_regs_reg_5_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_93_port);
   coeff_memory_reg_0_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_30);
   coeff_memory_reg_1_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_30);
   coeff_memory_reg_2_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_30);
   coeff_memory_reg_3_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_30);
   coeff_memory_reg_4_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_30);
   operand_regs_reg_2_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_190_port);
   operand_regs_reg_4_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_126_port);
   operand_regs_reg_6_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_62_port);
   operand_regs_reg_1_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_222_port);
   operand_regs_reg_7_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_30_port);
   operand_regs_reg_0_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_254_port);
   operand_regs_reg_1_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_221_port);
   operand_regs_reg_3_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_156_port);
   operand_regs_reg_5_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_92_port);
   coeff_memory_reg_0_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_29);
   coeff_memory_reg_1_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_29);
   coeff_memory_reg_2_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_29);
   coeff_memory_reg_3_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_29);
   coeff_memory_reg_4_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_29);
   operand_regs_reg_2_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_189_port);
   operand_regs_reg_4_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_125_port);
   operand_regs_reg_6_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_61_port);
   operand_regs_reg_7_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_29_port);
   operand_regs_reg_0_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_253_port);
   operand_regs_reg_1_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_220_port);
   operand_regs_reg_3_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_155_port);
   operand_regs_reg_5_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_91_port);
   coeff_memory_reg_0_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_28);
   coeff_memory_reg_1_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_28);
   coeff_memory_reg_2_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_28);
   coeff_memory_reg_3_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_28);
   coeff_memory_reg_4_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_28);
   operand_regs_reg_2_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_188_port);
   operand_regs_reg_4_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_124_port);
   operand_regs_reg_6_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_60_port);
   operand_regs_reg_7_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_28_port);
   operand_regs_reg_0_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_252_port);
   avs_readdata_reg_30 : DFFSPQ1 port map( D => n203, CK => clk, SB => resetn, 
                           Q => avs_readdata_30_port);
   avs_readdata_reg_28 : DFFSPQ1 port map( D => n205, CK => clk, SB => resetn, 
                           Q => avs_readdata_28_port);
   avs_readdata_reg_26 : DFFSPQ1 port map( D => n207, CK => clk, SB => resetn, 
                           Q => avs_readdata_26_port);
   avs_readdata_reg_24 : DFFSPQ1 port map( D => n209, CK => clk, SB => resetn, 
                           Q => avs_readdata_24_port);
   avs_readdata_reg_22 : DFFSPQ1 port map( D => n211, CK => clk, SB => resetn, 
                           Q => avs_readdata_22_port);
   avs_readdata_reg_20 : DFFSPQ1 port map( D => n213, CK => clk, SB => resetn, 
                           Q => avs_readdata_20_port);
   avs_readdata_reg_18 : DFFSPQ1 port map( D => n215, CK => clk, SB => resetn, 
                           Q => avs_readdata_18_port);
   avs_readdata_reg_16 : DFFSPQ1 port map( D => n217, CK => clk, SB => resetn, 
                           Q => avs_readdata_16_port);
   avs_readdata_reg_14 : DFFSPQ1 port map( D => n219, CK => clk, SB => resetn, 
                           Q => avs_readdata_14_port);
   avs_readdata_reg_12 : DFFSPQ1 port map( D => n221, CK => clk, SB => resetn, 
                           Q => avs_readdata_12_port);
   avs_readdata_reg_10 : DFFSPQ1 port map( D => n223, CK => clk, SB => resetn, 
                           Q => avs_readdata_10_port);
   avs_readdata_reg_8 : DFFSPQ1 port map( D => n225, CK => clk, SB => resetn, Q
                           => avs_readdata_8_port);
   avs_readdata_reg_6 : DFFSPQ1 port map( D => n227, CK => clk, SB => resetn, Q
                           => avs_readdata_6_port);
   avs_readdata_reg_4 : DFFSPQ1 port map( D => n229, CK => clk, SB => resetn, Q
                           => avs_readdata_4_port);
   avs_readdata_reg_2 : DFFSPQ1 port map( D => n231, CK => clk, SB => resetn, Q
                           => avs_readdata_2_port);
   avs_readdata_reg_0 : DFFSPQ1 port map( D => n233, CK => clk, SB => resetn, Q
                           => avs_readdata_0_port);
   operand_regs_reg_3_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_154_port);
   operand_regs_reg_5_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_90_port);
   operand_regs_reg_1_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_219_port);
   avs_readdata_reg_31 : DFFRPQ1 port map( D => n202, CK => clk, RB => resetn, 
                           Q => avs_readdata_31_port);
   avs_readdata_reg_29 : DFFRPQ1 port map( D => n204, CK => clk, RB => resetn, 
                           Q => avs_readdata_29_port);
   avs_readdata_reg_27 : DFFRPQ1 port map( D => n206, CK => clk, RB => resetn, 
                           Q => avs_readdata_27_port);
   avs_readdata_reg_25 : DFFRPQ1 port map( D => n208, CK => clk, RB => resetn, 
                           Q => avs_readdata_25_port);
   avs_readdata_reg_23 : DFFRPQ1 port map( D => n210, CK => clk, RB => resetn, 
                           Q => avs_readdata_23_port);
   avs_readdata_reg_21 : DFFRPQ1 port map( D => n212, CK => clk, RB => resetn, 
                           Q => avs_readdata_21_port);
   avs_readdata_reg_19 : DFFRPQ1 port map( D => n214, CK => clk, RB => resetn, 
                           Q => avs_readdata_19_port);
   avs_readdata_reg_17 : DFFRPQ1 port map( D => n216, CK => clk, RB => resetn, 
                           Q => avs_readdata_17_port);
   avs_readdata_reg_15 : DFFRPQ1 port map( D => n218, CK => clk, RB => resetn, 
                           Q => avs_readdata_15_port);
   avs_readdata_reg_13 : DFFRPQ1 port map( D => n220, CK => clk, RB => resetn, 
                           Q => avs_readdata_13_port);
   avs_readdata_reg_11 : DFFRPQ1 port map( D => n222, CK => clk, RB => resetn, 
                           Q => avs_readdata_11_port);
   avs_readdata_reg_9 : DFFRPQ1 port map( D => n224, CK => clk, RB => resetn, Q
                           => avs_readdata_9_port);
   avs_readdata_reg_7 : DFFRPQ1 port map( D => n226, CK => clk, RB => resetn, Q
                           => avs_readdata_7_port);
   avs_readdata_reg_5 : DFFRPQ1 port map( D => n228, CK => clk, RB => resetn, Q
                           => avs_readdata_5_port);
   avs_readdata_reg_3 : DFFRPQ1 port map( D => n230, CK => clk, RB => resetn, Q
                           => avs_readdata_3_port);
   avs_readdata_reg_1 : DFFRPQ1 port map( D => n232, CK => clk, RB => resetn, Q
                           => avs_readdata_1_port);
   stop_sim_reg : DFFRPQ1 port map( D => n157, CK => clk, RB => resetn, Q => 
                           stop_sim_port);
   operand_regs_reg_1_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_218_port);
   coeff_memory_reg_0_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_27);
   coeff_memory_reg_1_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_27);
   coeff_memory_reg_2_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_27);
   coeff_memory_reg_3_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_27);
   coeff_memory_reg_4_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_27);
   operand_regs_reg_2_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_187_port);
   operand_regs_reg_4_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_123_port);
   operand_regs_reg_6_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_59_port);
   operand_regs_reg_7_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_27_port);
   operand_regs_reg_0_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_251_port);
   operand_regs_reg_3_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_153_port);
   operand_regs_reg_5_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_89_port);
   coeff_memory_reg_0_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_26);
   coeff_memory_reg_1_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_26);
   coeff_memory_reg_2_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_26);
   coeff_memory_reg_3_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_26);
   coeff_memory_reg_4_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_26);
   operand_regs_reg_2_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_186_port);
   operand_regs_reg_4_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_122_port);
   operand_regs_reg_6_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_58_port);
   operand_regs_reg_7_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_26_port);
   operand_regs_reg_0_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_250_port);
   operand_regs_reg_1_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_217_port);
   operand_regs_reg_3_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_152_port);
   operand_regs_reg_5_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_88_port);
   operand_regs_reg_1_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_216_port);
   coeff_memory_reg_0_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_25);
   coeff_memory_reg_1_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_25);
   coeff_memory_reg_2_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_25);
   coeff_memory_reg_3_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_25);
   coeff_memory_reg_4_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_25);
   operand_regs_reg_2_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_185_port);
   operand_regs_reg_4_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_121_port);
   operand_regs_reg_6_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_57_port);
   operand_regs_reg_3_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_151_port);
   operand_regs_reg_5_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_87_port);
   operand_regs_reg_7_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_25_port);
   operand_regs_reg_0_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_249_port);
   operand_regs_reg_1_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_215_port);
   coeff_memory_reg_0_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_24);
   coeff_memory_reg_1_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_24);
   coeff_memory_reg_2_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_24);
   coeff_memory_reg_3_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_24);
   coeff_memory_reg_4_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_24);
   operand_regs_reg_2_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_184_port);
   operand_regs_reg_4_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_120_port);
   operand_regs_reg_6_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_56_port);
   operand_regs_reg_7_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_24_port);
   operand_regs_reg_0_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_248_port);
   coeff_memory_reg_0_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_23);
   coeff_memory_reg_1_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_23);
   coeff_memory_reg_2_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_23);
   coeff_memory_reg_3_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_23);
   coeff_memory_reg_4_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_23);
   operand_regs_reg_2_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_183_port);
   operand_regs_reg_4_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_119_port);
   operand_regs_reg_6_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_55_port);
   operand_regs_reg_7_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_23_port);
   operand_regs_reg_0_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_247_port);
   operand_regs_reg_3_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_150_port);
   operand_regs_reg_5_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_86_port);
   operand_regs_reg_3_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_149_port);
   operand_regs_reg_5_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_85_port);
   coeff_memory_reg_0_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_22);
   coeff_memory_reg_1_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_22);
   coeff_memory_reg_2_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_22);
   coeff_memory_reg_3_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_22);
   coeff_memory_reg_4_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_22);
   operand_regs_reg_2_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_182_port);
   operand_regs_reg_4_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_118_port);
   operand_regs_reg_6_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_54_port);
   operand_regs_reg_7_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_22_port);
   operand_regs_reg_0_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_246_port);
   operand_regs_reg_1_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_214_port);
   operand_regs_reg_3_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_148_port);
   operand_regs_reg_5_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_84_port);
   coeff_memory_reg_0_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_21);
   coeff_memory_reg_1_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_21);
   coeff_memory_reg_2_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_21);
   coeff_memory_reg_3_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_21);
   coeff_memory_reg_4_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_21);
   operand_regs_reg_2_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_181_port);
   operand_regs_reg_4_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_117_port);
   operand_regs_reg_6_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_53_port);
   operand_regs_reg_1_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_213_port);
   operand_regs_reg_3_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_147_port);
   operand_regs_reg_5_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_83_port);
   operand_regs_reg_7_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_21_port);
   operand_regs_reg_0_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_245_port);
   operand_regs_reg_3_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_144_port);
   operand_regs_reg_5_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_80_port);
   operand_regs_reg_3_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_146_port);
   operand_regs_reg_5_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_82_port);
   operand_regs_reg_3_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_143_port);
   operand_regs_reg_5_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_79_port);
   operand_regs_reg_3_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_139_port);
   operand_regs_reg_5_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_75_port);
   operand_regs_reg_3_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_145_port);
   operand_regs_reg_5_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_81_port);
   operand_regs_reg_3_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_142_port);
   operand_regs_reg_5_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_78_port);
   operand_regs_reg_3_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_141_port);
   operand_regs_reg_5_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_77_port);
   operand_regs_reg_3_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_140_port);
   operand_regs_reg_5_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_76_port);
   operand_regs_reg_1_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_212_port);
   coeff_memory_reg_0_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_20);
   coeff_memory_reg_1_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_20);
   coeff_memory_reg_2_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_20);
   coeff_memory_reg_3_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_20);
   coeff_memory_reg_4_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_20);
   operand_regs_reg_2_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_180_port);
   operand_regs_reg_4_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_116_port);
   operand_regs_reg_6_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_52_port);
   operand_regs_reg_1_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_211_port);
   operand_regs_reg_7_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_20_port);
   operand_regs_reg_0_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_244_port);
   operand_regs_reg_1_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_208_port);
   operand_regs_reg_3_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_138_port);
   operand_regs_reg_5_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_74_port);
   coeff_memory_reg_3_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n263,
                           CK => clk, RB => resetn, Q => coeff_memory_3_0);
   coeff_memory_reg_4_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n265,
                           CK => clk, RB => resetn, Q => coeff_memory_4_0);
   operand_regs_reg_1_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_210_port);
   coeff_memory_reg_0_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n267,
                           CK => clk, RB => resetn, Q => coeff_memory_0_0);
   operand_regs_reg_6_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n256,
                           CK => clk, RB => resetn, Q => operand_regs_32_port);
   coeff_memory_reg_0_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_19);
   coeff_memory_reg_1_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_19);
   coeff_memory_reg_2_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_19);
   coeff_memory_reg_3_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_19);
   coeff_memory_reg_4_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_19);
   coeff_memory_reg_1_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n266,
                           CK => clk, RB => resetn, Q => coeff_memory_1_0);
   coeff_memory_reg_2_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n264,
                           CK => clk, RB => resetn, Q => coeff_memory_2_0);
   operand_regs_reg_2_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_179_port);
   operand_regs_reg_4_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_115_port);
   operand_regs_reg_6_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_51_port);
   operand_regs_reg_2_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n258,
                           CK => clk, RB => resetn, Q => operand_regs_160_port)
                           ;
   operand_regs_reg_4_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n257,
                           CK => clk, RB => resetn, Q => operand_regs_96_port);
   operand_regs_reg_1_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_207_port);
   operand_regs_reg_7_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_19_port);
   operand_regs_reg_1_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_209_port);
   operand_regs_reg_0_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_243_port);
   coeff_memory_reg_0_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_18);
   coeff_memory_reg_1_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_18);
   coeff_memory_reg_2_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_18);
   coeff_memory_reg_3_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_18);
   coeff_memory_reg_4_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_18);
   operand_regs_reg_2_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_178_port);
   operand_regs_reg_4_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_114_port);
   operand_regs_reg_6_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_50_port);
   operand_regs_reg_3_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n261,
                           CK => clk, RB => resetn, Q => operand_regs_137_port)
                           ;
   operand_regs_reg_5_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n260,
                           CK => clk, RB => resetn, Q => operand_regs_73_port);
   operand_regs_reg_7_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_18_port);
   operand_regs_reg_0_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_242_port);
   operand_regs_reg_3_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n261,
                           CK => clk, RB => resetn, Q => operand_regs_132_port)
                           ;
   operand_regs_reg_5_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n260,
                           CK => clk, RB => resetn, Q => operand_regs_68_port);
   operand_regs_reg_3_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n261,
                           CK => clk, RB => resetn, Q => operand_regs_131_port)
                           ;
   operand_regs_reg_5_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n260,
                           CK => clk, RB => resetn, Q => operand_regs_67_port);
   operand_regs_reg_3_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n261,
                           CK => clk, RB => resetn, Q => operand_regs_128_port)
                           ;
   operand_regs_reg_5_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n260,
                           CK => clk, RB => resetn, Q => operand_regs_64_port);
   coeff_memory_reg_0_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_10);
   coeff_memory_reg_1_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_10);
   coeff_memory_reg_2_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_10);
   coeff_memory_reg_3_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_10);
   coeff_memory_reg_4_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_10);
   operand_regs_reg_2_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_170_port);
   operand_regs_reg_4_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_106_port);
   operand_regs_reg_6_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_42_port);
   operand_regs_reg_0_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_234_port);
   coeff_memory_reg_0_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_17);
   coeff_memory_reg_1_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_17);
   coeff_memory_reg_2_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_17);
   coeff_memory_reg_3_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_17);
   coeff_memory_reg_4_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_17);
   operand_regs_reg_2_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_177_port);
   operand_regs_reg_4_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_113_port);
   operand_regs_reg_6_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_49_port);
   operand_regs_reg_3_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n261,
                           CK => clk, RB => resetn, Q => operand_regs_133_port)
                           ;
   operand_regs_reg_5_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n260,
                           CK => clk, RB => resetn, Q => operand_regs_69_port);
   operand_regs_reg_7_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_17_port);
   operand_regs_reg_3_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n261,
                           CK => clk, RB => resetn, Q => operand_regs_129_port)
                           ;
   operand_regs_reg_5_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n260,
                           CK => clk, RB => resetn, Q => operand_regs_65_port);
   operand_regs_reg_0_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_241_port);
   coeff_memory_reg_0_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_16);
   coeff_memory_reg_1_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_16);
   coeff_memory_reg_2_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_16);
   coeff_memory_reg_3_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_16);
   coeff_memory_reg_4_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_16);
   operand_regs_reg_2_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_176_port);
   operand_regs_reg_4_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_112_port);
   operand_regs_reg_6_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_48_port);
   operand_regs_reg_3_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n261,
                           CK => clk, RB => resetn, Q => operand_regs_130_port)
                           ;
   operand_regs_reg_5_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n260,
                           CK => clk, RB => resetn, Q => operand_regs_66_port);
   coeff_memory_reg_0_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_14);
   coeff_memory_reg_1_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_14);
   coeff_memory_reg_2_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_14);
   coeff_memory_reg_3_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_14);
   coeff_memory_reg_4_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_14);
   operand_regs_reg_7_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_16_port);
   operand_regs_reg_3_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n261,
                           CK => clk, RB => resetn, Q => operand_regs_136_port)
                           ;
   operand_regs_reg_5_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n260,
                           CK => clk, RB => resetn, Q => operand_regs_72_port);
   operand_regs_reg_0_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n255,
                           CK => clk, RB => resetn, Q => operand_regs_224_port)
                           ;
   operand_regs_reg_0_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_240_port);
   operand_regs_reg_2_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_174_port);
   operand_regs_reg_4_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_110_port);
   operand_regs_reg_6_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_46_port);
   operand_regs_reg_3_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n261,
                           CK => clk, RB => resetn, Q => operand_regs_135_port)
                           ;
   operand_regs_reg_5_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n260,
                           CK => clk, RB => resetn, Q => operand_regs_71_port);
   operand_regs_reg_3_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n261,
                           CK => clk, RB => resetn, Q => operand_regs_134_port)
                           ;
   operand_regs_reg_5_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n260,
                           CK => clk, RB => resetn, Q => operand_regs_70_port);
   operand_regs_reg_0_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_238_port);
   operand_regs_reg_1_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_203_port);
   coeff_memory_reg_0_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_13);
   coeff_memory_reg_1_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_13);
   coeff_memory_reg_2_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_13);
   coeff_memory_reg_3_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_13);
   coeff_memory_reg_4_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_13);
   operand_regs_reg_7_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_14_port);
   operand_regs_reg_2_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_173_port);
   operand_regs_reg_4_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_109_port);
   operand_regs_reg_6_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_45_port);
   coeff_memory_reg_0_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_15);
   coeff_memory_reg_1_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_15);
   coeff_memory_reg_2_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_15);
   coeff_memory_reg_3_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_15);
   coeff_memory_reg_4_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_15);
   operand_regs_reg_2_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_175_port);
   operand_regs_reg_4_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_111_port);
   operand_regs_reg_6_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_47_port);
   coeff_memory_reg_0_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_12);
   coeff_memory_reg_1_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_12);
   coeff_memory_reg_2_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_12);
   coeff_memory_reg_3_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_12);
   coeff_memory_reg_4_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_12);
   operand_regs_reg_1_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_204_port);
   operand_regs_reg_7_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_13_port);
   operand_regs_reg_1_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_206_port);
   operand_regs_reg_0_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_237_port);
   operand_regs_reg_2_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_172_port);
   operand_regs_reg_4_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_108_port);
   operand_regs_reg_6_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_44_port);
   operand_regs_reg_1_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_205_port);
   operand_regs_reg_7_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_15_port);
   coeff_memory_reg_0_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n267,
                           CK => clk, RB => resetn, Q => coeff_memory_0_9);
   coeff_memory_reg_1_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n266,
                           CK => clk, RB => resetn, Q => coeff_memory_1_9);
   coeff_memory_reg_2_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n264,
                           CK => clk, RB => resetn, Q => coeff_memory_2_9);
   coeff_memory_reg_3_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n263,
                           CK => clk, RB => resetn, Q => coeff_memory_3_9);
   coeff_memory_reg_4_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n265,
                           CK => clk, RB => resetn, Q => coeff_memory_4_9);
   operand_regs_reg_2_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n258,
                           CK => clk, RB => resetn, Q => operand_regs_169_port)
                           ;
   operand_regs_reg_4_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n257,
                           CK => clk, RB => resetn, Q => operand_regs_105_port)
                           ;
   operand_regs_reg_6_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n256,
                           CK => clk, RB => resetn, Q => operand_regs_41_port);
   operand_regs_reg_0_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_239_port);
   operand_regs_reg_7_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n242,
                           CK => clk, RB => resetn, Q => operand_regs_0_port);
   operand_regs_reg_7_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_12_port);
   operand_regs_reg_0_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_236_port);
   operand_regs_reg_0_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n255,
                           CK => clk, RB => resetn, Q => operand_regs_233_port)
                           ;
   operand_regs_reg_7_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_10_port);
   operand_regs_reg_1_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n259,
                           CK => clk, RB => resetn, Q => operand_regs_196_port)
                           ;
   operand_regs_reg_1_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n259,
                           CK => clk, RB => resetn, Q => operand_regs_192_port)
                           ;
   coeff_memory_reg_0_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_11);
   coeff_memory_reg_1_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_11);
   coeff_memory_reg_2_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_11);
   coeff_memory_reg_3_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_11);
   coeff_memory_reg_4_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_11);
   operand_regs_reg_1_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n259,
                           CK => clk, RB => resetn, Q => operand_regs_195_port)
                           ;
   operand_regs_reg_2_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_171_port);
   operand_regs_reg_4_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_107_port);
   operand_regs_reg_6_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_43_port);
   operand_regs_reg_1_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_202_port);
   operand_regs_reg_7_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_11_port);
   operand_regs_reg_0_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_235_port);
   operand_regs_reg_1_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n259,
                           CK => clk, RB => resetn, Q => operand_regs_194_port)
                           ;
   operand_regs_reg_1_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n259,
                           CK => clk, RB => resetn, Q => operand_regs_193_port)
                           ;
   operand_regs_reg_7_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n242,
                           CK => clk, RB => resetn, Q => operand_regs_9_port);
   operand_regs_reg_1_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n259,
                           CK => clk, RB => resetn, Q => operand_regs_197_port)
                           ;
   operand_regs_reg_1_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n259,
                           CK => clk, RB => resetn, Q => operand_regs_201_port)
                           ;
   operand_regs_reg_1_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n259,
                           CK => clk, RB => resetn, Q => operand_regs_200_port)
                           ;
   operand_regs_reg_1_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n259,
                           CK => clk, RB => resetn, Q => operand_regs_199_port)
                           ;
   operand_regs_reg_1_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n259,
                           CK => clk, RB => resetn, Q => operand_regs_198_port)
                           ;
   coeff_memory_reg_0_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n267,
                           CK => clk, RB => resetn, Q => coeff_memory_0_8);
   coeff_memory_reg_1_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n266,
                           CK => clk, RB => resetn, Q => coeff_memory_1_8);
   coeff_memory_reg_2_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n264,
                           CK => clk, RB => resetn, Q => coeff_memory_2_8);
   coeff_memory_reg_3_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n263,
                           CK => clk, RB => resetn, Q => coeff_memory_3_8);
   coeff_memory_reg_4_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n265,
                           CK => clk, RB => resetn, Q => coeff_memory_4_8);
   operand_regs_reg_2_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n258,
                           CK => clk, RB => resetn, Q => operand_regs_168_port)
                           ;
   operand_regs_reg_4_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n257,
                           CK => clk, RB => resetn, Q => operand_regs_104_port)
                           ;
   operand_regs_reg_6_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n256,
                           CK => clk, RB => resetn, Q => operand_regs_40_port);
   coeff_memory_reg_0_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n267,
                           CK => clk, RB => resetn, Q => coeff_memory_0_4);
   coeff_memory_reg_1_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n266,
                           CK => clk, RB => resetn, Q => coeff_memory_1_4);
   coeff_memory_reg_2_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n264,
                           CK => clk, RB => resetn, Q => coeff_memory_2_4);
   coeff_memory_reg_3_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n263,
                           CK => clk, RB => resetn, Q => coeff_memory_3_4);
   coeff_memory_reg_4_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n265,
                           CK => clk, RB => resetn, Q => coeff_memory_4_4);
   operand_regs_reg_2_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n258,
                           CK => clk, RB => resetn, Q => operand_regs_164_port)
                           ;
   operand_regs_reg_4_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n257,
                           CK => clk, RB => resetn, Q => operand_regs_100_port)
                           ;
   operand_regs_reg_6_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n256,
                           CK => clk, RB => resetn, Q => operand_regs_36_port);
   operand_regs_reg_7_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n242,
                           CK => clk, RB => resetn, Q => operand_regs_8_port);
   operand_regs_reg_7_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n242,
                           CK => clk, RB => resetn, Q => operand_regs_4_port);
   operand_regs_reg_0_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n255,
                           CK => clk, RB => resetn, Q => operand_regs_232_port)
                           ;
   operand_regs_reg_0_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n255,
                           CK => clk, RB => resetn, Q => operand_regs_228_port)
                           ;
   coeff_memory_reg_0_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n267,
                           CK => clk, RB => resetn, Q => coeff_memory_0_6);
   coeff_memory_reg_1_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n266,
                           CK => clk, RB => resetn, Q => coeff_memory_1_6);
   coeff_memory_reg_2_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n264,
                           CK => clk, RB => resetn, Q => coeff_memory_2_6);
   coeff_memory_reg_3_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n263,
                           CK => clk, RB => resetn, Q => coeff_memory_3_6);
   coeff_memory_reg_4_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n265,
                           CK => clk, RB => resetn, Q => coeff_memory_4_6);
   operand_regs_reg_2_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n258,
                           CK => clk, RB => resetn, Q => operand_regs_166_port)
                           ;
   operand_regs_reg_4_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n257,
                           CK => clk, RB => resetn, Q => operand_regs_102_port)
                           ;
   operand_regs_reg_6_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n256,
                           CK => clk, RB => resetn, Q => operand_regs_38_port);
   operand_regs_reg_7_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n242,
                           CK => clk, RB => resetn, Q => operand_regs_6_port);
   operand_regs_reg_0_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n255,
                           CK => clk, RB => resetn, Q => operand_regs_230_port)
                           ;
   coeff_memory_reg_0_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n267,
                           CK => clk, RB => resetn, Q => coeff_memory_0_7);
   coeff_memory_reg_1_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n266,
                           CK => clk, RB => resetn, Q => coeff_memory_1_7);
   coeff_memory_reg_2_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n264,
                           CK => clk, RB => resetn, Q => coeff_memory_2_7);
   coeff_memory_reg_3_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n263,
                           CK => clk, RB => resetn, Q => coeff_memory_3_7);
   coeff_memory_reg_4_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n265,
                           CK => clk, RB => resetn, Q => coeff_memory_4_7);
   operand_regs_reg_2_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n258,
                           CK => clk, RB => resetn, Q => operand_regs_167_port)
                           ;
   operand_regs_reg_4_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n257,
                           CK => clk, RB => resetn, Q => operand_regs_103_port)
                           ;
   operand_regs_reg_6_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n256,
                           CK => clk, RB => resetn, Q => operand_regs_39_port);
   coeff_memory_reg_0_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n267,
                           CK => clk, RB => resetn, Q => coeff_memory_0_3);
   coeff_memory_reg_1_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n266,
                           CK => clk, RB => resetn, Q => coeff_memory_1_3);
   coeff_memory_reg_2_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n264,
                           CK => clk, RB => resetn, Q => coeff_memory_2_3);
   coeff_memory_reg_3_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n263,
                           CK => clk, RB => resetn, Q => coeff_memory_3_3);
   coeff_memory_reg_4_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n265,
                           CK => clk, RB => resetn, Q => coeff_memory_4_3);
   operand_regs_reg_2_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n258,
                           CK => clk, RB => resetn, Q => operand_regs_163_port)
                           ;
   operand_regs_reg_4_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n257,
                           CK => clk, RB => resetn, Q => operand_regs_99_port);
   operand_regs_reg_6_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n256,
                           CK => clk, RB => resetn, Q => operand_regs_35_port);
   coeff_memory_reg_0_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n267,
                           CK => clk, RB => resetn, Q => coeff_memory_0_2);
   coeff_memory_reg_1_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n266,
                           CK => clk, RB => resetn, Q => coeff_memory_1_2);
   coeff_memory_reg_2_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n264,
                           CK => clk, RB => resetn, Q => coeff_memory_2_2);
   coeff_memory_reg_3_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n263,
                           CK => clk, RB => resetn, Q => coeff_memory_3_2);
   coeff_memory_reg_4_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n265,
                           CK => clk, RB => resetn, Q => coeff_memory_4_2);
   operand_regs_reg_2_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n258,
                           CK => clk, RB => resetn, Q => operand_regs_162_port)
                           ;
   operand_regs_reg_4_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n257,
                           CK => clk, RB => resetn, Q => operand_regs_98_port);
   operand_regs_reg_6_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n256,
                           CK => clk, RB => resetn, Q => operand_regs_34_port);
   operand_regs_reg_7_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n242,
                           CK => clk, RB => resetn, Q => operand_regs_7_port);
   operand_regs_reg_7_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n242,
                           CK => clk, RB => resetn, Q => operand_regs_3_port);
   operand_regs_reg_0_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n255,
                           CK => clk, RB => resetn, Q => operand_regs_231_port)
                           ;
   operand_regs_reg_0_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n255,
                           CK => clk, RB => resetn, Q => operand_regs_227_port)
                           ;
   operand_regs_reg_7_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n242,
                           CK => clk, RB => resetn, Q => operand_regs_2_port);
   coeff_memory_reg_0_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n267,
                           CK => clk, RB => resetn, Q => coeff_memory_0_5);
   coeff_memory_reg_1_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n266,
                           CK => clk, RB => resetn, Q => coeff_memory_1_5);
   coeff_memory_reg_2_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n264,
                           CK => clk, RB => resetn, Q => coeff_memory_2_5);
   coeff_memory_reg_3_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n263,
                           CK => clk, RB => resetn, Q => coeff_memory_3_5);
   coeff_memory_reg_4_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n265,
                           CK => clk, RB => resetn, Q => coeff_memory_4_5);
   operand_regs_reg_2_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n258,
                           CK => clk, RB => resetn, Q => operand_regs_165_port)
                           ;
   operand_regs_reg_4_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n257,
                           CK => clk, RB => resetn, Q => operand_regs_101_port)
                           ;
   operand_regs_reg_6_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n256,
                           CK => clk, RB => resetn, Q => operand_regs_37_port);
   operand_regs_reg_0_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n255,
                           CK => clk, RB => resetn, Q => operand_regs_226_port)
                           ;
   operand_regs_reg_7_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n242,
                           CK => clk, RB => resetn, Q => operand_regs_5_port);
   operand_regs_reg_0_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n255,
                           CK => clk, RB => resetn, Q => operand_regs_229_port)
                           ;
   coeff_memory_reg_0_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n267,
                           CK => clk, RB => resetn, Q => coeff_memory_0_1);
   coeff_memory_reg_1_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n266,
                           CK => clk, RB => resetn, Q => coeff_memory_1_1);
   coeff_memory_reg_2_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n264,
                           CK => clk, RB => resetn, Q => coeff_memory_2_1);
   coeff_memory_reg_3_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n263,
                           CK => clk, RB => resetn, Q => coeff_memory_3_1);
   coeff_memory_reg_4_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n265,
                           CK => clk, RB => resetn, Q => coeff_memory_4_1);
   operand_regs_reg_2_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n258,
                           CK => clk, RB => resetn, Q => operand_regs_161_port)
                           ;
   operand_regs_reg_4_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n257,
                           CK => clk, RB => resetn, Q => operand_regs_97_port);
   operand_regs_reg_6_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n256,
                           CK => clk, RB => resetn, Q => operand_regs_33_port);
   operand_regs_reg_7_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n242,
                           CK => clk, RB => resetn, Q => operand_regs_1_port);
   operand_regs_reg_0_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n255,
                           CK => clk, RB => resetn, Q => operand_regs_225_port)
                           ;
   filt_mult_inputs_reg : DFERPQ1 port map( D => avs_writedata(0), CEB => n178,
                           CK => clk, RB => resetn, Q => filt_mult_inputs);
   siso_req_reg : DFERPQ1 port map( D => n806, CEB => n161, CK => clk, RB => 
                           resetn, Q => siso_req);
   siso_data_out_reg_0 : DFERPQ1 port map( D => N2888, CEB => n811, CK => clk, 
                           RB => resetn, Q => siso_data_out(0));
   siso_data_out_reg_15 : DFERPQ1 port map( D => N2903, CEB => n811, CK => clk,
                           RB => resetn, Q => siso_data_out(15));
   siso_data_out_reg_14 : DFERPQ1 port map( D => N2902, CEB => n811, CK => clk,
                           RB => resetn, Q => siso_data_out(14));
   siso_data_out_reg_13 : DFERPQ1 port map( D => N2901, CEB => n811, CK => clk,
                           RB => resetn, Q => siso_data_out(13));
   siso_data_out_reg_12 : DFERPQ1 port map( D => N2900, CEB => n811, CK => clk,
                           RB => resetn, Q => siso_data_out(12));
   siso_data_out_reg_11 : DFERPQ1 port map( D => N2899, CEB => n811, CK => clk,
                           RB => resetn, Q => siso_data_out(11));
   siso_data_out_reg_10 : DFERPQ1 port map( D => N2898, CEB => n811, CK => clk,
                           RB => resetn, Q => siso_data_out(10));
   siso_data_out_reg_9 : DFERPQ1 port map( D => N2897, CEB => n811, CK => clk, 
                           RB => resetn, Q => siso_data_out(9));
   siso_data_out_reg_8 : DFERPQ1 port map( D => N2896, CEB => n811, CK => clk, 
                           RB => resetn, Q => siso_data_out(8));
   siso_data_out_reg_7 : DFERPQ1 port map( D => N2895, CEB => n811, CK => clk, 
                           RB => resetn, Q => siso_data_out(7));
   siso_data_out_reg_6 : DFERPQ1 port map( D => N2894, CEB => n811, CK => clk, 
                           RB => resetn, Q => siso_data_out(6));
   siso_data_out_reg_5 : DFERPQ1 port map( D => N2893, CEB => n811, CK => clk, 
                           RB => resetn, Q => siso_data_out(5));
   siso_data_out_reg_4 : DFERPQ1 port map( D => N2892, CEB => n811, CK => clk, 
                           RB => resetn, Q => siso_data_out(4));
   siso_data_out_reg_3 : DFERPQ1 port map( D => N2891, CEB => n811, CK => clk, 
                           RB => resetn, Q => siso_data_out(3));
   siso_data_out_reg_2 : DFERPQ1 port map( D => N2890, CEB => n811, CK => clk, 
                           RB => resetn, Q => siso_data_out(2));
   siso_data_out_reg_1 : DFERPQ1 port map( D => N2889, CEB => n811, CK => clk, 
                           RB => resetn, Q => siso_data_out(1));
   siso_ready_reg : DFFRPQ1 port map( D => out_busy, CK => clk, RB => resetn, Q
                           => siso_ready);
   U642 : NAN3D1 port map( A1 => n309, A2 => avs_addr(0), A3 => n254, Z => n242
                           );
   U643 : AND2D1 port map( A1 => n313, A2 => avs_addr(0), Z => n243);
   U644 : AND2D1 port map( A1 => n561, A2 => N62, Z => n244);
   U645 : AND2D1 port map( A1 => n563, A2 => N62, Z => n245);
   U646 : NAN3D1 port map( A1 => n309, A2 => avs_addr(0), A3 => n110, Z => n246
                           );
   U647 : NAN2D1 port map( A1 => n110, A2 => n276, Z => n247);
   U648 : NAN2D1 port map( A1 => n110, A2 => n275, Z => n248);
   U649 : NAN2D1 port map( A1 => n110, A2 => n308, Z => n249);
   U650 : NAN2D1 port map( A1 => n110, A2 => n304, Z => n250);
   U651 : NAN2D1 port map( A1 => n110, A2 => n277, Z => n251);
   U652 : NAN2D1 port map( A1 => n110, A2 => n307, Z => n252);
   U653 : NAN2D1 port map( A1 => n110, A2 => n306, Z => n253);
   U654 : AND3D1 port map( A1 => operand_load, A2 => n104, A3 => n729, Z => 
                           n254);
   U655 : NAN2D1 port map( A1 => n275, A2 => n254, Z => n255);
   U656 : NAN2D1 port map( A1 => n277, A2 => n254, Z => n256);
   U657 : NAN2D1 port map( A1 => n276, A2 => n254, Z => n257);
   U658 : NAN2D1 port map( A1 => n307, A2 => n254, Z => n258);
   U659 : NAN2D1 port map( A1 => n308, A2 => n254, Z => n259);
   U660 : NAN2D1 port map( A1 => n304, A2 => n254, Z => n260);
   U661 : NAN2D1 port map( A1 => n306, A2 => n254, Z => n261);
   U662 : AND2D1 port map( A1 => n314, A2 => avs_addr(0), Z => n262);
   U663 : NAN2D1 port map( A1 => n306, A2 => n301, Z => n263);
   U664 : NAN2D1 port map( A1 => n307, A2 => n301, Z => n264);
   U665 : NAN2D1 port map( A1 => n276, A2 => n301, Z => n265);
   U666 : NAN2D1 port map( A1 => n308, A2 => n301, Z => n266);
   U667 : NAN2D1 port map( A1 => n275, A2 => n301, Z => n267);
   U668 : AND3D1 port map( A1 => N66, A2 => n300, A3 => read_comp_res, Z => 
                           n268);
   U669 : AND2D1 port map( A1 => n560, A2 => N62, Z => n269);
   U670 : AND2D1 port map( A1 => n562, A2 => N62, Z => n270);
   U671 : MUX2D1 port map( A0 => operand_regs_12_port, A1 => 
                           operand_regs_204_port, SL => n720, Z => n271);
   U672 : MUX2DL port map( A0 => operand_regs_13_port, A1 => 
                           operand_regs_205_port, SL => n719, Z => n272);
   U673 : MUX2DL port map( A0 => operand_regs_14_port, A1 => 
                           operand_regs_206_port, SL => n720, Z => n273);
   U674 : MUX2D1 port map( A0 => operand_regs_11_port, A1 => 
                           operand_regs_203_port, SL => n719, Z => n274);
   U675 : INVD1 port map( A => n724, Z => n710);
   U676 : INVD1 port map( A => n724, Z => n712);
   U677 : INVD1 port map( A => n724, Z => n711);
   U678 : INVD1 port map( A => n725, Z => n709);
   U679 : INVD1 port map( A => n725, Z => n707);
   U680 : INVD1 port map( A => n725, Z => n708);
   U681 : INVD1 port map( A => n726, Z => n706);
   U682 : INVD1 port map( A => n96, Z => n798);
   U683 : INVD1 port map( A => n702, Z => n724);
   U684 : INVD1 port map( A => n722, Z => n716);
   U685 : INVD1 port map( A => n723, Z => n714);
   U686 : INVD1 port map( A => n722, Z => n718);
   U687 : INVD1 port map( A => n723, Z => n715);
   U688 : INVD1 port map( A => n722, Z => n717);
   U689 : INVD1 port map( A => n702, Z => n725);
   U690 : INVD1 port map( A => n721, Z => n720);
   U691 : INVD1 port map( A => n721, Z => n719);
   U692 : INVD1 port map( A => n723, Z => n713);
   U693 : INVD1 port map( A => n702, Z => n726);
   U694 : INVD1 port map( A => n703, Z => n727);
   U695 : INVD1 port map( A => n703, Z => n728);
   U696 : INVD1 port map( A => n553, Z => n554);
   U697 : INVD1 port map( A => n558, Z => n559);
   U698 : INVD1 port map( A => n555, Z => n557);
   U699 : INVD1 port map( A => n555, Z => n556);
   U700 : INVD1 port map( A => n548, Z => n549);
   U701 : INVD1 port map( A => n548, Z => n550);
   U702 : INVD1 port map( A => n551, Z => n552);
   U703 : NAN2D1 port map( A1 => n275, A2 => n795, Z => n96);
   U704 : INVD1 port map( A => n74, Z => n797);
   U705 : NAN2D1 port map( A1 => n118, A2 => n807, Z => n176);
   U706 : NAN2D1 port map( A1 => n805, A2 => n118, Z => n174);
   U707 : INVD1 port map( A => n704, Z => n702);
   U708 : INVD1 port map( A => n701, Z => n722);
   U709 : INVD1 port map( A => n701, Z => n723);
   U710 : INVD1 port map( A => n701, Z => n721);
   U711 : INVD1 port map( A => n704, Z => n703);
   U712 : INVD1 port map( A => n300, Z => n700);
   U713 : INVD1 port map( A => n541, Z => n553);
   U714 : INVD1 port map( A => n543, Z => n558);
   U715 : INVD1 port map( A => n542, Z => n555);
   U716 : INVD1 port map( A => n699, Z => n698);
   U717 : INVD1 port map( A => n538, Z => n548);
   U718 : INVD1 port map( A => n539, Z => n551);
   U719 : OAI211D1 port map( A1 => n6300, A2 => n6400, B => n300, C => n65, Z 
                           => n14);
   U720 : NOR2D1 port map( A1 => n306, A2 => n307, Z => n6300);
   U721 : NOR3D1 port map( A1 => n797, A2 => N66, A3 => n798, Z => n65);
   U722 : INVD1 port map( A => n6400, Z => n795);
   U723 : NAN2D1 port map( A1 => n308, A2 => n795, Z => n74);
   U724 : AND3D1 port map( A1 => n796, A2 => n547, A3 => n762, Z => n275);
   U725 : AND2D1 port map( A1 => n111, A2 => n762, Z => n276);
   U726 : AND2D1 port map( A1 => n309, A2 => n762, Z => n277);
   U727 : NOR3D1 port map( A1 => n813, A2 => n810, A3 => n696, Z => n78);
   U728 : INVD1 port map( A => n81, Z => n801);
   U729 : INVD1 port map( A => n697, Z => n812);
   U730 : NOR2D1 port map( A1 => n809, A2 => n803, Z => n118);
   U731 : INVD1 port map( A => n88, Z => n807);
   U732 : NOR2D1 port map( A1 => n800, A2 => n91, Z => n89);
   U733 : INVD1 port map( A => n84, Z => n800);
   U734 : INVD1 port map( A => n155, Z => n804);
   U735 : NAN2D1 port map( A1 => n119, A2 => n115, Z => n171);
   U736 : NAN2D1 port map( A1 => n119, A2 => n101, Z => n162);
   U737 : NAN2D1 port map( A1 => n119, A2 => n118, Z => n170);
   U738 : NAN2D1 port map( A1 => n120, A2 => n119, Z => n163);
   U739 : NAN2D1 port map( A1 => n87, A2 => n84, Z => n86);
   U740 : NAN2D1 port map( A1 => n805, A2 => n101, Z => n166);
   U741 : INVD1 port map( A => n85, Z => n805);
   U742 : NAN2D1 port map( A1 => n120, A2 => n805, Z => n167);
   U743 : NAN2D1 port map( A1 => n805, A2 => n115, Z => n175);
   U744 : NAN2D1 port map( A1 => n87, A2 => n101, Z => n164);
   U745 : NAN2D1 port map( A1 => n115, A2 => n87, Z => n173);
   U746 : NAN2D1 port map( A1 => n120, A2 => n87, Z => n165);
   U747 : NAN2D1 port map( A1 => n118, A2 => n87, Z => n172);
   U748 : NAN2D1 port map( A1 => n807, A2 => n101, Z => n168);
   U749 : NAN2D1 port map( A1 => n115, A2 => n807, Z => n177);
   U750 : NAN2D1 port map( A1 => n120, A2 => n807, Z => n169);
   U751 : MUX2DL port map( A0 => operand_regs_33_port, A1 => coeff_memory_3_1, 
                           SL => n712, Z => N3010);
   U752 : MUX2DL port map( A0 => operand_regs_97_port, A1 => coeff_memory_2_1, 
                           SL => n710, Z => N2978);
   U753 : INVD1 port map( A => filt_mult_inputs, Z => n704);
   U754 : MUX2DL port map( A0 => operand_regs_1_port, A1 => coeff_memory_4_1, 
                           SL => n714, Z => N3042);
   U755 : MUX2DL port map( A0 => operand_regs_161_port, A1 => coeff_memory_1_1,
                           SL => n718, Z => N2946);
   U756 : MUX2DL port map( A0 => operand_regs_225_port, A1 => coeff_memory_0_1,
                           SL => n716, Z => N2914);
   U757 : INVD1 port map( A => n705, Z => n701);
   U758 : INVD1 port map( A => filt_mult_inputs, Z => n705);
   U759 : MUX2DL port map( A0 => operand_regs_37_port, A1 => coeff_memory_3_5, 
                           SL => n712, Z => N3014);
   U760 : MUX2DL port map( A0 => operand_regs_101_port, A1 => coeff_memory_2_5,
                           SL => n711, Z => N2982);
   U761 : MUX2DL port map( A0 => operand_regs_5_port, A1 => coeff_memory_4_5, 
                           SL => n714, Z => N3046);
   U762 : MUX2DL port map( A0 => operand_regs_165_port, A1 => coeff_memory_1_5,
                           SL => n718, Z => N2950);
   U763 : MUX2DL port map( A0 => operand_regs_229_port, A1 => coeff_memory_0_5,
                           SL => n715, Z => N2918);
   U764 : MUX2DL port map( A0 => operand_regs_34_port, A1 => coeff_memory_3_2, 
                           SL => n712, Z => N3011);
   U765 : MUX2DL port map( A0 => operand_regs_98_port, A1 => coeff_memory_2_2, 
                           SL => n710, Z => N2979);
   U766 : MUX2DL port map( A0 => operand_regs_35_port, A1 => coeff_memory_3_3, 
                           SL => n712, Z => N3012);
   U767 : MUX2DL port map( A0 => operand_regs_99_port, A1 => coeff_memory_2_3, 
                           SL => n710, Z => N2980);
   U768 : MUX2DL port map( A0 => operand_regs_2_port, A1 => coeff_memory_4_2, 
                           SL => n714, Z => N3043);
   U769 : MUX2DL port map( A0 => operand_regs_162_port, A1 => coeff_memory_1_2,
                           SL => n717, Z => N2947);
   U770 : MUX2DL port map( A0 => operand_regs_226_port, A1 => coeff_memory_0_2,
                           SL => n716, Z => N2915);
   U771 : MUX2DL port map( A0 => operand_regs_39_port, A1 => coeff_memory_3_7, 
                           SL => n712, Z => N3016);
   U772 : MUX2DL port map( A0 => operand_regs_103_port, A1 => coeff_memory_2_7,
                           SL => n711, Z => N2984);
   U773 : MUX2DL port map( A0 => operand_regs_3_port, A1 => coeff_memory_4_3, 
                           SL => n714, Z => N3044);
   U774 : MUX2DL port map( A0 => operand_regs_163_port, A1 => coeff_memory_1_3,
                           SL => n718, Z => N2948);
   U775 : MUX2DL port map( A0 => operand_regs_227_port, A1 => coeff_memory_0_3,
                           SL => n716, Z => N2916);
   U776 : MUX2DL port map( A0 => operand_regs_7_port, A1 => coeff_memory_4_7, 
                           SL => n714, Z => N3048);
   U777 : MUX2DL port map( A0 => operand_regs_167_port, A1 => coeff_memory_1_7,
                           SL => n718, Z => N2952);
   U778 : MUX2DL port map( A0 => operand_regs_231_port, A1 => coeff_memory_0_7,
                           SL => n715, Z => N2920);
   U779 : MUX2DL port map( A0 => operand_regs_38_port, A1 => coeff_memory_3_6, 
                           SL => n712, Z => N3015);
   U780 : MUX2DL port map( A0 => operand_regs_102_port, A1 => coeff_memory_2_6,
                           SL => n711, Z => N2983);
   U781 : MUX2DL port map( A0 => operand_regs_6_port, A1 => coeff_memory_4_6, 
                           SL => n714, Z => N3047);
   U782 : MUX2DL port map( A0 => operand_regs_166_port, A1 => coeff_memory_1_6,
                           SL => n717, Z => N2951);
   U783 : MUX2DL port map( A0 => operand_regs_230_port, A1 => coeff_memory_0_6,
                           SL => n715, Z => N2919);
   U784 : MUX2DL port map( A0 => operand_regs_36_port, A1 => coeff_memory_3_4, 
                           SL => n712, Z => N3013);
   U785 : MUX2DL port map( A0 => operand_regs_100_port, A1 => coeff_memory_2_4,
                           SL => n711, Z => N2981);
   U786 : MUX2DL port map( A0 => operand_regs_104_port, A1 => coeff_memory_2_8,
                           SL => n711, Z => N2985);
   U787 : MUX2DL port map( A0 => operand_regs_40_port, A1 => coeff_memory_3_8, 
                           SL => n709, Z => N3017);
   U788 : MUX2DL port map( A0 => operand_regs_4_port, A1 => coeff_memory_4_4, 
                           SL => n714, Z => N3045);
   U789 : MUX2DL port map( A0 => operand_regs_164_port, A1 => coeff_memory_1_4,
                           SL => n717, Z => N2949);
   U790 : MUX2DL port map( A0 => operand_regs_228_port, A1 => coeff_memory_0_4,
                           SL => n716, Z => N2917);
   U791 : MUX2DL port map( A0 => operand_regs_8_port, A1 => coeff_memory_4_8, 
                           SL => n714, Z => N3049);
   U792 : MUX2DL port map( A0 => operand_regs_168_port, A1 => coeff_memory_1_8,
                           SL => n717, Z => N2953);
   U793 : MUX2DL port map( A0 => operand_regs_232_port, A1 => coeff_memory_0_8,
                           SL => n715, Z => N2921);
   U794 : MUX2DL port map( A0 => operand_regs_6_port, A1 => 
                           operand_regs_198_port, SL => n720, Z => n278);
   U795 : MUX2DL port map( A0 => operand_regs_7_port, A1 => 
                           operand_regs_199_port, SL => n719, Z => n279);
   U796 : MUX2DL port map( A0 => operand_regs_43_port, A1 => coeff_memory_3_11,
                           SL => n711, Z => N3020);
   U797 : MUX2DL port map( A0 => operand_regs_107_port, A1 => coeff_memory_2_11
                           , SL => n711, Z => N2988);
   U798 : MUX2DL port map( A0 => operand_regs_8_port, A1 => 
                           operand_regs_200_port, SL => n720, Z => n280);
   U799 : MUX2DL port map( A0 => operand_regs_11_port, A1 => coeff_memory_4_11,
                           SL => n713, Z => N3052);
   U800 : MUX2DL port map( A0 => operand_regs_171_port, A1 => coeff_memory_1_11
                           , SL => n718, Z => N2956);
   U801 : MUX2DL port map( A0 => operand_regs_235_port, A1 => coeff_memory_0_11
                           , SL => n715, Z => N2924);
   U802 : MUX2DL port map( A0 => operand_regs_9_port, A1 => 
                           operand_regs_201_port, SL => n719, Z => n281);
   U803 : MUX2DL port map( A0 => operand_regs_5_port, A1 => 
                           operand_regs_197_port, SL => n719, Z => n282);
   U804 : MUX2DL port map( A0 => operand_regs_1_port, A1 => 
                           operand_regs_193_port, SL => n720, Z => n283);
   U805 : MUX2DL port map( A0 => operand_regs_2_port, A1 => 
                           operand_regs_194_port, SL => n720, Z => n284);
   U806 : MUX2DL port map( A0 => operand_regs_44_port, A1 => coeff_memory_3_12,
                           SL => n711, Z => N3021);
   U807 : MUX2DL port map( A0 => operand_regs_108_port, A1 => coeff_memory_2_12
                           , SL => n711, Z => N2989);
   U808 : MUX2DL port map( A0 => operand_regs_10_port, A1 => 
                           operand_regs_202_port, SL => n720, Z => n285);
   U809 : MUX2DL port map( A0 => operand_regs_41_port, A1 => coeff_memory_3_9, 
                           SL => n712, Z => N3018);
   U810 : MUX2DL port map( A0 => operand_regs_105_port, A1 => coeff_memory_2_9,
                           SL => n711, Z => N2986);
   U811 : MUX2DL port map( A0 => operand_regs_12_port, A1 => coeff_memory_4_12,
                           SL => n713, Z => N3053);
   U812 : MUX2DL port map( A0 => operand_regs_172_port, A1 => coeff_memory_1_12
                           , SL => n717, Z => N2957);
   U813 : MUX2DL port map( A0 => operand_regs_236_port, A1 => coeff_memory_0_12
                           , SL => n715, Z => N2925);
   U814 : MUX2DL port map( A0 => operand_regs_9_port, A1 => coeff_memory_4_9, 
                           SL => n713, Z => N3050);
   U815 : MUX2DL port map( A0 => operand_regs_169_port, A1 => coeff_memory_1_9,
                           SL => n718, Z => N2954);
   U816 : MUX2DL port map( A0 => operand_regs_233_port, A1 => coeff_memory_0_9,
                           SL => n715, Z => N2922);
   U817 : MUX2DL port map( A0 => operand_regs_3_port, A1 => 
                           operand_regs_195_port, SL => n720, Z => n286);
   U818 : MUX2DL port map( A0 => operand_regs_45_port, A1 => coeff_memory_3_13,
                           SL => n711, Z => N3022);
   U819 : MUX2DL port map( A0 => operand_regs_109_port, A1 => coeff_memory_2_13
                           , SL => n711, Z => N2990);
   U820 : MUX2DL port map( A0 => operand_regs_47_port, A1 => coeff_memory_3_15,
                           SL => n711, Z => N3024);
   U821 : MUX2DL port map( A0 => operand_regs_111_port, A1 => coeff_memory_2_15
                           , SL => n712, Z => N2992);
   U822 : MUX2DL port map( A0 => operand_regs_4_port, A1 => 
                           operand_regs_196_port, SL => n720, Z => n287);
   U823 : MUX2DL port map( A0 => operand_regs_13_port, A1 => coeff_memory_4_13,
                           SL => n713, Z => N3054);
   U824 : MUX2DL port map( A0 => operand_regs_173_port, A1 => coeff_memory_1_13
                           , SL => n718, Z => N2958);
   U825 : MUX2DL port map( A0 => operand_regs_237_port, A1 => coeff_memory_0_13
                           , SL => n715, Z => N2926);
   U826 : MUX2DL port map( A0 => operand_regs_15_port, A1 => coeff_memory_4_15,
                           SL => n713, Z => N3056);
   U827 : MUX2DL port map( A0 => operand_regs_175_port, A1 => coeff_memory_1_15
                           , SL => n718, Z => N2960);
   U828 : MUX2DL port map( A0 => operand_regs_239_port, A1 => coeff_memory_0_15
                           , SL => n715, Z => N2928);
   U829 : MUX2DL port map( A0 => operand_regs_192_port, A1 => 
                           operand_regs_0_port, SL => n721, Z => n288);
   U830 : INVD1 port map( A => operand_regs_198_port, Z => n755);
   U831 : INVD1 port map( A => operand_regs_199_port, Z => n754);
   U832 : MUX2DL port map( A0 => operand_regs_46_port, A1 => coeff_memory_3_14,
                           SL => n711, Z => N3023);
   U833 : MUX2DL port map( A0 => operand_regs_110_port, A1 => coeff_memory_2_14
                           , SL => n711, Z => N2991);
   U834 : INVD1 port map( A => operand_regs_200_port, Z => n753);
   U835 : MUX2DL port map( A0 => operand_regs_14_port, A1 => coeff_memory_4_14,
                           SL => n713, Z => N3055);
   U836 : MUX2DL port map( A0 => operand_regs_174_port, A1 => coeff_memory_1_14
                           , SL => n717, Z => N2959);
   U837 : MUX2DL port map( A0 => operand_regs_238_port, A1 => coeff_memory_0_14
                           , SL => n715, Z => N2927);
   U838 : INVD1 port map( A => operand_regs_194_port, Z => n759);
   U839 : INVD1 port map( A => operand_regs_193_port, Z => n760);
   U840 : INVD1 port map( A => operand_regs_197_port, Z => n756);
   U841 : MUX2DL port map( A0 => operand_regs_48_port, A1 => coeff_memory_3_16,
                           SL => n709, Z => N3025);
   U842 : MUX2DL port map( A0 => operand_regs_16_port, A1 => coeff_memory_4_16,
                           SL => n713, Z => N3057);
   U843 : MUX2DL port map( A0 => operand_regs_112_port, A1 => coeff_memory_2_16
                           , SL => n717, Z => N2993);
   U844 : MUX2DL port map( A0 => operand_regs_176_port, A1 => coeff_memory_1_16
                           , SL => n717, Z => N2961);
   U845 : MUX2DL port map( A0 => operand_regs_240_port, A1 => coeff_memory_0_16
                           , SL => n715, Z => N2929);
   U846 : MUX2DL port map( A0 => operand_regs_49_port, A1 => coeff_memory_3_17,
                           SL => n709, Z => N3026);
   U847 : MUX2DL port map( A0 => operand_regs_17_port, A1 => coeff_memory_4_17,
                           SL => n713, Z => N3058);
   U848 : MUX2DL port map( A0 => operand_regs_113_port, A1 => coeff_memory_2_17
                           , SL => n719, Z => N2994);
   U849 : MUX2DL port map( A0 => operand_regs_177_port, A1 => coeff_memory_1_17
                           , SL => n717, Z => N2962);
   U850 : MUX2DL port map( A0 => operand_regs_241_port, A1 => coeff_memory_0_17
                           , SL => n715, Z => N2930);
   U851 : MUX2DL port map( A0 => operand_regs_42_port, A1 => coeff_memory_3_10,
                           SL => n711, Z => N3019);
   U852 : MUX2DL port map( A0 => operand_regs_106_port, A1 => coeff_memory_2_10
                           , SL => n711, Z => N2987);
   U853 : INVD1 port map( A => operand_regs_195_port, Z => n758);
   U854 : MUX2DL port map( A0 => operand_regs_10_port, A1 => coeff_memory_4_10,
                           SL => n713, Z => N3051);
   U855 : MUX2DL port map( A0 => operand_regs_170_port, A1 => coeff_memory_1_10
                           , SL => n717, Z => N2955);
   U856 : MUX2DL port map( A0 => operand_regs_234_port, A1 => coeff_memory_0_10
                           , SL => n715, Z => N2923);
   U857 : INVD1 port map( A => operand_regs_192_port, Z => n761);
   U858 : INVD1 port map( A => operand_regs_196_port, Z => n757);
   U859 : MUX2DL port map( A0 => operand_regs_50_port, A1 => coeff_memory_3_18,
                           SL => n709, Z => N3027);
   U860 : MUX2DL port map( A0 => operand_regs_18_port, A1 => coeff_memory_4_18,
                           SL => n713, Z => N3059);
   U861 : MUX2DL port map( A0 => operand_regs_114_port, A1 => coeff_memory_2_18
                           , SL => n718, Z => N2995);
   U862 : MUX2DL port map( A0 => operand_regs_178_port, A1 => coeff_memory_1_18
                           , SL => n717, Z => N2963);
   U863 : MUX2DL port map( A0 => operand_regs_242_port, A1 => coeff_memory_0_18
                           , SL => n715, Z => N2931);
   U864 : INVD1 port map( A => operand_regs_201_port, Z => n752);
   U865 : MUX2DL port map( A0 => operand_regs_96_port, A1 => coeff_memory_2_0, 
                           SL => n710, Z => N2977);
   U866 : MUX2DL port map( A0 => operand_regs_51_port, A1 => coeff_memory_3_19,
                           SL => n710, Z => N3028);
   U867 : MUX2DL port map( A0 => operand_regs_32_port, A1 => coeff_memory_3_0, 
                           SL => n712, Z => N3009);
   U868 : MUX2DL port map( A0 => operand_regs_160_port, A1 => coeff_memory_1_0,
                           SL => n717, Z => N2945);
   U869 : MUX2DL port map( A0 => operand_regs_19_port, A1 => coeff_memory_4_19,
                           SL => n713, Z => N3060);
   U870 : MUX2DL port map( A0 => operand_regs_115_port, A1 => coeff_memory_2_19
                           , SL => n719, Z => N2996);
   U871 : MUX2DL port map( A0 => operand_regs_179_port, A1 => coeff_memory_1_19
                           , SL => n717, Z => N2964);
   U872 : MUX2DL port map( A0 => operand_regs_243_port, A1 => coeff_memory_0_19
                           , SL => n715, Z => N2932);
   U873 : MUX2DL port map( A0 => operand_regs_224_port, A1 => coeff_memory_0_0,
                           SL => n716, Z => N2913);
   U874 : MUX2DL port map( A0 => operand_regs_0_port, A1 => coeff_memory_4_0, 
                           SL => n714, Z => N3041);
   U875 : INVD1 port map( A => operand_regs_202_port, Z => n751);
   U876 : MUX2DL port map( A0 => operand_regs_17_port, A1 => 
                           operand_regs_209_port, SL => n719, Z => n289);
   U877 : MUX2DL port map( A0 => operand_regs_18_port, A1 => 
                           operand_regs_210_port, SL => n720, Z => n290);
   U878 : INVD1 port map( A => operand_regs_204_port, Z => n749);
   U879 : MUX2DL port map( A0 => operand_regs_15_port, A1 => 
                           operand_regs_207_port, SL => n719, Z => n291);
   U880 : INVD1 port map( A => operand_regs_203_port, Z => n750);
   U881 : MUX2DL port map( A0 => operand_regs_16_port, A1 => 
                           operand_regs_208_port, SL => n720, Z => n292);
   U882 : MUX2DL port map( A0 => operand_regs_52_port, A1 => coeff_memory_3_20,
                           SL => n710, Z => N3029);
   U883 : INVD1 port map( A => operand_regs_205_port, Z => n748);
   U884 : MUX2DL port map( A0 => operand_regs_20_port, A1 => coeff_memory_4_20,
                           SL => n713, Z => N3061);
   U885 : MUX2DL port map( A0 => operand_regs_116_port, A1 => coeff_memory_2_20
                           , SL => n718, Z => N2997);
   U886 : MUX2DL port map( A0 => operand_regs_180_port, A1 => coeff_memory_1_20
                           , SL => n717, Z => N2965);
   U887 : MUX2DL port map( A0 => operand_regs_244_port, A1 => coeff_memory_0_20
                           , SL => n715, Z => N2933);
   U888 : INVD1 port map( A => operand_regs_206_port, Z => n747);
   U889 : INVD1 port map( A => operand_regs_209_port, Z => n744);
   U890 : MUX2DL port map( A0 => operand_regs_19_port, A1 => 
                           operand_regs_211_port, SL => n719, Z => n293);
   U891 : INVD1 port map( A => operand_regs_207_port, Z => n746);
   U892 : MUX2DL port map( A0 => operand_regs_20_port, A1 => 
                           operand_regs_212_port, SL => n720, Z => n294);
   U893 : INVD1 port map( A => operand_regs_210_port, Z => n743);
   U894 : INVD1 port map( A => operand_regs_208_port, Z => n745);
   U895 : INVD1 port map( A => operand_regs_211_port, Z => n742);
   U896 : INVD1 port map( A => operand_regs_212_port, Z => n741);
   U897 : MUX2DL port map( A0 => operand_regs_53_port, A1 => coeff_memory_3_21,
                           SL => n710, Z => N3030);
   U898 : MUX2DL port map( A0 => operand_regs_21_port, A1 => coeff_memory_4_21,
                           SL => n713, Z => N3062);
   U899 : MUX2DL port map( A0 => operand_regs_117_port, A1 => coeff_memory_2_21
                           , SL => n719, Z => N2998);
   U900 : MUX2DL port map( A0 => operand_regs_181_port, A1 => coeff_memory_1_21
                           , SL => n716, Z => N2966);
   U901 : MUX2DL port map( A0 => operand_regs_245_port, A1 => coeff_memory_0_21
                           , SL => n715, Z => N2934);
   U902 : MUX2DL port map( A0 => operand_regs_21_port, A1 => 
                           operand_regs_213_port, SL => n719, Z => n295);
   U903 : MUX2DL port map( A0 => operand_regs_54_port, A1 => coeff_memory_3_22,
                           SL => n710, Z => N3031);
   U904 : MUX2DL port map( A0 => operand_regs_22_port, A1 => coeff_memory_4_22,
                           SL => n713, Z => N3063);
   U905 : MUX2DL port map( A0 => operand_regs_118_port, A1 => coeff_memory_2_22
                           , SL => n717, Z => N2999);
   U906 : MUX2DL port map( A0 => operand_regs_182_port, A1 => coeff_memory_1_22
                           , SL => n716, Z => N2967);
   U907 : MUX2DL port map( A0 => operand_regs_246_port, A1 => coeff_memory_0_22
                           , SL => n714, Z => N2935);
   U908 : MUX2DL port map( A0 => operand_regs_22_port, A1 => 
                           operand_regs_214_port, SL => n720, Z => n296);
   U909 : INVD1 port map( A => operand_regs_213_port, Z => n740);
   U910 : INVD1 port map( A => operand_regs_214_port, Z => n739);
   U911 : MUX2DL port map( A0 => operand_regs_55_port, A1 => coeff_memory_3_23,
                           SL => n710, Z => N3032);
   U912 : MUX2DL port map( A0 => operand_regs_23_port, A1 => coeff_memory_4_23,
                           SL => n713, Z => N3064);
   U913 : MUX2DL port map( A0 => operand_regs_119_port, A1 => coeff_memory_2_23
                           , SL => n718, Z => N3000);
   U914 : MUX2DL port map( A0 => operand_regs_183_port, A1 => coeff_memory_1_23
                           , SL => n716, Z => N2968);
   U915 : MUX2DL port map( A0 => operand_regs_247_port, A1 => coeff_memory_0_23
                           , SL => n714, Z => N2936);
   U916 : MUX2DL port map( A0 => operand_regs_56_port, A1 => coeff_memory_3_24,
                           SL => n710, Z => N3033);
   U917 : MUX2DL port map( A0 => operand_regs_24_port, A1 => coeff_memory_4_24,
                           SL => n713, Z => N3065);
   U918 : MUX2DL port map( A0 => operand_regs_120_port, A1 => coeff_memory_2_24
                           , SL => n718, Z => N3001);
   U919 : MUX2DL port map( A0 => operand_regs_184_port, A1 => coeff_memory_1_24
                           , SL => n716, Z => N2969);
   U920 : MUX2DL port map( A0 => operand_regs_248_port, A1 => coeff_memory_0_24
                           , SL => n714, Z => N2937);
   U921 : MUX2DL port map( A0 => operand_regs_23_port, A1 => 
                           operand_regs_215_port, SL => n719, Z => n297);
   U922 : INVD1 port map( A => operand_regs_215_port, Z => n738);
   U923 : MUX2DL port map( A0 => operand_regs_57_port, A1 => coeff_memory_3_25,
                           SL => n710, Z => N3034);
   U924 : MUX2DL port map( A0 => operand_regs_25_port, A1 => coeff_memory_4_25,
                           SL => n713, Z => N3066);
   U925 : MUX2DL port map( A0 => operand_regs_121_port, A1 => coeff_memory_2_25
                           , SL => n718, Z => N3002);
   U926 : MUX2DL port map( A0 => operand_regs_185_port, A1 => coeff_memory_1_25
                           , SL => n716, Z => N2970);
   U927 : MUX2DL port map( A0 => operand_regs_249_port, A1 => coeff_memory_0_25
                           , SL => n714, Z => N2938);
   U928 : NOR3M1D1 port map( A1 => n104, A2 => coeff_load, A3 => operand_load, 
                           Z => n110);
   U929 : AND2D1 port map( A1 => N66, A2 => avs_write, Z => n104);
   U930 : MUX2DL port map( A0 => operand_regs_24_port, A1 => 
                           operand_regs_216_port, SL => n720, Z => n298);
   U931 : INVD1 port map( A => operand_regs_216_port, Z => n737);
   U932 : MUX2DL port map( A0 => operand_regs_25_port, A1 => 
                           operand_regs_217_port, SL => n719, Z => n299);
   U933 : MUX2DL port map( A0 => operand_regs_26_port, A1 => coeff_memory_4_26,
                           SL => n712, Z => N3067);
   U934 : MUX2DL port map( A0 => operand_regs_58_port, A1 => coeff_memory_3_26,
                           SL => n710, Z => N3035);
   U935 : MUX2DL port map( A0 => operand_regs_122_port, A1 => coeff_memory_2_26
                           , SL => n718, Z => N3003);
   U936 : MUX2DL port map( A0 => operand_regs_186_port, A1 => coeff_memory_1_26
                           , SL => n716, Z => N2971);
   U937 : MUX2DL port map( A0 => operand_regs_250_port, A1 => coeff_memory_0_26
                           , SL => n714, Z => N2939);
   U938 : INVD1 port map( A => coeff_load, Z => n729);
   U939 : INVD1 port map( A => operand_regs_217_port, Z => n736);
   U940 : NAN4D1 port map( A1 => n5900, A2 => n14, A3 => n6000, A4 => n6100, Z 
                           => n233);
   U941 : NAN2M1D1 port map( A1 => n70, A2 => n300, Z => n5900);
   U942 : NAN2D1 port map( A1 => N2009, A2 => n268, Z => n6000);
   U943 : INVD1 port map( A => avs_write, Z => n799);
   U944 : AND2D1 port map( A1 => avs_read, A2 => n799, Z => n300);
   U945 : INVD1 port map( A => n12, Z => n699);
   U946 : NOR3M1D1 port map( A1 => N66, A2 => n700, A3 => read_comp_res, Z => 
                           n12);
   U947 : NAN3D1 port map( A1 => n56, A2 => n14, A3 => n57, Z => n231);
   U948 : NAN2D1 port map( A1 => N2007, A2 => n268, Z => n56);
   U949 : NAN3D1 port map( A1 => n452, A2 => n451, A3 => n453, Z => N2007);
   U950 : NAN3D1 port map( A1 => n53, A2 => n14, A3 => n54, Z => n229);
   U951 : NAN2D1 port map( A1 => N2005, A2 => n268, Z => n53);
   U952 : NAN3D1 port map( A1 => n458, A2 => n457, A3 => n459, Z => N2005);
   U953 : NAN3D1 port map( A1 => n50, A2 => n14, A3 => n51, Z => n227);
   U954 : NAN2D1 port map( A1 => N2003, A2 => n268, Z => n50);
   U955 : NAN3D1 port map( A1 => n464, A2 => n463, A3 => n465, Z => N2003);
   U956 : NAN3D1 port map( A1 => n47, A2 => n14, A3 => n48, Z => n225);
   U957 : NAN2D1 port map( A1 => N2001, A2 => n268, Z => n47);
   U958 : NAN3D1 port map( A1 => n470, A2 => n469, A3 => n471, Z => N2001);
   U959 : NAN3D1 port map( A1 => n44, A2 => n14, A3 => n45, Z => n223);
   U960 : NAN2D1 port map( A1 => N1999, A2 => n268, Z => n44);
   U961 : NAN3D1 port map( A1 => n476, A2 => n475, A3 => n477, Z => N1999);
   U962 : NAN3D1 port map( A1 => n41, A2 => n14, A3 => n42, Z => n221);
   U963 : NAN2D1 port map( A1 => N1997, A2 => n268, Z => n41);
   U964 : NAN3D1 port map( A1 => n482, A2 => n481, A3 => n483, Z => N1997);
   U965 : NAN3D1 port map( A1 => n38, A2 => n14, A3 => n39, Z => n219);
   U966 : NAN2D1 port map( A1 => N1995, A2 => n268, Z => n38);
   U967 : NAN3D1 port map( A1 => n488, A2 => n487, A3 => n489, Z => N1995);
   U968 : NAN3D1 port map( A1 => n35, A2 => n14, A3 => n36, Z => n217);
   U969 : NAN2D1 port map( A1 => N1993, A2 => n268, Z => n35);
   U970 : NAN3D1 port map( A1 => n494, A2 => n493, A3 => n495, Z => N1993);
   U971 : NAN3D1 port map( A1 => n13, A2 => n14, A3 => n15, Z => n203);
   U972 : NAN2D1 port map( A1 => N1979, A2 => n268, Z => n13);
   U973 : NAN3D1 port map( A1 => n536, A2 => n535, A3 => n537, Z => N1979);
   U974 : INVD1 port map( A => avs_addr(2), Z => n547);
   U975 : NAN3D1 port map( A1 => n32, A2 => n14, A3 => n33, Z => n215);
   U976 : NAN2D1 port map( A1 => N1991, A2 => n268, Z => n32);
   U977 : NAN3D1 port map( A1 => n500, A2 => n499, A3 => n501, Z => N1991);
   U978 : NAN3D1 port map( A1 => n29, A2 => n14, A3 => n30, Z => n213);
   U979 : NAN2D1 port map( A1 => N1989, A2 => n268, Z => n29);
   U980 : NAN3D1 port map( A1 => n506, A2 => n505, A3 => n507, Z => N1989);
   U981 : NAN3D1 port map( A1 => n26, A2 => n14, A3 => n27, Z => n211);
   U982 : NAN2D1 port map( A1 => N1987, A2 => n268, Z => n26);
   U983 : NAN3D1 port map( A1 => n512, A2 => n511, A3 => n513, Z => N1987);
   U984 : NAN3D1 port map( A1 => n23, A2 => n14, A3 => n24, Z => n209);
   U985 : NAN2D1 port map( A1 => N1985, A2 => n268, Z => n23);
   U986 : NAN3D1 port map( A1 => n518, A2 => n517, A3 => n519, Z => N1985);
   U987 : NAN3D1 port map( A1 => n20, A2 => n14, A3 => n21, Z => n207);
   U988 : NAN2D1 port map( A1 => N1983, A2 => n268, Z => n20);
   U989 : NAN3D1 port map( A1 => n524, A2 => n523, A3 => n525, Z => N1983);
   U990 : NAN3D1 port map( A1 => n17, A2 => n14, A3 => n18, Z => n205);
   U991 : NAN2D1 port map( A1 => N1981, A2 => n268, Z => n17);
   U992 : NAN3D1 port map( A1 => n530, A2 => n529, A3 => n531, Z => N1981);
   U993 : OAI21M20D1 port map( A1 => avs_readdata_1_port, A2 => n700, B => n58,
                           Z => n232);
   U994 : NAN3D1 port map( A1 => n449, A2 => n448, A3 => n450, Z => N2008);
   U995 : OAI21M20D1 port map( A1 => avs_readdata_3_port, A2 => n700, B => n55,
                           Z => n230);
   U996 : NAN3D1 port map( A1 => n455, A2 => n454, A3 => n456, Z => N2006);
   U997 : OAI21M20D1 port map( A1 => avs_readdata_5_port, A2 => n700, B => n52,
                           Z => n228);
   U998 : NAN3D1 port map( A1 => n461, A2 => n460, A3 => n462, Z => N2004);
   U999 : OAI21M20D1 port map( A1 => avs_readdata_7_port, A2 => n700, B => n49,
                           Z => n226);
   U1000 : NAN3D1 port map( A1 => n467, A2 => n466, A3 => n468, Z => N2002);
   U1001 : OAI21M20D1 port map( A1 => avs_readdata_15_port, A2 => n700, B => 
                           n37, Z => n218);
   U1002 : NAN3D1 port map( A1 => n491, A2 => n490, A3 => n492, Z => N1994);
   U1003 : OAI21M20D1 port map( A1 => avs_readdata_17_port, A2 => n700, B => 
                           n34, Z => n216);
   U1004 : NAN3D1 port map( A1 => n497, A2 => n496, A3 => n498, Z => N1992);
   U1005 : OAI21M20D1 port map( A1 => avs_readdata_19_port, A2 => n700, B => 
                           n31, Z => n214);
   U1006 : NAN3D1 port map( A1 => n503, A2 => n502, A3 => n504, Z => N1990);
   U1007 : OAI21M20D1 port map( A1 => avs_readdata_21_port, A2 => n700, B => 
                           n28, Z => n212);
   U1008 : NAN3D1 port map( A1 => n509, A2 => n508, A3 => n510, Z => N1988);
   U1009 : OAI21M20D1 port map( A1 => avs_readdata_23_port, A2 => n700, B => 
                           n25, Z => n210);
   U1010 : NAN3D1 port map( A1 => n515, A2 => n514, A3 => n516, Z => N1986);
   U1011 : OAI21M20D1 port map( A1 => avs_readdata_25_port, A2 => n700, B => 
                           n22, Z => n208);
   U1012 : NAN3D1 port map( A1 => n521, A2 => n520, A3 => n522, Z => N1984);
   U1013 : OAI21M20D1 port map( A1 => avs_readdata_27_port, A2 => n700, B => 
                           n19, Z => n206);
   U1014 : NAN3D1 port map( A1 => n527, A2 => n526, A3 => n528, Z => N1982);
   U1015 : OAI21M20D1 port map( A1 => avs_readdata_29_port, A2 => n700, B => 
                           n16, Z => n204);
   U1016 : NAN3D1 port map( A1 => n533, A2 => n532, A3 => n534, Z => N1980);
   U1017 : OAI21M20D1 port map( A1 => avs_readdata_31_port, A2 => n700, B => 
                           n10, Z => n202);
   U1018 : OAI21M20D1 port map( A1 => avs_readdata_9_port, A2 => n700, B => n46
                           , Z => n224);
   U1019 : NAN3D1 port map( A1 => n473, A2 => n472, A3 => n474, Z => N2000);
   U1020 : OAI21M20D1 port map( A1 => avs_readdata_11_port, A2 => n700, B => 
                           n43, Z => n222);
   U1021 : NAN3D1 port map( A1 => n479, A2 => n478, A3 => n480, Z => N1998);
   U1022 : OAI21M20D1 port map( A1 => avs_readdata_13_port, A2 => n700, B => 
                           n40, Z => n220);
   U1023 : NAN3D1 port map( A1 => n485, A2 => n484, A3 => n486, Z => N1996);
   U1024 : AND2D1 port map( A1 => coeff_load, A2 => n104, Z => n301);
   U1025 : MUX2DL port map( A0 => operand_regs_27_port, A1 => coeff_memory_4_27
                           , SL => n712, Z => N3068);
   U1026 : MUX2DL port map( A0 => operand_regs_59_port, A1 => coeff_memory_3_27
                           , SL => n710, Z => N3036);
   U1027 : MUX2DL port map( A0 => operand_regs_123_port, A1 => 
                           coeff_memory_2_27, SL => n718, Z => N3004);
   U1028 : MUX2DL port map( A0 => operand_regs_187_port, A1 => 
                           coeff_memory_1_27, SL => n716, Z => N2972);
   U1029 : MUX2DL port map( A0 => operand_regs_251_port, A1 => 
                           coeff_memory_0_27, SL => n714, Z => N2940);
   U1030 : NAN3D1 port map( A1 => n545, A2 => n544, A3 => n546, Z => N1978);
   U1031 : NAN2D1 port map( A1 => comp_res_31_port, A2 => n554, Z => n545);
   U1032 : AOI22M10D1 port map( B1 => in_buf_63_port, B2 => n540, A1 => n553, 
                           A2 => in_buf_127_port, Z => n442);
   U1033 : NAN3D1 port map( A1 => n446, A2 => n445, A3 => n447, Z => N2009);
   U1034 : NAN2D1 port map( A1 => comp_res_0_port, A2 => n554, Z => n446);
   U1035 : MUX2DL port map( A0 => operand_regs_26_port, A1 => 
                           operand_regs_218_port, SL => n720, Z => n302);
   U1036 : NAN2D1 port map( A1 => comp_res_25_port, A2 => n554, Z => n521);
   U1037 : NAN2D1 port map( A1 => comp_res_27_port, A2 => n554, Z => n527);
   U1038 : NAN2D1 port map( A1 => comp_res_29_port, A2 => n554, Z => n533);
   U1039 : NAN2D1 port map( A1 => comp_res_1_port, A2 => n554, Z => n449);
   U1040 : NAN2D1 port map( A1 => comp_res_3_port, A2 => n541, Z => n455);
   U1041 : NAN2D1 port map( A1 => comp_res_5_port, A2 => n541, Z => n461);
   U1042 : NAN2D1 port map( A1 => comp_res_7_port, A2 => n554, Z => n467);
   U1043 : NAN2D1 port map( A1 => comp_res_9_port, A2 => n541, Z => n473);
   U1044 : NAN2D1 port map( A1 => comp_res_11_port, A2 => n554, Z => n479);
   U1045 : NAN2D1 port map( A1 => comp_res_13_port, A2 => n554, Z => n485);
   U1046 : NAN2D1 port map( A1 => comp_res_15_port, A2 => n554, Z => n491);
   U1047 : NAN2D1 port map( A1 => comp_res_17_port, A2 => n554, Z => n497);
   U1048 : NAN2D1 port map( A1 => comp_res_19_port, A2 => n554, Z => n503);
   U1049 : NAN2D1 port map( A1 => comp_res_21_port, A2 => n554, Z => n509);
   U1050 : NAN2D1 port map( A1 => comp_res_23_port, A2 => n554, Z => n515);
   U1051 : NAN2D1 port map( A1 => comp_res_24_port, A2 => n554, Z => n518);
   U1052 : NAN2D1 port map( A1 => comp_res_26_port, A2 => n554, Z => n524);
   U1053 : NAN2D1 port map( A1 => comp_res_28_port, A2 => n554, Z => n530);
   U1054 : NAN2D1 port map( A1 => comp_res_30_port, A2 => n554, Z => n536);
   U1055 : NAN2D1 port map( A1 => comp_res_2_port, A2 => n541, Z => n452);
   U1056 : NAN2D1 port map( A1 => comp_res_4_port, A2 => n541, Z => n458);
   U1057 : NAN2D1 port map( A1 => comp_res_6_port, A2 => n541, Z => n464);
   U1058 : NAN2D1 port map( A1 => comp_res_8_port, A2 => n541, Z => n470);
   U1059 : NAN2D1 port map( A1 => comp_res_10_port, A2 => n541, Z => n476);
   U1060 : NAN2D1 port map( A1 => comp_res_12_port, A2 => n541, Z => n482);
   U1061 : NAN2D1 port map( A1 => comp_res_14_port, A2 => n541, Z => n488);
   U1062 : NAN2D1 port map( A1 => comp_res_16_port, A2 => n541, Z => n494);
   U1063 : NAN2D1 port map( A1 => comp_res_18_port, A2 => n541, Z => n500);
   U1064 : NAN2D1 port map( A1 => comp_res_20_port, A2 => n541, Z => n506);
   U1065 : NAN2D1 port map( A1 => comp_res_22_port, A2 => n541, Z => n512);
   U1066 : INVD1 port map( A => operand_regs_218_port, Z => n735);
   U1067 : MUX2DL port map( A0 => operand_regs_27_port, A1 => 
                           operand_regs_219_port, SL => n719, Z => n303);
   U1068 : MUX2DL port map( A0 => operand_regs_28_port, A1 => coeff_memory_4_28
                           , SL => n712, Z => N3069);
   U1069 : MUX2DL port map( A0 => operand_regs_60_port, A1 => coeff_memory_3_28
                           , SL => n710, Z => N3037);
   U1070 : MUX2DL port map( A0 => operand_regs_124_port, A1 => 
                           coeff_memory_2_28, SL => n717, Z => N3005);
   U1071 : MUX2DL port map( A0 => operand_regs_188_port, A1 => 
                           coeff_memory_1_28, SL => n716, Z => N2973);
   U1072 : MUX2DL port map( A0 => operand_regs_252_port, A1 => 
                           coeff_memory_0_28, SL => n714, Z => N2941);
   U1073 : NOR2D1 port map( A1 => avs_addr(5), A2 => avs_addr(4), Z => n114);
   U1074 : INVD1 port map( A => operand_regs_219_port, Z => n734);
   U1075 : INVD1 port map( A => avs_addr(0), Z => n762);
   U1076 : AND2D1 port map( A1 => avs_addr(2), A2 => n796, Z => n111);
   U1077 : INVD1 port map( A => avs_addr(1), Z => n796);
   U1078 : AND2D1 port map( A1 => n111, A2 => avs_addr(0), Z => n304);
   U1079 : MUX2DL port map( A0 => operand_regs_28_port, A1 => 
                           operand_regs_220_port, SL => n720, Z => n305);
   U1080 : AND3D1 port map( A1 => avs_addr(0), A2 => avs_addr(1), A3 => n547, Z
                           => n306);
   U1081 : AND3D1 port map( A1 => avs_addr(1), A2 => n547, A3 => n762, Z => 
                           n307);
   U1082 : AND3D1 port map( A1 => avs_addr(0), A2 => n796, A3 => n547, Z => 
                           n308);
   U1083 : AND2D1 port map( A1 => avs_addr(2), A2 => avs_addr(1), Z => n309);
   U1084 : MUX2DL port map( A0 => operand_regs_29_port, A1 => coeff_memory_4_29
                           , SL => n712, Z => N3070);
   U1085 : MUX2DL port map( A0 => operand_regs_61_port, A1 => coeff_memory_3_29
                           , SL => n710, Z => N3038);
   U1086 : MUX2DL port map( A0 => operand_regs_125_port, A1 => 
                           coeff_memory_2_29, SL => n718, Z => N3006);
   U1087 : MUX2DL port map( A0 => operand_regs_189_port, A1 => 
                           coeff_memory_1_29, SL => n716, Z => N2974);
   U1088 : MUX2DL port map( A0 => operand_regs_253_port, A1 => 
                           coeff_memory_0_29, SL => n714, Z => N2942);
   U1089 : INVD1 port map( A => operand_regs_220_port, Z => n733);
   U1090 : NOR2D1 port map( A1 => n92, A2 => n799, Z => n240);
   U1091 : NOR2D1 port map( A1 => n95, A2 => n799, Z => n241);
   U1092 : NAN3D1 port map( A1 => avs_write, A2 => n795, A3 => n304, Z => n179)
                           ;
   U1093 : MUX2DL port map( A0 => operand_regs_29_port, A1 => 
                           operand_regs_221_port, SL => n719, Z => n310);
   U1094 : AO31D1 port map( A1 => avs_write, A2 => n795, A3 => n276, B => 
                           stop_sim_port, Z => n157);
   U1095 : MUX2DL port map( A0 => operand_regs_30_port, A1 => coeff_memory_4_30
                           , SL => n712, Z => N3071);
   U1096 : MUX2DL port map( A0 => operand_regs_62_port, A1 => coeff_memory_3_30
                           , SL => n710, Z => N3039);
   U1097 : MUX2DL port map( A0 => operand_regs_126_port, A1 => 
                           coeff_memory_2_30, SL => n717, Z => N3007);
   U1098 : MUX2DL port map( A0 => operand_regs_190_port, A1 => 
                           coeff_memory_1_30, SL => n716, Z => N2975);
   U1099 : MUX2DL port map( A0 => operand_regs_254_port, A1 => 
                           coeff_memory_0_30, SL => n716, Z => N2943);
   U1100 : MUX2DL port map( A0 => operand_regs_30_port, A1 => 
                           operand_regs_222_port, SL => n720, Z => n311);
   U1101 : INVD1 port map( A => operand_regs_223_port, Z => n730);
   U1102 : INVD1 port map( A => operand_regs_221_port, Z => n732);
   U1103 : INVD1 port map( A => operand_regs_222_port, Z => n731);
   U1104 : MUX2DL port map( A0 => operand_regs_31_port, A1 => coeff_memory_4_31
                           , SL => n712, Z => N3072);
   U1105 : MUX2DL port map( A0 => operand_regs_63_port, A1 => coeff_memory_3_31
                           , SL => n710, Z => N3040);
   U1106 : MUX2DL port map( A0 => operand_regs_255_port, A1 => 
                           coeff_memory_0_31, SL => n712, Z => N2944);
   U1107 : MUX2DL port map( A0 => operand_regs_127_port, A1 => 
                           coeff_memory_2_31, SL => n718, Z => N3008);
   U1108 : MUX2DL port map( A0 => operand_regs_191_port, A1 => 
                           coeff_memory_1_31, SL => n716, Z => N2976);
   U1109 : MUX2DL port map( A0 => operand_regs_31_port, A1 => 
                           operand_regs_223_port, SL => n719, Z => n312);
   U1110 : AO22D1 port map( A1 => N2876, A2 => n697, B1 => N2859, B2 => n812, Z
                           => N2894);
   U1111 : AO22D1 port map( A1 => N2875, A2 => n697, B1 => N2858, B2 => n812, Z
                           => N2895);
   U1112 : AO22D1 port map( A1 => N2874, A2 => n697, B1 => N2857, B2 => n812, Z
                           => N2896);
   U1113 : AO22D1 port map( A1 => N2873, A2 => n697, B1 => N2856, B2 => n812, Z
                           => N2897);
   U1114 : AO22D1 port map( A1 => N2872, A2 => n697, B1 => N2855, B2 => n812, Z
                           => N2898);
   U1115 : AO22D1 port map( A1 => N2871, A2 => n697, B1 => N2854, B2 => n812, Z
                           => N2899);
   U1116 : AO22D1 port map( A1 => N2870, A2 => n697, B1 => N2853, B2 => n812, Z
                           => N2900);
   U1117 : AO22D1 port map( A1 => N2869, A2 => n697, B1 => N2852, B2 => n812, Z
                           => N2901);
   U1118 : AO22D1 port map( A1 => N2868, A2 => n697, B1 => N2851, B2 => n812, Z
                           => N2902);
   U1119 : AO22D1 port map( A1 => N2867, A2 => n697, B1 => N2850, B2 => n812, Z
                           => N2903);
   U1120 : AO22D1 port map( A1 => N2881, A2 => n697, B1 => N2864, B2 => n812, Z
                           => N2889);
   U1121 : AO22D1 port map( A1 => N2880, A2 => n697, B1 => N2863, B2 => n812, Z
                           => N2890);
   U1122 : AO22D1 port map( A1 => N2879, A2 => n697, B1 => N2862, B2 => n812, Z
                           => N2891);
   U1123 : AO22D1 port map( A1 => N2878, A2 => n697, B1 => N2861, B2 => n812, Z
                           => N2892);
   U1124 : AO22D1 port map( A1 => N2877, A2 => n697, B1 => N2860, B2 => n812, Z
                           => N2893);
   U1125 : AO22D1 port map( A1 => N2882, A2 => n697, B1 => N2865, B2 => n812, Z
                           => N2888);
   U1126 : INVD1 port map( A => N64, Z => n696);
   U1127 : NOR2D1 port map( A1 => n801, A2 => out_busy, Z => n79);
   U1128 : NAN3D1 port map( A1 => n81, A2 => out_busy, A3 => N62, Z => n4);
   U1129 : INVD1 port map( A => N62, Z => n810);
   U1130 : BUFD1 port map( A => odd1, Z => n697);
   U1131 : INVD1 port map( A => out_busy, Z => n811);
   U1132 : INVD1 port map( A => odd, Z => n803);
   U1133 : NAN3D1 port map( A1 => in_counter_1_port, A2 => in_busy, A3 => 
                           in_counter_0_port, Z => n88);
   U1134 : NOR2D1 port map( A1 => n806, A2 => in_counter_0_port, Z => n155);
   U1135 : OAI21M20D1 port map( A1 => n806, A2 => in_trigger, B => n100, Z => 
                           n84);
   U1136 : INVD1 port map( A => in_busy, Z => n806);
   U1137 : INVD1 port map( A => in_counter_2_port, Z => n809);
   U1138 : INVD1 port map( A => N63, Z => n813);
   U1139 : NOR2D1 port map( A1 => n804, A2 => in_counter_1_port, Z => n119);
   U1140 : NAN2D1 port map( A1 => in_counter_1_port, A2 => n155, Z => n85);
   U1141 : AND3D1 port map( A1 => in_counter_0_port, A2 => in_busy, A3 => n808,
                           Z => n87);
   U1142 : INVD1 port map( A => in_counter_1_port, Z => n808);
   U1143 : NAN2D1 port map( A1 => n78, A2 => n697, Z => n77);
   U1144 : NOR2D1 port map( A1 => n803, A2 => in_counter_2_port, Z => n101);
   U1145 : NOR2D1 port map( A1 => n809, A2 => odd, Z => n115);
   U1146 : NOR2D1 port map( A1 => odd, A2 => in_counter_2_port, Z => n120);
   U1147 : INVD1 port map( A => out_trigger, Z => n802);
   U1148 : NOR2D1 port map( A1 => n547, A2 => avs_addr(1), Z => n313);
   U1149 : NOR2D1 port map( A1 => n547, A2 => n796, Z => n314);
   U1150 : AOI22D1 port map( A1 => in_buf_64_port, A2 => n243, B1 => 
                           in_buf_0_port, B2 => n262, Z => n320);
   U1151 : NOR2D1 port map( A1 => avs_addr(1), A2 => avs_addr(2), Z => n315);
   U1152 : AND2D1 port map( A1 => n315, A2 => avs_addr(0), Z => n539);
   U1153 : NOR2D1 port map( A1 => n796, A2 => avs_addr(2), Z => n316);
   U1154 : AND2D1 port map( A1 => n316, A2 => avs_addr(0), Z => n538);
   U1155 : AOI22D1 port map( A1 => in_buf_192_port, A2 => n552, B1 => 
                           in_buf_128_port, B2 => n550, Z => n319);
   U1156 : NOR2M1D1 port map( A1 => n313, A2 => avs_addr(0), Z => n541);
   U1157 : NOR2M1D1 port map( A1 => n314, A2 => avs_addr(0), Z => n540);
   U1158 : AOI22D1 port map( A1 => in_buf_96_port, A2 => n554, B1 => 
                           in_buf_32_port, B2 => n540, Z => n318);
   U1159 : NOR2M1D1 port map( A1 => n315, A2 => avs_addr(0), Z => n543);
   U1160 : NOR2M1D1 port map( A1 => n316, A2 => avs_addr(0), Z => n542);
   U1161 : AOI22D1 port map( A1 => in_buf_224_port, A2 => n559, B1 => 
                           in_buf_160_port, B2 => n557, Z => n317);
   U1162 : NAN4D1 port map( A1 => n320, A2 => n319, A3 => n318, A4 => n317, Z 
                           => N2041);
   U1163 : AOI22D1 port map( A1 => in_buf_65_port, A2 => n243, B1 => 
                           in_buf_1_port, B2 => n262, Z => n324);
   U1164 : AOI22D1 port map( A1 => in_buf_193_port, A2 => n539, B1 => 
                           in_buf_129_port, B2 => n538, Z => n323);
   U1165 : AOI22D1 port map( A1 => in_buf_97_port, A2 => n554, B1 => 
                           in_buf_33_port, B2 => n540, Z => n322);
   U1166 : AOI22D1 port map( A1 => in_buf_225_port, A2 => n543, B1 => 
                           in_buf_161_port, B2 => n542, Z => n321);
   U1167 : NAN4D1 port map( A1 => n324, A2 => n323, A3 => n322, A4 => n321, Z 
                           => N2040);
   U1168 : AOI22D1 port map( A1 => in_buf_66_port, A2 => n243, B1 => 
                           in_buf_2_port, B2 => n262, Z => n328);
   U1169 : AOI22D1 port map( A1 => in_buf_194_port, A2 => n539, B1 => 
                           in_buf_130_port, B2 => n538, Z => n327);
   U1170 : AOI22D1 port map( A1 => in_buf_98_port, A2 => n554, B1 => 
                           in_buf_34_port, B2 => n540, Z => n326);
   U1171 : AOI22D1 port map( A1 => in_buf_226_port, A2 => n543, B1 => 
                           in_buf_162_port, B2 => n542, Z => n325);
   U1172 : NAN4D1 port map( A1 => n328, A2 => n327, A3 => n326, A4 => n325, Z 
                           => N2039);
   U1173 : AOI22D1 port map( A1 => in_buf_67_port, A2 => n243, B1 => 
                           in_buf_3_port, B2 => n262, Z => n332);
   U1174 : AOI22D1 port map( A1 => in_buf_195_port, A2 => n539, B1 => 
                           in_buf_131_port, B2 => n538, Z => n331);
   U1175 : AOI22D1 port map( A1 => in_buf_99_port, A2 => n554, B1 => 
                           in_buf_35_port, B2 => n540, Z => n330);
   U1176 : AOI22D1 port map( A1 => in_buf_227_port, A2 => n543, B1 => 
                           in_buf_163_port, B2 => n542, Z => n329);
   U1177 : NAN4D1 port map( A1 => n332, A2 => n331, A3 => n330, A4 => n329, Z 
                           => N2038);
   U1178 : AOI22D1 port map( A1 => in_buf_68_port, A2 => n243, B1 => 
                           in_buf_4_port, B2 => n262, Z => n336);
   U1179 : AOI22D1 port map( A1 => in_buf_196_port, A2 => n539, B1 => 
                           in_buf_132_port, B2 => n538, Z => n335);
   U1180 : AOI22D1 port map( A1 => in_buf_100_port, A2 => n554, B1 => 
                           in_buf_36_port, B2 => n540, Z => n334);
   U1181 : AOI22D1 port map( A1 => in_buf_228_port, A2 => n543, B1 => 
                           in_buf_164_port, B2 => n542, Z => n333);
   U1182 : NAN4D1 port map( A1 => n336, A2 => n335, A3 => n334, A4 => n333, Z 
                           => N2037);
   U1183 : AOI22D1 port map( A1 => in_buf_69_port, A2 => n243, B1 => 
                           in_buf_5_port, B2 => n262, Z => n340);
   U1184 : AOI22D1 port map( A1 => in_buf_197_port, A2 => n539, B1 => 
                           in_buf_133_port, B2 => n538, Z => n339);
   U1185 : AOI22D1 port map( A1 => in_buf_101_port, A2 => n554, B1 => 
                           in_buf_37_port, B2 => n540, Z => n338);
   U1186 : AOI22D1 port map( A1 => in_buf_229_port, A2 => n543, B1 => 
                           in_buf_165_port, B2 => n542, Z => n337);
   U1187 : NAN4D1 port map( A1 => n340, A2 => n339, A3 => n338, A4 => n337, Z 
                           => N2036);
   U1188 : AOI22D1 port map( A1 => in_buf_70_port, A2 => n243, B1 => 
                           in_buf_6_port, B2 => n262, Z => n344);
   U1189 : AOI22D1 port map( A1 => in_buf_198_port, A2 => n539, B1 => 
                           in_buf_134_port, B2 => n538, Z => n343);
   U1190 : AOI22D1 port map( A1 => in_buf_102_port, A2 => n554, B1 => 
                           in_buf_38_port, B2 => n540, Z => n342);
   U1191 : AOI22D1 port map( A1 => in_buf_230_port, A2 => n543, B1 => 
                           in_buf_166_port, B2 => n542, Z => n341);
   U1192 : NAN4D1 port map( A1 => n344, A2 => n343, A3 => n342, A4 => n341, Z 
                           => N2035);
   U1193 : AOI22D1 port map( A1 => in_buf_71_port, A2 => n243, B1 => 
                           in_buf_7_port, B2 => n262, Z => n348);
   U1194 : AOI22D1 port map( A1 => in_buf_199_port, A2 => n539, B1 => 
                           in_buf_135_port, B2 => n538, Z => n347);
   U1195 : AOI22D1 port map( A1 => in_buf_103_port, A2 => n554, B1 => 
                           in_buf_39_port, B2 => n540, Z => n346);
   U1196 : AOI22D1 port map( A1 => in_buf_231_port, A2 => n543, B1 => 
                           in_buf_167_port, B2 => n542, Z => n345);
   U1197 : NAN4D1 port map( A1 => n348, A2 => n347, A3 => n346, A4 => n345, Z 
                           => N2034);
   U1198 : AOI22D1 port map( A1 => in_buf_72_port, A2 => n243, B1 => 
                           in_buf_8_port, B2 => n262, Z => n352);
   U1199 : AOI22D1 port map( A1 => in_buf_200_port, A2 => n539, B1 => 
                           in_buf_136_port, B2 => n538, Z => n351);
   U1200 : AOI22D1 port map( A1 => in_buf_104_port, A2 => n541, B1 => 
                           in_buf_40_port, B2 => n540, Z => n350);
   U1201 : AOI22D1 port map( A1 => in_buf_232_port, A2 => n543, B1 => 
                           in_buf_168_port, B2 => n542, Z => n349);
   U1202 : NAN4D1 port map( A1 => n352, A2 => n351, A3 => n350, A4 => n349, Z 
                           => N2033);
   U1203 : AOI22D1 port map( A1 => in_buf_73_port, A2 => n243, B1 => 
                           in_buf_9_port, B2 => n262, Z => n356);
   U1204 : AOI22D1 port map( A1 => in_buf_201_port, A2 => n539, B1 => 
                           in_buf_137_port, B2 => n538, Z => n355);
   U1205 : AOI22D1 port map( A1 => in_buf_105_port, A2 => n541, B1 => 
                           in_buf_41_port, B2 => n540, Z => n354);
   U1206 : AOI22D1 port map( A1 => in_buf_233_port, A2 => n543, B1 => 
                           in_buf_169_port, B2 => n542, Z => n353);
   U1207 : NAN4D1 port map( A1 => n356, A2 => n355, A3 => n354, A4 => n353, Z 
                           => N2032);
   U1208 : AOI22D1 port map( A1 => in_buf_74_port, A2 => n243, B1 => 
                           in_buf_10_port, B2 => n262, Z => n360);
   U1209 : AOI22D1 port map( A1 => in_buf_202_port, A2 => n539, B1 => 
                           in_buf_138_port, B2 => n538, Z => n359);
   U1210 : AOI22D1 port map( A1 => in_buf_106_port, A2 => n541, B1 => 
                           in_buf_42_port, B2 => n540, Z => n358);
   U1211 : AOI22D1 port map( A1 => in_buf_234_port, A2 => n559, B1 => 
                           in_buf_170_port, B2 => n542, Z => n357);
   U1212 : NAN4D1 port map( A1 => n360, A2 => n359, A3 => n358, A4 => n357, Z 
                           => N2031);
   U1213 : AOI22D1 port map( A1 => in_buf_75_port, A2 => n243, B1 => 
                           in_buf_11_port, B2 => n262, Z => n364);
   U1214 : AOI22D1 port map( A1 => in_buf_203_port, A2 => n539, B1 => 
                           in_buf_139_port, B2 => n538, Z => n363);
   U1215 : AOI22D1 port map( A1 => in_buf_107_port, A2 => n541, B1 => 
                           in_buf_43_port, B2 => n540, Z => n362);
   U1216 : AOI22D1 port map( A1 => in_buf_235_port, A2 => n543, B1 => 
                           in_buf_171_port, B2 => n542, Z => n361);
   U1217 : NAN4D1 port map( A1 => n364, A2 => n363, A3 => n362, A4 => n361, Z 
                           => N2030);
   U1218 : AOI22D1 port map( A1 => in_buf_76_port, A2 => n243, B1 => 
                           in_buf_12_port, B2 => n262, Z => n368);
   U1219 : AOI22D1 port map( A1 => in_buf_204_port, A2 => n539, B1 => 
                           in_buf_140_port, B2 => n538, Z => n367);
   U1220 : AOI22D1 port map( A1 => in_buf_108_port, A2 => n554, B1 => 
                           in_buf_44_port, B2 => n540, Z => n366);
   U1221 : AOI22D1 port map( A1 => in_buf_236_port, A2 => n559, B1 => 
                           in_buf_172_port, B2 => n557, Z => n365);
   U1222 : NAN4D1 port map( A1 => n368, A2 => n367, A3 => n366, A4 => n365, Z 
                           => N2029);
   U1223 : AOI22D1 port map( A1 => in_buf_77_port, A2 => n243, B1 => 
                           in_buf_13_port, B2 => n262, Z => n372);
   U1224 : AOI22D1 port map( A1 => in_buf_205_port, A2 => n552, B1 => 
                           in_buf_141_port, B2 => n550, Z => n371);
   U1225 : AOI22D1 port map( A1 => in_buf_109_port, A2 => n541, B1 => 
                           in_buf_45_port, B2 => n540, Z => n370);
   U1226 : AOI22D1 port map( A1 => in_buf_237_port, A2 => n559, B1 => 
                           in_buf_173_port, B2 => n556, Z => n369);
   U1227 : NAN4D1 port map( A1 => n372, A2 => n371, A3 => n370, A4 => n369, Z 
                           => N2028);
   U1228 : AOI22D1 port map( A1 => in_buf_78_port, A2 => n243, B1 => 
                           in_buf_14_port, B2 => n262, Z => n376);
   U1229 : AOI22D1 port map( A1 => in_buf_206_port, A2 => n552, B1 => 
                           in_buf_142_port, B2 => n550, Z => n375);
   U1230 : AOI22D1 port map( A1 => in_buf_110_port, A2 => n541, B1 => 
                           in_buf_46_port, B2 => n540, Z => n374);
   U1231 : AOI22D1 port map( A1 => in_buf_238_port, A2 => n559, B1 => 
                           in_buf_174_port, B2 => n542, Z => n373);
   U1232 : NAN4D1 port map( A1 => n376, A2 => n375, A3 => n374, A4 => n373, Z 
                           => N2027);
   U1233 : AOI22D1 port map( A1 => in_buf_79_port, A2 => n243, B1 => 
                           in_buf_15_port, B2 => n262, Z => n380);
   U1234 : AOI22D1 port map( A1 => in_buf_207_port, A2 => n552, B1 => 
                           in_buf_143_port, B2 => n550, Z => n379);
   U1235 : AOI22D1 port map( A1 => in_buf_111_port, A2 => n541, B1 => 
                           in_buf_47_port, B2 => n540, Z => n378);
   U1236 : AOI22D1 port map( A1 => in_buf_239_port, A2 => n559, B1 => 
                           in_buf_175_port, B2 => n542, Z => n377);
   U1237 : NAN4D1 port map( A1 => n380, A2 => n379, A3 => n378, A4 => n377, Z 
                           => N2026);
   U1238 : AOI22D1 port map( A1 => in_buf_80_port, A2 => n243, B1 => 
                           in_buf_16_port, B2 => n262, Z => n384);
   U1239 : AOI22D1 port map( A1 => in_buf_208_port, A2 => n552, B1 => 
                           in_buf_144_port, B2 => n550, Z => n383);
   U1240 : AOI22D1 port map( A1 => in_buf_112_port, A2 => n541, B1 => 
                           in_buf_48_port, B2 => n540, Z => n382);
   U1241 : AOI22D1 port map( A1 => in_buf_240_port, A2 => n559, B1 => 
                           in_buf_176_port, B2 => n542, Z => n381);
   U1242 : NAN4D1 port map( A1 => n384, A2 => n383, A3 => n382, A4 => n381, Z 
                           => N2025);
   U1243 : AOI22D1 port map( A1 => in_buf_81_port, A2 => n243, B1 => 
                           in_buf_17_port, B2 => n262, Z => n388);
   U1244 : AOI22D1 port map( A1 => in_buf_209_port, A2 => n552, B1 => 
                           in_buf_145_port, B2 => n550, Z => n387);
   U1245 : AOI22D1 port map( A1 => in_buf_113_port, A2 => n541, B1 => 
                           in_buf_49_port, B2 => n540, Z => n386);
   U1246 : AOI22D1 port map( A1 => in_buf_241_port, A2 => n559, B1 => 
                           in_buf_177_port, B2 => n542, Z => n385);
   U1247 : NAN4D1 port map( A1 => n388, A2 => n387, A3 => n386, A4 => n385, Z 
                           => N2024);
   U1248 : AOI22D1 port map( A1 => in_buf_82_port, A2 => n243, B1 => 
                           in_buf_18_port, B2 => n262, Z => n392);
   U1249 : AOI22D1 port map( A1 => in_buf_210_port, A2 => n552, B1 => 
                           in_buf_146_port, B2 => n550, Z => n391);
   U1250 : AOI22D1 port map( A1 => in_buf_114_port, A2 => n541, B1 => 
                           in_buf_50_port, B2 => n540, Z => n390);
   U1251 : AOI22D1 port map( A1 => in_buf_242_port, A2 => n559, B1 => 
                           in_buf_178_port, B2 => n542, Z => n389);
   U1252 : NAN4D1 port map( A1 => n392, A2 => n391, A3 => n390, A4 => n389, Z 
                           => N2023);
   U1253 : AOI22D1 port map( A1 => in_buf_83_port, A2 => n243, B1 => 
                           in_buf_19_port, B2 => n262, Z => n396);
   U1254 : AOI22D1 port map( A1 => in_buf_211_port, A2 => n552, B1 => 
                           in_buf_147_port, B2 => n550, Z => n395);
   U1255 : AOI22D1 port map( A1 => in_buf_115_port, A2 => n541, B1 => 
                           in_buf_51_port, B2 => n540, Z => n394);
   U1256 : AOI22D1 port map( A1 => in_buf_243_port, A2 => n559, B1 => 
                           in_buf_179_port, B2 => n542, Z => n393);
   U1257 : NAN4D1 port map( A1 => n396, A2 => n395, A3 => n394, A4 => n393, Z 
                           => N2022);
   U1258 : AOI22D1 port map( A1 => in_buf_84_port, A2 => n243, B1 => 
                           in_buf_20_port, B2 => n262, Z => n400);
   U1259 : AOI22D1 port map( A1 => in_buf_212_port, A2 => n552, B1 => 
                           in_buf_148_port, B2 => n550, Z => n399);
   U1260 : AOI22D1 port map( A1 => in_buf_116_port, A2 => n541, B1 => 
                           in_buf_52_port, B2 => n540, Z => n398);
   U1261 : AOI22D1 port map( A1 => in_buf_244_port, A2 => n559, B1 => 
                           in_buf_180_port, B2 => n542, Z => n397);
   U1262 : NAN4D1 port map( A1 => n400, A2 => n399, A3 => n398, A4 => n397, Z 
                           => N2021);
   U1263 : AOI22D1 port map( A1 => in_buf_85_port, A2 => n243, B1 => 
                           in_buf_21_port, B2 => n262, Z => n404);
   U1264 : AOI22D1 port map( A1 => in_buf_213_port, A2 => n552, B1 => 
                           in_buf_149_port, B2 => n550, Z => n403);
   U1265 : AOI22D1 port map( A1 => in_buf_117_port, A2 => n541, B1 => 
                           in_buf_53_port, B2 => n540, Z => n402);
   U1266 : AOI22D1 port map( A1 => in_buf_245_port, A2 => n559, B1 => 
                           in_buf_181_port, B2 => n542, Z => n401);
   U1267 : NAN4D1 port map( A1 => n404, A2 => n403, A3 => n402, A4 => n401, Z 
                           => N2020);
   U1268 : AOI22D1 port map( A1 => in_buf_86_port, A2 => n243, B1 => 
                           in_buf_22_port, B2 => n262, Z => n408);
   U1269 : AOI22D1 port map( A1 => in_buf_214_port, A2 => n552, B1 => 
                           in_buf_150_port, B2 => n550, Z => n407);
   U1270 : AOI22D1 port map( A1 => in_buf_118_port, A2 => n541, B1 => 
                           in_buf_54_port, B2 => n540, Z => n406);
   U1271 : AOI22D1 port map( A1 => in_buf_246_port, A2 => n559, B1 => 
                           in_buf_182_port, B2 => n542, Z => n405);
   U1272 : NAN4D1 port map( A1 => n408, A2 => n407, A3 => n406, A4 => n405, Z 
                           => N2019);
   U1273 : AOI22D1 port map( A1 => in_buf_87_port, A2 => n243, B1 => 
                           in_buf_23_port, B2 => n262, Z => n412);
   U1274 : AOI22D1 port map( A1 => in_buf_215_port, A2 => n552, B1 => 
                           in_buf_151_port, B2 => n550, Z => n411);
   U1275 : AOI22D1 port map( A1 => in_buf_119_port, A2 => n541, B1 => 
                           in_buf_55_port, B2 => n540, Z => n410);
   U1276 : AOI22D1 port map( A1 => in_buf_247_port, A2 => n559, B1 => 
                           in_buf_183_port, B2 => n542, Z => n409);
   U1277 : NAN4D1 port map( A1 => n412, A2 => n411, A3 => n410, A4 => n409, Z 
                           => N2018);
   U1278 : AOI22D1 port map( A1 => in_buf_88_port, A2 => n243, B1 => 
                           in_buf_24_port, B2 => n262, Z => n416);
   U1279 : AOI22D1 port map( A1 => in_buf_216_port, A2 => n552, B1 => 
                           in_buf_152_port, B2 => n550, Z => n415);
   U1280 : AOI22D1 port map( A1 => in_buf_120_port, A2 => n541, B1 => 
                           in_buf_56_port, B2 => n540, Z => n414);
   U1281 : AOI22D1 port map( A1 => in_buf_248_port, A2 => n559, B1 => 
                           in_buf_184_port, B2 => n542, Z => n413);
   U1282 : NAN4D1 port map( A1 => n416, A2 => n415, A3 => n414, A4 => n413, Z 
                           => N2017);
   U1283 : AOI22D1 port map( A1 => in_buf_89_port, A2 => n243, B1 => 
                           in_buf_25_port, B2 => n262, Z => n420);
   U1284 : AOI22D1 port map( A1 => in_buf_217_port, A2 => n552, B1 => 
                           in_buf_153_port, B2 => n550, Z => n419);
   U1285 : AOI22D1 port map( A1 => in_buf_121_port, A2 => n541, B1 => 
                           in_buf_57_port, B2 => n540, Z => n418);
   U1286 : AOI22D1 port map( A1 => in_buf_249_port, A2 => n559, B1 => 
                           in_buf_185_port, B2 => n556, Z => n417);
   U1287 : NAN4D1 port map( A1 => n420, A2 => n419, A3 => n418, A4 => n417, Z 
                           => N2016);
   U1288 : AOI22D1 port map( A1 => in_buf_90_port, A2 => n243, B1 => 
                           in_buf_26_port, B2 => n262, Z => n424);
   U1289 : AOI22D1 port map( A1 => in_buf_218_port, A2 => n552, B1 => 
                           in_buf_154_port, B2 => n549, Z => n423);
   U1290 : AOI22D1 port map( A1 => in_buf_122_port, A2 => n541, B1 => 
                           in_buf_58_port, B2 => n540, Z => n422);
   U1291 : AOI22D1 port map( A1 => in_buf_250_port, A2 => n543, B1 => 
                           in_buf_186_port, B2 => n557, Z => n421);
   U1292 : NAN4D1 port map( A1 => n424, A2 => n423, A3 => n422, A4 => n421, Z 
                           => N2015);
   U1293 : AOI22D1 port map( A1 => in_buf_91_port, A2 => n243, B1 => 
                           in_buf_27_port, B2 => n262, Z => n428);
   U1294 : AOI22D1 port map( A1 => in_buf_219_port, A2 => n539, B1 => 
                           in_buf_155_port, B2 => n549, Z => n427);
   U1295 : AOI22D1 port map( A1 => in_buf_123_port, A2 => n541, B1 => 
                           in_buf_59_port, B2 => n540, Z => n426);
   U1296 : AOI22D1 port map( A1 => in_buf_251_port, A2 => n543, B1 => 
                           in_buf_187_port, B2 => n557, Z => n425);
   U1297 : NAN4D1 port map( A1 => n428, A2 => n427, A3 => n426, A4 => n425, Z 
                           => N2014);
   U1298 : AOI22D1 port map( A1 => in_buf_92_port, A2 => n243, B1 => 
                           in_buf_28_port, B2 => n262, Z => n432);
   U1299 : AOI22D1 port map( A1 => in_buf_220_port, A2 => n539, B1 => 
                           in_buf_156_port, B2 => n549, Z => n431);
   U1300 : AOI22D1 port map( A1 => in_buf_124_port, A2 => n541, B1 => 
                           in_buf_60_port, B2 => n540, Z => n430);
   U1301 : AOI22D1 port map( A1 => in_buf_252_port, A2 => n543, B1 => 
                           in_buf_188_port, B2 => n557, Z => n429);
   U1302 : NAN4D1 port map( A1 => n432, A2 => n431, A3 => n430, A4 => n429, Z 
                           => N2013);
   U1303 : AOI22D1 port map( A1 => in_buf_93_port, A2 => n243, B1 => 
                           in_buf_29_port, B2 => n262, Z => n436);
   U1304 : AOI22D1 port map( A1 => in_buf_221_port, A2 => n539, B1 => 
                           in_buf_157_port, B2 => n549, Z => n435);
   U1305 : AOI22D1 port map( A1 => in_buf_125_port, A2 => n541, B1 => 
                           in_buf_61_port, B2 => n540, Z => n434);
   U1306 : AOI22D1 port map( A1 => in_buf_253_port, A2 => n543, B1 => 
                           in_buf_189_port, B2 => n557, Z => n433);
   U1307 : NAN4D1 port map( A1 => n436, A2 => n435, A3 => n434, A4 => n433, Z 
                           => N2012);
   U1308 : AOI22D1 port map( A1 => in_buf_94_port, A2 => n243, B1 => 
                           in_buf_30_port, B2 => n262, Z => n440);
   U1309 : AOI22D1 port map( A1 => in_buf_222_port, A2 => n552, B1 => 
                           in_buf_158_port, B2 => n549, Z => n439);
   U1310 : AOI22D1 port map( A1 => in_buf_126_port, A2 => n541, B1 => 
                           in_buf_62_port, B2 => n540, Z => n438);
   U1311 : AOI22D1 port map( A1 => in_buf_254_port, A2 => n559, B1 => 
                           in_buf_190_port, B2 => n557, Z => n437);
   U1312 : NAN4D1 port map( A1 => n440, A2 => n439, A3 => n438, A4 => n437, Z 
                           => N2011);
   U1313 : AOI22D1 port map( A1 => in_buf_95_port, A2 => n243, B1 => 
                           in_buf_31_port, B2 => n262, Z => n444);
   U1314 : AOI22D1 port map( A1 => in_buf_223_port, A2 => n539, B1 => 
                           in_buf_159_port, B2 => n549, Z => n443);
   U1315 : AOI22D1 port map( A1 => in_buf_255_port, A2 => n543, B1 => 
                           in_buf_191_port, B2 => n557, Z => n441);
   U1316 : NAN4D1 port map( A1 => n444, A2 => n443, A3 => n442, A4 => n441, Z 
                           => N2010);
   U1317 : AOI22D1 port map( A1 => comp_res_96_port, A2 => n539, B1 => 
                           comp_res_32_port, B2 => n549, Z => n447);
   U1318 : AOI22D1 port map( A1 => comp_res_128_port, A2 => n543, B1 => 
                           comp_res_64_port, B2 => n557, Z => n445);
   U1319 : AOI22D1 port map( A1 => comp_res_97_port, A2 => n539, B1 => 
                           comp_res_33_port, B2 => n549, Z => n450);
   U1320 : AOI22D1 port map( A1 => comp_res_129_port, A2 => n543, B1 => 
                           comp_res_65_port, B2 => n557, Z => n448);
   U1321 : AOI22D1 port map( A1 => comp_res_98_port, A2 => n539, B1 => 
                           comp_res_34_port, B2 => n549, Z => n453);
   U1322 : AOI22D1 port map( A1 => comp_res_130_port, A2 => n543, B1 => 
                           comp_res_66_port, B2 => n557, Z => n451);
   U1323 : AOI22D1 port map( A1 => comp_res_99_port, A2 => n539, B1 => 
                           comp_res_35_port, B2 => n549, Z => n456);
   U1324 : AOI22D1 port map( A1 => comp_res_131_port, A2 => n543, B1 => 
                           comp_res_67_port, B2 => n557, Z => n454);
   U1325 : AOI22D1 port map( A1 => comp_res_100_port, A2 => n539, B1 => 
                           comp_res_36_port, B2 => n549, Z => n459);
   U1326 : AOI22D1 port map( A1 => comp_res_132_port, A2 => n543, B1 => 
                           comp_res_68_port, B2 => n557, Z => n457);
   U1327 : AOI22D1 port map( A1 => comp_res_101_port, A2 => n539, B1 => 
                           comp_res_37_port, B2 => n549, Z => n462);
   U1328 : AOI22D1 port map( A1 => comp_res_133_port, A2 => n543, B1 => 
                           comp_res_69_port, B2 => n557, Z => n460);
   U1329 : AOI22D1 port map( A1 => comp_res_102_port, A2 => n539, B1 => 
                           comp_res_38_port, B2 => n549, Z => n465);
   U1330 : AOI22D1 port map( A1 => comp_res_134_port, A2 => n543, B1 => 
                           comp_res_70_port, B2 => n557, Z => n463);
   U1331 : AOI22D1 port map( A1 => comp_res_103_port, A2 => n539, B1 => 
                           comp_res_39_port, B2 => n550, Z => n468);
   U1332 : AOI22D1 port map( A1 => comp_res_135_port, A2 => n543, B1 => 
                           comp_res_71_port, B2 => n556, Z => n466);
   U1333 : AOI22D1 port map( A1 => comp_res_104_port, A2 => n539, B1 => 
                           comp_res_40_port, B2 => n538, Z => n471);
   U1334 : AOI22D1 port map( A1 => comp_res_136_port, A2 => n559, B1 => 
                           comp_res_72_port, B2 => n542, Z => n469);
   U1335 : AOI22D1 port map( A1 => comp_res_105_port, A2 => n539, B1 => 
                           comp_res_41_port, B2 => n550, Z => n474);
   U1336 : AOI22D1 port map( A1 => comp_res_137_port, A2 => n543, B1 => 
                           comp_res_73_port, B2 => n542, Z => n472);
   U1337 : AOI22D1 port map( A1 => comp_res_106_port, A2 => n539, B1 => 
                           comp_res_42_port, B2 => n549, Z => n477);
   U1338 : AOI22D1 port map( A1 => comp_res_138_port, A2 => n559, B1 => 
                           comp_res_74_port, B2 => n542, Z => n475);
   U1339 : AOI22D1 port map( A1 => comp_res_107_port, A2 => n552, B1 => 
                           comp_res_43_port, B2 => n538, Z => n480);
   U1340 : AOI22D1 port map( A1 => comp_res_139_port, A2 => n543, B1 => 
                           comp_res_75_port, B2 => n557, Z => n478);
   U1341 : AOI22D1 port map( A1 => comp_res_108_port, A2 => n539, B1 => 
                           comp_res_44_port, B2 => n550, Z => n483);
   U1342 : AOI22D1 port map( A1 => comp_res_140_port, A2 => n559, B1 => 
                           comp_res_76_port, B2 => n542, Z => n481);
   U1343 : AOI22D1 port map( A1 => comp_res_109_port, A2 => n539, B1 => 
                           comp_res_45_port, B2 => n549, Z => n486);
   U1344 : AOI22D1 port map( A1 => comp_res_141_port, A2 => n543, B1 => 
                           comp_res_77_port, B2 => n542, Z => n484);
   U1345 : AOI22D1 port map( A1 => comp_res_110_port, A2 => n539, B1 => 
                           comp_res_46_port, B2 => n538, Z => n489);
   U1346 : AOI22D1 port map( A1 => comp_res_142_port, A2 => n559, B1 => 
                           comp_res_78_port, B2 => n557, Z => n487);
   U1347 : AOI22D1 port map( A1 => comp_res_111_port, A2 => n539, B1 => 
                           comp_res_47_port, B2 => n549, Z => n492);
   U1348 : AOI22D1 port map( A1 => comp_res_143_port, A2 => n543, B1 => 
                           comp_res_79_port, B2 => n556, Z => n490);
   U1349 : AOI22D1 port map( A1 => comp_res_112_port, A2 => n539, B1 => 
                           comp_res_48_port, B2 => n538, Z => n495);
   U1350 : AOI22D1 port map( A1 => comp_res_144_port, A2 => n543, B1 => 
                           comp_res_80_port, B2 => n542, Z => n493);
   U1351 : AOI22D1 port map( A1 => comp_res_113_port, A2 => n539, B1 => 
                           comp_res_49_port, B2 => n538, Z => n498);
   U1352 : AOI22D1 port map( A1 => comp_res_145_port, A2 => n543, B1 => 
                           comp_res_81_port, B2 => n556, Z => n496);
   U1353 : AOI22D1 port map( A1 => comp_res_114_port, A2 => n539, B1 => 
                           comp_res_50_port, B2 => n549, Z => n501);
   U1354 : AOI22D1 port map( A1 => comp_res_146_port, A2 => n559, B1 => 
                           comp_res_82_port, B2 => n556, Z => n499);
   U1355 : AOI22D1 port map( A1 => comp_res_115_port, A2 => n539, B1 => 
                           comp_res_51_port, B2 => n549, Z => n504);
   U1356 : AOI22D1 port map( A1 => comp_res_147_port, A2 => n543, B1 => 
                           comp_res_83_port, B2 => n556, Z => n502);
   U1357 : AOI22D1 port map( A1 => comp_res_116_port, A2 => n539, B1 => 
                           comp_res_52_port, B2 => n538, Z => n507);
   U1358 : AOI22D1 port map( A1 => comp_res_148_port, A2 => n543, B1 => 
                           comp_res_84_port, B2 => n556, Z => n505);
   U1359 : AOI22D1 port map( A1 => comp_res_117_port, A2 => n539, B1 => 
                           comp_res_53_port, B2 => n538, Z => n510);
   U1360 : AOI22D1 port map( A1 => comp_res_149_port, A2 => n543, B1 => 
                           comp_res_85_port, B2 => n556, Z => n508);
   U1361 : AOI22D1 port map( A1 => comp_res_118_port, A2 => n539, B1 => 
                           comp_res_54_port, B2 => n538, Z => n513);
   U1362 : AOI22D1 port map( A1 => comp_res_150_port, A2 => n543, B1 => 
                           comp_res_86_port, B2 => n556, Z => n511);
   U1363 : AOI22D1 port map( A1 => comp_res_119_port, A2 => n539, B1 => 
                           comp_res_55_port, B2 => n538, Z => n516);
   U1364 : AOI22D1 port map( A1 => comp_res_151_port, A2 => n543, B1 => 
                           comp_res_87_port, B2 => n556, Z => n514);
   U1365 : AOI22D1 port map( A1 => comp_res_120_port, A2 => n539, B1 => 
                           comp_res_56_port, B2 => n538, Z => n519);
   U1366 : AOI22D1 port map( A1 => comp_res_152_port, A2 => n543, B1 => 
                           comp_res_88_port, B2 => n556, Z => n517);
   U1367 : AOI22D1 port map( A1 => comp_res_121_port, A2 => n539, B1 => 
                           comp_res_57_port, B2 => n538, Z => n522);
   U1368 : AOI22D1 port map( A1 => comp_res_153_port, A2 => n559, B1 => 
                           comp_res_89_port, B2 => n556, Z => n520);
   U1369 : AOI22D1 port map( A1 => comp_res_122_port, A2 => n539, B1 => 
                           comp_res_58_port, B2 => n538, Z => n525);
   U1370 : AOI22D1 port map( A1 => comp_res_154_port, A2 => n543, B1 => 
                           comp_res_90_port, B2 => n556, Z => n523);
   U1371 : AOI22D1 port map( A1 => comp_res_123_port, A2 => n552, B1 => 
                           comp_res_59_port, B2 => n538, Z => n528);
   U1372 : AOI22D1 port map( A1 => comp_res_155_port, A2 => n543, B1 => 
                           comp_res_91_port, B2 => n556, Z => n526);
   U1373 : AOI22D1 port map( A1 => comp_res_124_port, A2 => n539, B1 => 
                           comp_res_60_port, B2 => n538, Z => n531);
   U1374 : AOI22D1 port map( A1 => comp_res_156_port, A2 => n559, B1 => 
                           comp_res_92_port, B2 => n556, Z => n529);
   U1375 : AOI22D1 port map( A1 => comp_res_125_port, A2 => n539, B1 => 
                           comp_res_61_port, B2 => n538, Z => n534);
   U1376 : AOI22D1 port map( A1 => comp_res_157_port, A2 => n543, B1 => 
                           comp_res_93_port, B2 => n556, Z => n532);
   U1377 : AOI22D1 port map( A1 => comp_res_126_port, A2 => n539, B1 => 
                           comp_res_62_port, B2 => n538, Z => n537);
   U1378 : AOI22D1 port map( A1 => comp_res_158_port, A2 => n559, B1 => 
                           comp_res_94_port, B2 => n556, Z => n535);
   U1379 : AOI22D1 port map( A1 => comp_res_127_port, A2 => n539, B1 => 
                           comp_res_63_port, B2 => n550, Z => n546);
   U1380 : AOI22D1 port map( A1 => comp_res_159_port, A2 => n543, B1 => 
                           comp_res_95_port, B2 => n556, Z => n544);
   U1381 : NOR2D1 port map( A1 => n696, A2 => N63, Z => n560);
   U1382 : NOR2D1 port map( A1 => n696, A2 => n813, Z => n561);
   U1383 : AOI22D1 port map( A1 => out_buf_80_port, A2 => n269, B1 => 
                           out_buf_16_port, B2 => n244, Z => n567);
   U1384 : NOR2D1 port map( A1 => N63, A2 => N64, Z => n562);
   U1385 : NOR2D1 port map( A1 => n813, A2 => N64, Z => n563);
   U1386 : AOI22D1 port map( A1 => out_buf_208_port, A2 => n270, B1 => 
                           out_buf_144_port, B2 => n245, Z => n566);
   U1387 : NOR2M1D1 port map( A1 => n560, A2 => N62, Z => n689);
   U1388 : NOR2M1D1 port map( A1 => n561, A2 => N62, Z => n688);
   U1389 : AOI22D1 port map( A1 => out_buf_112_port, A2 => n689, B1 => 
                           out_buf_48_port, B2 => n688, Z => n565);
   U1390 : NOR2M1D1 port map( A1 => n562, A2 => N62, Z => n691);
   U1391 : NOR2M1D1 port map( A1 => n563, A2 => N62, Z => n690);
   U1392 : AOI22D1 port map( A1 => out_buf_240_port, A2 => n691, B1 => 
                           out_buf_176_port, B2 => n690, Z => n564);
   U1393 : NAN4D1 port map( A1 => n567, A2 => n566, A3 => n565, A4 => n564, Z 
                           => N2882);
   U1394 : AOI22D1 port map( A1 => out_buf_81_port, A2 => n269, B1 => 
                           out_buf_17_port, B2 => n244, Z => n571);
   U1395 : AOI22D1 port map( A1 => out_buf_209_port, A2 => n270, B1 => 
                           out_buf_145_port, B2 => n245, Z => n570);
   U1396 : AOI22D1 port map( A1 => out_buf_113_port, A2 => n689, B1 => 
                           out_buf_49_port, B2 => n688, Z => n569);
   U1397 : AOI22D1 port map( A1 => out_buf_241_port, A2 => n691, B1 => 
                           out_buf_177_port, B2 => n690, Z => n568);
   U1398 : NAN4D1 port map( A1 => n571, A2 => n570, A3 => n569, A4 => n568, Z 
                           => N2881);
   U1399 : AOI22D1 port map( A1 => out_buf_82_port, A2 => n269, B1 => 
                           out_buf_18_port, B2 => n244, Z => n575);
   U1400 : AOI22D1 port map( A1 => out_buf_210_port, A2 => n270, B1 => 
                           out_buf_146_port, B2 => n245, Z => n574);
   U1401 : AOI22D1 port map( A1 => out_buf_114_port, A2 => n689, B1 => 
                           out_buf_50_port, B2 => n688, Z => n573);
   U1402 : AOI22D1 port map( A1 => out_buf_242_port, A2 => n691, B1 => 
                           out_buf_178_port, B2 => n690, Z => n572);
   U1403 : NAN4D1 port map( A1 => n575, A2 => n574, A3 => n573, A4 => n572, Z 
                           => N2880);
   U1404 : AOI22D1 port map( A1 => out_buf_83_port, A2 => n269, B1 => 
                           out_buf_19_port, B2 => n244, Z => n579);
   U1405 : AOI22D1 port map( A1 => out_buf_211_port, A2 => n270, B1 => 
                           out_buf_147_port, B2 => n245, Z => n578);
   U1406 : AOI22D1 port map( A1 => out_buf_115_port, A2 => n689, B1 => 
                           out_buf_51_port, B2 => n688, Z => n577);
   U1407 : AOI22D1 port map( A1 => out_buf_243_port, A2 => n691, B1 => 
                           out_buf_179_port, B2 => n690, Z => n576);
   U1408 : NAN4D1 port map( A1 => n579, A2 => n578, A3 => n577, A4 => n576, Z 
                           => N2879);
   U1409 : AOI22D1 port map( A1 => out_buf_84_port, A2 => n269, B1 => 
                           out_buf_20_port, B2 => n244, Z => n583);
   U1410 : AOI22D1 port map( A1 => out_buf_212_port, A2 => n270, B1 => 
                           out_buf_148_port, B2 => n245, Z => n582);
   U1411 : AOI22D1 port map( A1 => out_buf_116_port, A2 => n689, B1 => 
                           out_buf_52_port, B2 => n688, Z => n581);
   U1412 : AOI22D1 port map( A1 => out_buf_244_port, A2 => n691, B1 => 
                           out_buf_180_port, B2 => n690, Z => n580);
   U1413 : NAN4D1 port map( A1 => n583, A2 => n582, A3 => n581, A4 => n580, Z 
                           => N2878);
   U1414 : AOI22D1 port map( A1 => out_buf_85_port, A2 => n269, B1 => 
                           out_buf_21_port, B2 => n244, Z => n587);
   U1415 : AOI22D1 port map( A1 => out_buf_213_port, A2 => n270, B1 => 
                           out_buf_149_port, B2 => n245, Z => n586);
   U1416 : AOI22D1 port map( A1 => out_buf_117_port, A2 => n689, B1 => 
                           out_buf_53_port, B2 => n688, Z => n585);
   U1417 : AOI22D1 port map( A1 => out_buf_245_port, A2 => n691, B1 => 
                           out_buf_181_port, B2 => n690, Z => n584);
   U1418 : NAN4D1 port map( A1 => n587, A2 => n586, A3 => n585, A4 => n584, Z 
                           => N2877);
   U1419 : AOI22D1 port map( A1 => out_buf_86_port, A2 => n269, B1 => 
                           out_buf_22_port, B2 => n244, Z => n591);
   U1420 : AOI22D1 port map( A1 => out_buf_214_port, A2 => n270, B1 => 
                           out_buf_150_port, B2 => n245, Z => n5901);
   U1421 : AOI22D1 port map( A1 => out_buf_118_port, A2 => n689, B1 => 
                           out_buf_54_port, B2 => n688, Z => n589);
   U1422 : AOI22D1 port map( A1 => out_buf_246_port, A2 => n691, B1 => 
                           out_buf_182_port, B2 => n690, Z => n588);
   U1423 : NAN4D1 port map( A1 => n591, A2 => n5901, A3 => n589, A4 => n588, Z 
                           => N2876);
   U1424 : AOI22D1 port map( A1 => out_buf_87_port, A2 => n269, B1 => 
                           out_buf_23_port, B2 => n244, Z => n595);
   U1425 : AOI22D1 port map( A1 => out_buf_215_port, A2 => n270, B1 => 
                           out_buf_151_port, B2 => n245, Z => n594);
   U1426 : AOI22D1 port map( A1 => out_buf_119_port, A2 => n689, B1 => 
                           out_buf_55_port, B2 => n688, Z => n593);
   U1427 : AOI22D1 port map( A1 => out_buf_247_port, A2 => n691, B1 => 
                           out_buf_183_port, B2 => n690, Z => n592);
   U1428 : NAN4D1 port map( A1 => n595, A2 => n594, A3 => n593, A4 => n592, Z 
                           => N2875);
   U1429 : AOI22D1 port map( A1 => out_buf_88_port, A2 => n269, B1 => 
                           out_buf_24_port, B2 => n244, Z => n599);
   U1430 : AOI22D1 port map( A1 => out_buf_216_port, A2 => n270, B1 => 
                           out_buf_152_port, B2 => n245, Z => n598);
   U1431 : AOI22D1 port map( A1 => out_buf_120_port, A2 => n689, B1 => 
                           out_buf_56_port, B2 => n688, Z => n597);
   U1432 : AOI22D1 port map( A1 => out_buf_248_port, A2 => n691, B1 => 
                           out_buf_184_port, B2 => n690, Z => n596);
   U1433 : NAN4D1 port map( A1 => n599, A2 => n598, A3 => n597, A4 => n596, Z 
                           => N2874);
   U1434 : AOI22D1 port map( A1 => out_buf_89_port, A2 => n269, B1 => 
                           out_buf_25_port, B2 => n244, Z => n603);
   U1435 : AOI22D1 port map( A1 => out_buf_217_port, A2 => n270, B1 => 
                           out_buf_153_port, B2 => n245, Z => n602);
   U1436 : AOI22D1 port map( A1 => out_buf_121_port, A2 => n689, B1 => 
                           out_buf_57_port, B2 => n688, Z => n601);
   U1437 : AOI22D1 port map( A1 => out_buf_249_port, A2 => n691, B1 => 
                           out_buf_185_port, B2 => n690, Z => n6001);
   U1438 : NAN4D1 port map( A1 => n603, A2 => n602, A3 => n601, A4 => n6001, Z 
                           => N2873);
   U1439 : AOI22D1 port map( A1 => out_buf_90_port, A2 => n269, B1 => 
                           out_buf_26_port, B2 => n244, Z => n607);
   U1440 : AOI22D1 port map( A1 => out_buf_218_port, A2 => n270, B1 => 
                           out_buf_154_port, B2 => n245, Z => n606);
   U1441 : AOI22D1 port map( A1 => out_buf_122_port, A2 => n689, B1 => 
                           out_buf_58_port, B2 => n688, Z => n605);
   U1442 : AOI22D1 port map( A1 => out_buf_250_port, A2 => n691, B1 => 
                           out_buf_186_port, B2 => n690, Z => n604);
   U1443 : NAN4D1 port map( A1 => n607, A2 => n606, A3 => n605, A4 => n604, Z 
                           => N2872);
   U1444 : AOI22D1 port map( A1 => out_buf_91_port, A2 => n269, B1 => 
                           out_buf_27_port, B2 => n244, Z => n611);
   U1445 : AOI22D1 port map( A1 => out_buf_219_port, A2 => n270, B1 => 
                           out_buf_155_port, B2 => n245, Z => n6101);
   U1446 : AOI22D1 port map( A1 => out_buf_123_port, A2 => n689, B1 => 
                           out_buf_59_port, B2 => n688, Z => n609);
   U1447 : AOI22D1 port map( A1 => out_buf_251_port, A2 => n691, B1 => 
                           out_buf_187_port, B2 => n690, Z => n608);
   U1448 : NAN4D1 port map( A1 => n611, A2 => n6101, A3 => n609, A4 => n608, Z 
                           => N2871);
   U1449 : AOI22D1 port map( A1 => out_buf_92_port, A2 => n269, B1 => 
                           out_buf_28_port, B2 => n244, Z => n615);
   U1450 : AOI22D1 port map( A1 => out_buf_220_port, A2 => n270, B1 => 
                           out_buf_156_port, B2 => n245, Z => n614);
   U1451 : AOI22D1 port map( A1 => out_buf_124_port, A2 => n689, B1 => 
                           out_buf_60_port, B2 => n688, Z => n613);
   U1452 : AOI22D1 port map( A1 => out_buf_252_port, A2 => n691, B1 => 
                           out_buf_188_port, B2 => n690, Z => n612);
   U1453 : NAN4D1 port map( A1 => n615, A2 => n614, A3 => n613, A4 => n612, Z 
                           => N2870);
   U1454 : AOI22D1 port map( A1 => out_buf_93_port, A2 => n269, B1 => 
                           out_buf_29_port, B2 => n244, Z => n619);
   U1455 : AOI22D1 port map( A1 => out_buf_221_port, A2 => n270, B1 => 
                           out_buf_157_port, B2 => n245, Z => n618);
   U1456 : AOI22D1 port map( A1 => out_buf_125_port, A2 => n689, B1 => 
                           out_buf_61_port, B2 => n688, Z => n617);
   U1457 : AOI22D1 port map( A1 => out_buf_253_port, A2 => n691, B1 => 
                           out_buf_189_port, B2 => n690, Z => n616);
   U1458 : NAN4D1 port map( A1 => n619, A2 => n618, A3 => n617, A4 => n616, Z 
                           => N2869);
   U1459 : AOI22D1 port map( A1 => out_buf_94_port, A2 => n269, B1 => 
                           out_buf_30_port, B2 => n244, Z => n623);
   U1460 : AOI22D1 port map( A1 => out_buf_222_port, A2 => n270, B1 => 
                           out_buf_158_port, B2 => n245, Z => n622);
   U1461 : AOI22D1 port map( A1 => out_buf_126_port, A2 => n689, B1 => 
                           out_buf_62_port, B2 => n688, Z => n621);
   U1462 : AOI22D1 port map( A1 => out_buf_254_port, A2 => n691, B1 => 
                           out_buf_190_port, B2 => n690, Z => n620);
   U1463 : NAN4D1 port map( A1 => n623, A2 => n622, A3 => n621, A4 => n620, Z 
                           => N2868);
   U1464 : AOI22D1 port map( A1 => out_buf_95_port, A2 => n269, B1 => 
                           out_buf_31_port, B2 => n244, Z => n627);
   U1465 : AOI22D1 port map( A1 => out_buf_223_port, A2 => n270, B1 => 
                           out_buf_159_port, B2 => n245, Z => n626);
   U1466 : AOI22D1 port map( A1 => out_buf_127_port, A2 => n689, B1 => 
                           out_buf_63_port, B2 => n688, Z => n625);
   U1467 : AOI22D1 port map( A1 => out_buf_255_port, A2 => n691, B1 => 
                           out_buf_191_port, B2 => n690, Z => n624);
   U1468 : NAN4D1 port map( A1 => n627, A2 => n626, A3 => n625, A4 => n624, Z 
                           => N2867);
   U1469 : AOI22D1 port map( A1 => out_buf_64_port, A2 => n269, B1 => 
                           out_buf_0_port, B2 => n244, Z => n631);
   U1470 : AOI22D1 port map( A1 => out_buf_192_port, A2 => n270, B1 => 
                           out_buf_128_port, B2 => n245, Z => n6301);
   U1471 : AOI22D1 port map( A1 => out_buf_96_port, A2 => n689, B1 => 
                           out_buf_32_port, B2 => n688, Z => n629);
   U1472 : AOI22D1 port map( A1 => out_buf_224_port, A2 => n691, B1 => 
                           out_buf_160_port, B2 => n690, Z => n628);
   U1473 : NAN4D1 port map( A1 => n631, A2 => n6301, A3 => n629, A4 => n628, Z 
                           => N2865);
   U1474 : AOI22D1 port map( A1 => out_buf_65_port, A2 => n269, B1 => 
                           out_buf_1_port, B2 => n244, Z => n635);
   U1475 : AOI22D1 port map( A1 => out_buf_193_port, A2 => n270, B1 => 
                           out_buf_129_port, B2 => n245, Z => n634);
   U1476 : AOI22D1 port map( A1 => out_buf_97_port, A2 => n689, B1 => 
                           out_buf_33_port, B2 => n688, Z => n633);
   U1477 : AOI22D1 port map( A1 => out_buf_225_port, A2 => n691, B1 => 
                           out_buf_161_port, B2 => n690, Z => n632);
   U1478 : NAN4D1 port map( A1 => n635, A2 => n634, A3 => n633, A4 => n632, Z 
                           => N2864);
   U1479 : AOI22D1 port map( A1 => out_buf_66_port, A2 => n269, B1 => 
                           out_buf_2_port, B2 => n244, Z => n639);
   U1480 : AOI22D1 port map( A1 => out_buf_194_port, A2 => n270, B1 => 
                           out_buf_130_port, B2 => n245, Z => n638);
   U1481 : AOI22D1 port map( A1 => out_buf_98_port, A2 => n689, B1 => 
                           out_buf_34_port, B2 => n688, Z => n637);
   U1482 : AOI22D1 port map( A1 => out_buf_226_port, A2 => n691, B1 => 
                           out_buf_162_port, B2 => n690, Z => n636);
   U1483 : NAN4D1 port map( A1 => n639, A2 => n638, A3 => n637, A4 => n636, Z 
                           => N2863);
   U1484 : AOI22D1 port map( A1 => out_buf_67_port, A2 => n269, B1 => 
                           out_buf_3_port, B2 => n244, Z => n643);
   U1485 : AOI22D1 port map( A1 => out_buf_195_port, A2 => n270, B1 => 
                           out_buf_131_port, B2 => n245, Z => n642);
   U1486 : AOI22D1 port map( A1 => out_buf_99_port, A2 => n689, B1 => 
                           out_buf_35_port, B2 => n688, Z => n641);
   U1487 : AOI22D1 port map( A1 => out_buf_227_port, A2 => n691, B1 => 
                           out_buf_163_port, B2 => n690, Z => n6401);
   U1488 : NAN4D1 port map( A1 => n643, A2 => n642, A3 => n641, A4 => n6401, Z 
                           => N2862);
   U1489 : AOI22D1 port map( A1 => out_buf_68_port, A2 => n269, B1 => 
                           out_buf_4_port, B2 => n244, Z => n647);
   U1490 : AOI22D1 port map( A1 => out_buf_196_port, A2 => n270, B1 => 
                           out_buf_132_port, B2 => n245, Z => n646);
   U1491 : AOI22D1 port map( A1 => out_buf_100_port, A2 => n689, B1 => 
                           out_buf_36_port, B2 => n688, Z => n645);
   U1492 : AOI22D1 port map( A1 => out_buf_228_port, A2 => n691, B1 => 
                           out_buf_164_port, B2 => n690, Z => n644);
   U1493 : NAN4D1 port map( A1 => n647, A2 => n646, A3 => n645, A4 => n644, Z 
                           => N2861);
   U1494 : AOI22D1 port map( A1 => out_buf_69_port, A2 => n269, B1 => 
                           out_buf_5_port, B2 => n244, Z => n651);
   U1495 : AOI22D1 port map( A1 => out_buf_197_port, A2 => n270, B1 => 
                           out_buf_133_port, B2 => n245, Z => n650);
   U1496 : AOI22D1 port map( A1 => out_buf_101_port, A2 => n689, B1 => 
                           out_buf_37_port, B2 => n688, Z => n649);
   U1497 : AOI22D1 port map( A1 => out_buf_229_port, A2 => n691, B1 => 
                           out_buf_165_port, B2 => n690, Z => n648);
   U1498 : NAN4D1 port map( A1 => n651, A2 => n650, A3 => n649, A4 => n648, Z 
                           => N2860);
   U1499 : AOI22D1 port map( A1 => out_buf_70_port, A2 => n269, B1 => 
                           out_buf_6_port, B2 => n244, Z => n655);
   U1500 : AOI22D1 port map( A1 => out_buf_198_port, A2 => n270, B1 => 
                           out_buf_134_port, B2 => n245, Z => n654);
   U1501 : AOI22D1 port map( A1 => out_buf_102_port, A2 => n689, B1 => 
                           out_buf_38_port, B2 => n688, Z => n653);
   U1502 : AOI22D1 port map( A1 => out_buf_230_port, A2 => n691, B1 => 
                           out_buf_166_port, B2 => n690, Z => n652);
   U1503 : NAN4D1 port map( A1 => n655, A2 => n654, A3 => n653, A4 => n652, Z 
                           => N2859);
   U1504 : AOI22D1 port map( A1 => out_buf_71_port, A2 => n269, B1 => 
                           out_buf_7_port, B2 => n244, Z => n659);
   U1505 : AOI22D1 port map( A1 => out_buf_199_port, A2 => n270, B1 => 
                           out_buf_135_port, B2 => n245, Z => n658);
   U1506 : AOI22D1 port map( A1 => out_buf_103_port, A2 => n689, B1 => 
                           out_buf_39_port, B2 => n688, Z => n657);
   U1507 : AOI22D1 port map( A1 => out_buf_231_port, A2 => n691, B1 => 
                           out_buf_167_port, B2 => n690, Z => n656);
   U1508 : NAN4D1 port map( A1 => n659, A2 => n658, A3 => n657, A4 => n656, Z 
                           => N2858);
   U1509 : AOI22D1 port map( A1 => out_buf_72_port, A2 => n269, B1 => 
                           out_buf_8_port, B2 => n244, Z => n663);
   U1510 : AOI22D1 port map( A1 => out_buf_200_port, A2 => n270, B1 => 
                           out_buf_136_port, B2 => n245, Z => n662);
   U1511 : AOI22D1 port map( A1 => out_buf_104_port, A2 => n689, B1 => 
                           out_buf_40_port, B2 => n688, Z => n661);
   U1512 : AOI22D1 port map( A1 => out_buf_232_port, A2 => n691, B1 => 
                           out_buf_168_port, B2 => n690, Z => n660);
   U1513 : NAN4D1 port map( A1 => n663, A2 => n662, A3 => n661, A4 => n660, Z 
                           => N2857);
   U1514 : AOI22D1 port map( A1 => out_buf_73_port, A2 => n269, B1 => 
                           out_buf_9_port, B2 => n244, Z => n667);
   U1515 : AOI22D1 port map( A1 => out_buf_201_port, A2 => n270, B1 => 
                           out_buf_137_port, B2 => n245, Z => n666);
   U1516 : AOI22D1 port map( A1 => out_buf_105_port, A2 => n689, B1 => 
                           out_buf_41_port, B2 => n688, Z => n665);
   U1517 : AOI22D1 port map( A1 => out_buf_233_port, A2 => n691, B1 => 
                           out_buf_169_port, B2 => n690, Z => n664);
   U1518 : NAN4D1 port map( A1 => n667, A2 => n666, A3 => n665, A4 => n664, Z 
                           => N2856);
   U1519 : AOI22D1 port map( A1 => out_buf_74_port, A2 => n269, B1 => 
                           out_buf_10_port, B2 => n244, Z => n671);
   U1520 : AOI22D1 port map( A1 => out_buf_202_port, A2 => n270, B1 => 
                           out_buf_138_port, B2 => n245, Z => n670);
   U1521 : AOI22D1 port map( A1 => out_buf_106_port, A2 => n689, B1 => 
                           out_buf_42_port, B2 => n688, Z => n669);
   U1522 : AOI22D1 port map( A1 => out_buf_234_port, A2 => n691, B1 => 
                           out_buf_170_port, B2 => n690, Z => n668);
   U1523 : NAN4D1 port map( A1 => n671, A2 => n670, A3 => n669, A4 => n668, Z 
                           => N2855);
   U1524 : AOI22D1 port map( A1 => out_buf_75_port, A2 => n269, B1 => 
                           out_buf_11_port, B2 => n244, Z => n675);
   U1525 : AOI22D1 port map( A1 => out_buf_203_port, A2 => n270, B1 => 
                           out_buf_139_port, B2 => n245, Z => n674);
   U1526 : AOI22D1 port map( A1 => out_buf_107_port, A2 => n689, B1 => 
                           out_buf_43_port, B2 => n688, Z => n673);
   U1527 : AOI22D1 port map( A1 => out_buf_235_port, A2 => n691, B1 => 
                           out_buf_171_port, B2 => n690, Z => n672);
   U1528 : NAN4D1 port map( A1 => n675, A2 => n674, A3 => n673, A4 => n672, Z 
                           => N2854);
   U1529 : AOI22D1 port map( A1 => out_buf_76_port, A2 => n269, B1 => 
                           out_buf_12_port, B2 => n244, Z => n679);
   U1530 : AOI22D1 port map( A1 => out_buf_204_port, A2 => n270, B1 => 
                           out_buf_140_port, B2 => n245, Z => n678);
   U1531 : AOI22D1 port map( A1 => out_buf_108_port, A2 => n689, B1 => 
                           out_buf_44_port, B2 => n688, Z => n677);
   U1532 : AOI22D1 port map( A1 => out_buf_236_port, A2 => n691, B1 => 
                           out_buf_172_port, B2 => n690, Z => n676);
   U1533 : NAN4D1 port map( A1 => n679, A2 => n678, A3 => n677, A4 => n676, Z 
                           => N2853);
   U1534 : AOI22D1 port map( A1 => out_buf_77_port, A2 => n269, B1 => 
                           out_buf_13_port, B2 => n244, Z => n683);
   U1535 : AOI22D1 port map( A1 => out_buf_205_port, A2 => n270, B1 => 
                           out_buf_141_port, B2 => n245, Z => n682);
   U1536 : AOI22D1 port map( A1 => out_buf_109_port, A2 => n689, B1 => 
                           out_buf_45_port, B2 => n688, Z => n681);
   U1537 : AOI22D1 port map( A1 => out_buf_237_port, A2 => n691, B1 => 
                           out_buf_173_port, B2 => n690, Z => n680);
   U1538 : NAN4D1 port map( A1 => n683, A2 => n682, A3 => n681, A4 => n680, Z 
                           => N2852);
   U1539 : AOI22D1 port map( A1 => out_buf_78_port, A2 => n269, B1 => 
                           out_buf_14_port, B2 => n244, Z => n687);
   U1540 : AOI22D1 port map( A1 => out_buf_206_port, A2 => n270, B1 => 
                           out_buf_142_port, B2 => n245, Z => n686);
   U1541 : AOI22D1 port map( A1 => out_buf_110_port, A2 => n689, B1 => 
                           out_buf_46_port, B2 => n688, Z => n685);
   U1542 : AOI22D1 port map( A1 => out_buf_238_port, A2 => n691, B1 => 
                           out_buf_174_port, B2 => n690, Z => n684);
   U1543 : NAN4D1 port map( A1 => n687, A2 => n686, A3 => n685, A4 => n684, Z 
                           => N2851);
   U1544 : AOI22D1 port map( A1 => out_buf_79_port, A2 => n269, B1 => 
                           out_buf_15_port, B2 => n244, Z => n695);
   U1545 : AOI22D1 port map( A1 => out_buf_207_port, A2 => n270, B1 => 
                           out_buf_143_port, B2 => n245, Z => n694);
   U1546 : AOI22D1 port map( A1 => out_buf_111_port, A2 => n689, B1 => 
                           out_buf_47_port, B2 => n688, Z => n693);
   U1547 : AOI22D1 port map( A1 => out_buf_239_port, A2 => n691, B1 => 
                           out_buf_175_port, B2 => n690, Z => n692);
   U1548 : NAN4D1 port map( A1 => n695, A2 => n694, A3 => n693, A4 => n692, Z 
                           => N2850);
   U1549 : NAN2D1 port map( A1 => n114, A2 => avs_addr(3), Z => n6400);
   U1550 : NAN3D1 port map( A1 => avs_write, A2 => n277, A3 => n795, Z => n178)
                           ;
   U1551 : NAN2D1 port map( A1 => operand_regs_255_port, A2 => n709, Z => n763)
                           ;
   U1552 : OAI21D1 port map( A1 => n713, A2 => n730, B => n763, Z => N3104);
   U1553 : NAN2D1 port map( A1 => operand_regs_254_port, A2 => n709, Z => n764)
                           ;
   U1554 : OAI21D1 port map( A1 => n706, A2 => n731, B => n764, Z => N3103);
   U1555 : NAN2D1 port map( A1 => operand_regs_253_port, A2 => n709, Z => n765)
                           ;
   U1556 : OAI21D1 port map( A1 => n708, A2 => n732, B => n765, Z => N3102);
   U1557 : NAN2D1 port map( A1 => operand_regs_252_port, A2 => n709, Z => n766)
                           ;
   U1558 : OAI21D1 port map( A1 => n706, A2 => n733, B => n766, Z => N3101);
   U1559 : NAN2D1 port map( A1 => operand_regs_251_port, A2 => n709, Z => n767)
                           ;
   U1560 : OAI21D1 port map( A1 => n706, A2 => n734, B => n767, Z => N3100);
   U1561 : NAN2D1 port map( A1 => operand_regs_250_port, A2 => n709, Z => n768)
                           ;
   U1562 : OAI21D1 port map( A1 => n713, A2 => n735, B => n768, Z => N3099);
   U1563 : NAN2D1 port map( A1 => operand_regs_249_port, A2 => n709, Z => n769)
                           ;
   U1564 : OAI21D1 port map( A1 => n707, A2 => n736, B => n769, Z => N3098);
   U1565 : NAN2D1 port map( A1 => operand_regs_248_port, A2 => n709, Z => n770)
                           ;
   U1566 : OAI21D1 port map( A1 => n708, A2 => n737, B => n770, Z => N3097);
   U1567 : NAN2D1 port map( A1 => operand_regs_247_port, A2 => n709, Z => n771)
                           ;
   U1568 : OAI21D1 port map( A1 => n707, A2 => n738, B => n771, Z => N3096);
   U1569 : NAN2D1 port map( A1 => operand_regs_246_port, A2 => n709, Z => n772)
                           ;
   U1570 : OAI21D1 port map( A1 => n713, A2 => n739, B => n772, Z => N3095);
   U1571 : NAN2D1 port map( A1 => operand_regs_245_port, A2 => n709, Z => n773)
                           ;
   U1572 : OAI21D1 port map( A1 => n707, A2 => n740, B => n773, Z => N3094);
   U1573 : NAN2D1 port map( A1 => operand_regs_244_port, A2 => n708, Z => n774)
                           ;
   U1574 : OAI21D1 port map( A1 => n707, A2 => n741, B => n774, Z => N3093);
   U1575 : NAN2D1 port map( A1 => operand_regs_243_port, A2 => n708, Z => n775)
                           ;
   U1576 : OAI21D1 port map( A1 => n707, A2 => n742, B => n775, Z => N3092);
   U1577 : NAN2D1 port map( A1 => operand_regs_242_port, A2 => n708, Z => n776)
                           ;
   U1578 : OAI21D1 port map( A1 => n707, A2 => n743, B => n776, Z => N3091);
   U1579 : NAN2D1 port map( A1 => operand_regs_241_port, A2 => n708, Z => n777)
                           ;
   U1580 : OAI21D1 port map( A1 => n708, A2 => n744, B => n777, Z => N3090);
   U1581 : NAN2D1 port map( A1 => operand_regs_240_port, A2 => n708, Z => n778)
                           ;
   U1582 : OAI21D1 port map( A1 => n706, A2 => n745, B => n778, Z => N3089);
   U1583 : NAN2D1 port map( A1 => operand_regs_239_port, A2 => n708, Z => n779)
                           ;
   U1584 : OAI21D1 port map( A1 => n708, A2 => n746, B => n779, Z => N3088);
   U1585 : NAN2D1 port map( A1 => operand_regs_238_port, A2 => n708, Z => n780)
                           ;
   U1586 : OAI21D1 port map( A1 => n706, A2 => n747, B => n780, Z => N3087);
   U1587 : NAN2D1 port map( A1 => operand_regs_237_port, A2 => n708, Z => n781)
                           ;
   U1588 : OAI21D1 port map( A1 => n708, A2 => n748, B => n781, Z => N3086);
   U1589 : NAN2D1 port map( A1 => operand_regs_236_port, A2 => n707, Z => n782)
                           ;
   U1590 : OAI21D1 port map( A1 => n708, A2 => n749, B => n782, Z => N3085);
   U1591 : NAN2D1 port map( A1 => operand_regs_235_port, A2 => n708, Z => n783)
                           ;
   U1592 : OAI21D1 port map( A1 => n713, A2 => n750, B => n783, Z => N3084);
   U1593 : NAN2D1 port map( A1 => operand_regs_234_port, A2 => n708, Z => n784)
                           ;
   U1594 : OAI21D1 port map( A1 => n708, A2 => n751, B => n784, Z => N3083);
   U1595 : NAN2D1 port map( A1 => operand_regs_233_port, A2 => n708, Z => n785)
                           ;
   U1596 : OAI21D1 port map( A1 => n713, A2 => n752, B => n785, Z => N3082);
   U1597 : NAN2D1 port map( A1 => operand_regs_232_port, A2 => n707, Z => n786)
                           ;
   U1598 : OAI21D1 port map( A1 => n708, A2 => n753, B => n786, Z => N3081);
   U1599 : NAN2D1 port map( A1 => operand_regs_231_port, A2 => n708, Z => n787)
                           ;
   U1600 : OAI21D1 port map( A1 => n706, A2 => n754, B => n787, Z => N3080);
   U1601 : NAN2D1 port map( A1 => operand_regs_230_port, A2 => n707, Z => n788)
                           ;
   U1602 : OAI21D1 port map( A1 => n706, A2 => n755, B => n788, Z => N3079);
   U1603 : NAN2D1 port map( A1 => operand_regs_229_port, A2 => n708, Z => n789)
                           ;
   U1604 : OAI21D1 port map( A1 => n706, A2 => n756, B => n789, Z => N3078);
   U1605 : NAN2D1 port map( A1 => operand_regs_228_port, A2 => n707, Z => n790)
                           ;
   U1606 : OAI21D1 port map( A1 => n706, A2 => n757, B => n790, Z => N3077);
   U1607 : NAN2D1 port map( A1 => operand_regs_227_port, A2 => n707, Z => n791)
                           ;
   U1608 : OAI21D1 port map( A1 => n706, A2 => n758, B => n791, Z => N3076);
   U1609 : NAN2D1 port map( A1 => operand_regs_226_port, A2 => n708, Z => n792)
                           ;
   U1610 : OAI21D1 port map( A1 => n706, A2 => n759, B => n792, Z => N3075);
   U1611 : NAN2D1 port map( A1 => operand_regs_225_port, A2 => n707, Z => n793)
                           ;
   U1612 : OAI21D1 port map( A1 => n706, A2 => n760, B => n793, Z => N3074);
   U1613 : NAN2D1 port map( A1 => operand_regs_224_port, A2 => n707, Z => n794)
                           ;
   U1614 : OAI21D1 port map( A1 => n706, A2 => n761, B => n794, Z => N3073);
   U1615 : OAI21M20D1 port map( A1 => operand_regs_159_port, A2 => n726, B => 
                           n763, Z => N3136);
   U1616 : OAI21M20D1 port map( A1 => operand_regs_158_port, A2 => n726, B => 
                           n764, Z => N3135);
   U1617 : OAI21M20D1 port map( A1 => operand_regs_157_port, A2 => n726, B => 
                           n765, Z => N3134);
   U1618 : OAI21M20D1 port map( A1 => operand_regs_156_port, A2 => n726, B => 
                           n766, Z => N3133);
   U1619 : OAI21M20D1 port map( A1 => operand_regs_155_port, A2 => n726, B => 
                           n767, Z => N3132);
   U1620 : OAI21M20D1 port map( A1 => operand_regs_154_port, A2 => n728, B => 
                           n768, Z => N3131);
   U1621 : OAI21M20D1 port map( A1 => operand_regs_153_port, A2 => n728, B => 
                           n769, Z => N3130);
   U1622 : OAI21M20D1 port map( A1 => operand_regs_152_port, A2 => n728, B => 
                           n770, Z => N3129);
   U1623 : OAI21M20D1 port map( A1 => operand_regs_151_port, A2 => n728, B => 
                           n771, Z => N3128);
   U1624 : OAI21M20D1 port map( A1 => operand_regs_150_port, A2 => n727, B => 
                           n772, Z => N3127);
   U1625 : OAI21M20D1 port map( A1 => operand_regs_149_port, A2 => n728, B => 
                           n773, Z => N3126);
   U1626 : OAI21M20D1 port map( A1 => operand_regs_148_port, A2 => n728, B => 
                           n774, Z => N3125);
   U1627 : OAI21M20D1 port map( A1 => operand_regs_147_port, A2 => n727, B => 
                           n775, Z => N3124);
   U1628 : OAI21M20D1 port map( A1 => operand_regs_146_port, A2 => n727, B => 
                           n776, Z => N3123);
   U1629 : OAI21M20D1 port map( A1 => operand_regs_145_port, A2 => n727, B => 
                           n777, Z => N3122);
   U1630 : OAI21M20D1 port map( A1 => operand_regs_144_port, A2 => n728, B => 
                           n778, Z => N3121);
   U1631 : OAI21M20D1 port map( A1 => operand_regs_143_port, A2 => n727, B => 
                           n779, Z => N3120);
   U1632 : OAI21M20D1 port map( A1 => operand_regs_142_port, A2 => n727, B => 
                           n780, Z => N3119);
   U1633 : OAI21M20D1 port map( A1 => operand_regs_141_port, A2 => n728, B => 
                           n781, Z => N3118);
   U1634 : OAI21M20D1 port map( A1 => operand_regs_140_port, A2 => n727, B => 
                           n782, Z => N3117);
   U1635 : OAI21M20D1 port map( A1 => operand_regs_139_port, A2 => n728, B => 
                           n783, Z => N3116);
   U1636 : OAI21M20D1 port map( A1 => operand_regs_138_port, A2 => n727, B => 
                           n784, Z => N3115);
   U1637 : OAI21M20D1 port map( A1 => operand_regs_137_port, A2 => n728, B => 
                           n785, Z => N3114);
   U1638 : OAI21M20D1 port map( A1 => operand_regs_136_port, A2 => n727, B => 
                           n786, Z => N3113);
   U1639 : OAI21M20D1 port map( A1 => operand_regs_135_port, A2 => n727, B => 
                           n787, Z => N3112);
   U1640 : OAI21M20D1 port map( A1 => operand_regs_134_port, A2 => n727, B => 
                           n788, Z => N3111);
   U1641 : OAI21M20D1 port map( A1 => operand_regs_133_port, A2 => n727, B => 
                           n789, Z => N3110);
   U1642 : OAI21M20D1 port map( A1 => operand_regs_132_port, A2 => n727, B => 
                           n790, Z => N3109);
   U1643 : OAI21M20D1 port map( A1 => operand_regs_131_port, A2 => n727, B => 
                           n791, Z => N3108);
   U1644 : OAI21M20D1 port map( A1 => operand_regs_130_port, A2 => n727, B => 
                           n792, Z => N3107);
   U1645 : OAI21M20D1 port map( A1 => operand_regs_129_port, A2 => n727, B => 
                           n793, Z => N3106);
   U1646 : OAI21M20D1 port map( A1 => operand_regs_128_port, A2 => n727, B => 
                           n794, Z => N3105);
   U1647 : OAI21M20D1 port map( A1 => operand_regs_95_port, A2 => n728, B => 
                           n763, Z => N3168);
   U1648 : OAI21M20D1 port map( A1 => operand_regs_94_port, A2 => n727, B => 
                           n764, Z => N3167);
   U1649 : OAI21M20D1 port map( A1 => operand_regs_93_port, A2 => n728, B => 
                           n765, Z => N3166);
   U1650 : OAI21M20D1 port map( A1 => operand_regs_92_port, A2 => n727, B => 
                           n766, Z => N3165);
   U1651 : OAI21M20D1 port map( A1 => operand_regs_91_port, A2 => n728, B => 
                           n767, Z => N3164);
   U1652 : OAI21M20D1 port map( A1 => operand_regs_90_port, A2 => n728, B => 
                           n768, Z => N3163);
   U1653 : OAI21M20D1 port map( A1 => operand_regs_89_port, A2 => n727, B => 
                           n769, Z => N3162);
   U1654 : OAI21M20D1 port map( A1 => operand_regs_88_port, A2 => n727, B => 
                           n770, Z => N3161);
   U1655 : OAI21M20D1 port map( A1 => operand_regs_87_port, A2 => n728, B => 
                           n771, Z => N3160);
   U1656 : OAI21M20D1 port map( A1 => operand_regs_86_port, A2 => n728, B => 
                           n772, Z => N3159);
   U1657 : OAI21M20D1 port map( A1 => operand_regs_85_port, A2 => n727, B => 
                           n773, Z => N3158);
   U1658 : OAI21M20D1 port map( A1 => operand_regs_84_port, A2 => n728, B => 
                           n774, Z => N3157);
   U1659 : OAI21M20D1 port map( A1 => operand_regs_83_port, A2 => n727, B => 
                           n775, Z => N3156);
   U1660 : OAI21M20D1 port map( A1 => operand_regs_82_port, A2 => n727, B => 
                           n776, Z => N3155);
   U1661 : OAI21M20D1 port map( A1 => operand_regs_81_port, A2 => n727, B => 
                           n777, Z => N3154);
   U1662 : OAI21M20D1 port map( A1 => operand_regs_80_port, A2 => n727, B => 
                           n778, Z => N3153);
   U1663 : OAI21M20D1 port map( A1 => operand_regs_79_port, A2 => n727, B => 
                           n779, Z => N3152);
   U1664 : OAI21M20D1 port map( A1 => operand_regs_78_port, A2 => n727, B => 
                           n780, Z => N3151);
   U1665 : OAI21M20D1 port map( A1 => operand_regs_77_port, A2 => n727, B => 
                           n781, Z => N3150);
   U1666 : OAI21M20D1 port map( A1 => operand_regs_76_port, A2 => n727, B => 
                           n782, Z => N3149);
   U1667 : OAI21M20D1 port map( A1 => operand_regs_75_port, A2 => n727, B => 
                           n783, Z => N3148);
   U1668 : OAI21M20D1 port map( A1 => operand_regs_74_port, A2 => n727, B => 
                           n784, Z => N3147);
   U1669 : OAI21M20D1 port map( A1 => operand_regs_73_port, A2 => n727, B => 
                           n785, Z => N3146);
   U1670 : OAI21M20D1 port map( A1 => operand_regs_72_port, A2 => n727, B => 
                           n786, Z => N3145);
   U1671 : OAI21M20D1 port map( A1 => operand_regs_71_port, A2 => n727, B => 
                           n787, Z => N3144);
   U1672 : OAI21M20D1 port map( A1 => operand_regs_70_port, A2 => n728, B => 
                           n788, Z => N3143);
   U1673 : OAI21M20D1 port map( A1 => operand_regs_69_port, A2 => n728, B => 
                           n789, Z => N3142);
   U1674 : OAI21M20D1 port map( A1 => operand_regs_68_port, A2 => n728, B => 
                           n790, Z => N3141);
   U1675 : OAI21M20D1 port map( A1 => operand_regs_67_port, A2 => n728, B => 
                           n791, Z => N3140);
   U1676 : OAI21M20D1 port map( A1 => operand_regs_66_port, A2 => n728, B => 
                           n792, Z => N3139);
   U1677 : OAI21M20D1 port map( A1 => operand_regs_65_port, A2 => n728, B => 
                           n793, Z => N3138);
   U1678 : OAI21M20D1 port map( A1 => operand_regs_64_port, A2 => n728, B => 
                           n794, Z => N3137);
   U1679 : NOR3D1 port map( A1 => avs_addr(3), A2 => avs_addr(5), A3 => 
                           avs_addr(4), Z => N66);
   mult_21_C241_U1395 : INVD1 port map( A => N2944, Z => mult_21_C241_n1066);
   mult_21_C241_U1394 : BUFD1 port map( A => N3084, Z => mult_21_C241_n1540);
   mult_21_C241_U1393 : BUFD1 port map( A => N3083, Z => mult_21_C241_n1539);
   mult_21_C241_U1392 : BUFD1 port map( A => N3082, Z => mult_21_C241_n1538);
   mult_21_C241_U1391 : INVD1 port map( A => N3073, Z => mult_21_C241_n1549);
   mult_21_C241_U1390 : INVD1 port map( A => N3075, Z => mult_21_C241_n1547);
   mult_21_C241_U1389 : AO21D1 port map( A1 => N2942, A2 => N2943, B => 
                           mult_21_C241_n1066, Z => mult_21_C241_n105);
   mult_21_C241_U1388 : INVD1 port map( A => N2942, Z => mult_21_C241_n1067);
   mult_21_C241_U1387 : AO21D1 port map( A1 => N2940, A2 => N2941, B => 
                           mult_21_C241_n1067, Z => mult_21_C241_n101);
   mult_21_C241_U1386 : EXOR2D1 port map( A1 => mult_21_C241_n1307, A2 => 
                           mult_21_C241_n1337, Z => mult_21_C241_n343);
   mult_21_C241_U1385 : INVD1 port map( A => N2940, Z => mult_21_C241_n1068);
   mult_21_C241_U1384 : AO21D1 port map( A1 => N2938, A2 => N2939, B => 
                           mult_21_C241_n1068, Z => mult_21_C241_n96);
   mult_21_C241_U1383 : ADHALFDL port map( A => mult_21_C241_n1309, B => 
                           mult_21_C241_n1339, CO => mult_21_C241_n400, S => 
                           mult_21_C241_n401);
   mult_21_C241_U1382 : AO21D1 port map( A1 => N2936, A2 => N2937, B => 
                           mult_21_C241_n1069, Z => mult_21_C241_n91);
   mult_21_C241_U1381 : INVD1 port map( A => N2938, Z => mult_21_C241_n1069);
   mult_21_C241_U1380 : ADHALFDL port map( A => mult_21_C241_n1311, B => 
                           mult_21_C241_n1341, CO => mult_21_C241_n454, S => 
                           mult_21_C241_n455);
   mult_21_C241_U1379 : OAI21D1 port map( A1 => N2936, A2 => N2937, B => 
                           mult_21_C241_n1069, Z => mult_21_C241_n89);
   mult_21_C241_U1378 : ADHALFDL port map( A => mult_21_C241_n1313, B => 
                           mult_21_C241_n1343, CO => mult_21_C241_n504, S => 
                           mult_21_C241_n505);
   mult_21_C241_U1377 : AO21D1 port map( A1 => N2934, A2 => N2935, B => 
                           mult_21_C241_n1070, Z => mult_21_C241_n86);
   mult_21_C241_U1376 : INVD1 port map( A => N2936, Z => mult_21_C241_n1070);
   mult_21_C241_U1375 : OAI21D1 port map( A1 => N2934, A2 => N2935, B => 
                           mult_21_C241_n1070, Z => mult_21_C241_n84);
   mult_21_C241_U1374 : AO21D1 port map( A1 => N2932, A2 => N2933, B => 
                           mult_21_C241_n1071, Z => mult_21_C241_n81);
   mult_21_C241_U1373 : INVD1 port map( A => N2934, Z => mult_21_C241_n1071);
   mult_21_C241_U1372 : OAI21D1 port map( A1 => N2932, A2 => N2933, B => 
                           mult_21_C241_n1071, Z => mult_21_C241_n79);
   mult_21_C241_U1371 : EXNOR2D1 port map( A1 => N2934, A2 => N2935, Z => 
                           mult_21_C241_n88);
   mult_21_C241_U1370 : AO21D1 port map( A1 => N2930, A2 => N2931, B => 
                           mult_21_C241_n1072, Z => mult_21_C241_n76);
   mult_21_C241_U1369 : OAI21D1 port map( A1 => N2922, A2 => N2923, B => 
                           mult_21_C241_n1076, Z => mult_21_C241_n42);
   mult_21_C241_U1368 : INVD1 port map( A => N2932, Z => mult_21_C241_n1072);
   mult_21_C241_U1367 : OAI21D1 port map( A1 => N2930, A2 => N2931, B => 
                           mult_21_C241_n1072, Z => mult_21_C241_n73);
   mult_21_C241_U1366 : INVD1 port map( A => N2924, Z => mult_21_C241_n1076);
   mult_21_C241_U1365 : AO21D1 port map( A1 => N2922, A2 => N2923, B => 
                           mult_21_C241_n1076, Z => mult_21_C241_n45);
   mult_21_C241_U1364 : OAI21D1 port map( A1 => N2928, A2 => N2929, B => 
                           mult_21_C241_n1073, Z => mult_21_C241_n66);
   mult_21_C241_U1363 : INVD1 port map( A => N2930, Z => mult_21_C241_n1073);
   mult_21_C241_U1362 : OAI21D1 port map( A1 => N2926, A2 => N2927, B => 
                           mult_21_C241_n1074, Z => mult_21_C241_n58);
   mult_21_C241_U1361 : INVD1 port map( A => N2928, Z => mult_21_C241_n1074);
   mult_21_C241_U1360 : AO21D1 port map( A1 => N2928, A2 => N2929, B => 
                           mult_21_C241_n1073, Z => mult_21_C241_n69);
   mult_21_C241_U1359 : AO21D1 port map( A1 => N2926, A2 => N2927, B => 
                           mult_21_C241_n1074, Z => mult_21_C241_n61);
   mult_21_C241_U1358 : OAI21D1 port map( A1 => N2924, A2 => N2925, B => 
                           mult_21_C241_n1075, Z => mult_21_C241_n50);
   mult_21_C241_U1357 : AO21D1 port map( A1 => N2920, A2 => N2921, B => 
                           mult_21_C241_n1077, Z => mult_21_C241_n38);
   mult_21_C241_U1356 : AO21D1 port map( A1 => N2916, A2 => N2917, B => 
                           mult_21_C241_n1079, Z => mult_21_C241_n22);
   mult_21_C241_U1355 : ADHALFDL port map( A => mult_21_C241_n1315, B => 
                           mult_21_C241_n1345, CO => mult_21_C241_n550, S => 
                           mult_21_C241_n551);
   mult_21_C241_U1354 : INVD1 port map( A => N2926, Z => mult_21_C241_n1075);
   mult_21_C241_U1353 : AO21D1 port map( A1 => N2924, A2 => N2925, B => 
                           mult_21_C241_n1075, Z => mult_21_C241_n53);
   mult_21_C241_U1352 : INVD1 port map( A => N2913, Z => mult_21_C241_n8);
   mult_21_C241_U1351 : EXNOR2D1 port map( A1 => N2932, A2 => N2933, Z => 
                           mult_21_C241_n83);
   mult_21_C241_U1350 : AO21D1 port map( A1 => N2918, A2 => N2919, B => 
                           mult_21_C241_n1078, Z => mult_21_C241_n30);
   mult_21_C241_U1349 : INVD1 port map( A => mult_21_C241_n1549, Z => 
                           mult_21_C241_n1548);
   mult_21_C241_U1348 : INVD1 port map( A => mult_21_C241_n1547, Z => 
                           mult_21_C241_n1546);
   mult_21_C241_U1347 : AO21D1 port map( A1 => N2914, A2 => N2915, B => 
                           mult_21_C241_n1080, Z => mult_21_C241_n14);
   mult_21_C241_U1346 : EXNOR2D1 port map( A1 => N2930, A2 => N2931, Z => 
                           mult_21_C241_n78);
   mult_21_C241_U1345 : EXNOR2D1 port map( A1 => N2922, A2 => N2923, Z => 
                           mult_21_C241_n48);
   mult_21_C241_U1344 : INVD1 port map( A => N2918, Z => mult_21_C241_n1079);
   mult_21_C241_U1343 : EXNOR2D1 port map( A1 => N2928, A2 => N2929, Z => 
                           mult_21_C241_n71);
   mult_21_C241_U1342 : EXNOR2D1 port map( A1 => N2926, A2 => N2927, Z => 
                           mult_21_C241_n63);
   mult_21_C241_U1341 : INVD1 port map( A => N2922, Z => mult_21_C241_n1077);
   mult_21_C241_U1340 : INVD1 port map( A => N2914, Z => mult_21_C241_n6);
   mult_21_C241_U1339 : NAN2D1 port map( A1 => N2913, A2 => mult_21_C241_n6, Z 
                           => mult_21_C241_n3);
   mult_21_C241_U1338 : INVD1 port map( A => N2920, Z => mult_21_C241_n1078);
   mult_21_C241_U1337 : EXNOR2D1 port map( A1 => N2924, A2 => N2925, Z => 
                           mult_21_C241_n56);
   mult_21_C241_U1336 : INVD1 port map( A => N2916, Z => mult_21_C241_n1080);
   mult_21_C241_U1335 : OA21D1 port map( A1 => N2918, A2 => N2919, B => 
                           mult_21_C241_n1078, Z => mult_21_C241_n1537);
   mult_21_C241_U1334 : ADHALFDL port map( A => mult_21_C241_n1325, B => 
                           mult_21_C241_n1355, CO => mult_21_C241_n720, S => 
                           mult_21_C241_n721);
   mult_21_C241_U1333 : ADHALFDL port map( A => mult_21_C241_n1321, B => 
                           mult_21_C241_n1351, CO => mult_21_C241_n664, S => 
                           mult_21_C241_n665);
   mult_21_C241_U1332 : ADHALFDL port map( A => mult_21_C241_n1319, B => 
                           mult_21_C241_n1349, CO => mult_21_C241_n630, S => 
                           mult_21_C241_n631);
   mult_21_C241_U1331 : ADHALFDL port map( A => mult_21_C241_n1327, B => 
                           mult_21_C241_n1357, CO => mult_21_C241_n742, S => 
                           mult_21_C241_n743);
   mult_21_C241_U1330 : ADHALFDL port map( A => mult_21_C241_n1317, B => 
                           mult_21_C241_n1347, CO => mult_21_C241_n592, S => 
                           mult_21_C241_n593);
   mult_21_C241_U1329 : EXOR2D1 port map( A1 => N2920, A2 => N2921, Z => 
                           mult_21_C241_n1536);
   mult_21_C241_U1328 : EXOR2D1 port map( A1 => N2916, A2 => N2917, Z => 
                           mult_21_C241_n1535);
   mult_21_C241_U1327 : EXOR2D1 port map( A1 => N2918, A2 => N2919, Z => 
                           mult_21_C241_n1534);
   mult_21_C241_U1326 : ADHALFDL port map( A => mult_21_C241_n1323, B => 
                           mult_21_C241_n1353, CO => mult_21_C241_n694, S => 
                           mult_21_C241_n695);
   mult_21_C241_U1325 : EXOR2D1 port map( A1 => N2914, A2 => N2915, Z => 
                           mult_21_C241_n1533);
   mult_21_C241_U1324 : ADHALFDL port map( A => mult_21_C241_n1329, B => 
                           mult_21_C241_n1359, CO => mult_21_C241_n760, S => 
                           mult_21_C241_n761);
   mult_21_C241_U1323 : ADHALFDL port map( A => mult_21_C241_n1098, B => 
                           mult_21_C241_n1081, CO => mult_21_C241_n372, S => 
                           mult_21_C241_n373);
   mult_21_C241_U1322 : ADHALFDL port map( A => mult_21_C241_n1102, B => 
                           mult_21_C241_n1082, CO => mult_21_C241_n428, S => 
                           mult_21_C241_n429);
   mult_21_C241_U1321 : ADHALFDL port map( A => mult_21_C241_n1108, B => 
                           mult_21_C241_n1083, CO => mult_21_C241_n480, S => 
                           mult_21_C241_n481);
   mult_21_C241_U1320 : ADHALFDL port map( A => mult_21_C241_n1116, B => 
                           mult_21_C241_n1084, CO => mult_21_C241_n528, S => 
                           mult_21_C241_n529);
   mult_21_C241_U1319 : ADHALFDL port map( A => mult_21_C241_n1126, B => 
                           mult_21_C241_n1085, CO => mult_21_C241_n572, S => 
                           mult_21_C241_n573);
   mult_21_C241_U1318 : INVD1 port map( A => mult_21_C241_n1367, Z => 
                           mult_21_C241_n303);
   mult_21_C241_U1317 : ADHALFDL port map( A => mult_21_C241_n1138, B => 
                           mult_21_C241_n1086, CO => mult_21_C241_n612, S => 
                           mult_21_C241_n613);
   mult_21_C241_U1316 : ADHALFDL port map( A => mult_21_C241_n1186, B => 
                           mult_21_C241_n1089, CO => mult_21_C241_n708, S => 
                           mult_21_C241_n709);
   mult_21_C241_U1315 : ADHALFDL port map( A => mult_21_C241_n1228, B => 
                           mult_21_C241_n1091, CO => mult_21_C241_n752, S => 
                           mult_21_C241_n753);
   mult_21_C241_U1314 : ADHALFDL port map( A => mult_21_C241_n1152, B => 
                           mult_21_C241_n1087, CO => mult_21_C241_n648, S => 
                           mult_21_C241_n649);
   mult_21_C241_U1313 : ADHALFDL port map( A => mult_21_C241_n1168, B => 
                           mult_21_C241_n1088, CO => mult_21_C241_n680, S => 
                           mult_21_C241_n681);
   mult_21_C241_U1312 : ADHALFDL port map( A => mult_21_C241_n1206, B => 
                           mult_21_C241_n1090, CO => mult_21_C241_n732, S => 
                           mult_21_C241_n733);
   mult_21_C241_U1311 : INVD1 port map( A => mult_21_C241_n1537, Z => 
                           mult_21_C241_n1543);
   mult_21_C241_U1310 : ADHALFDL port map( A => mult_21_C241_n1306, B => 
                           mult_21_C241_n1094, CO => mult_21_C241_n788, S => 
                           mult_21_C241_n789);
   mult_21_C241_U1309 : ADHALFDL port map( A => mult_21_C241_n1333, B => 
                           mult_21_C241_n1363, CO => mult_21_C241_n784, S => 
                           mult_21_C241_n785);
   mult_21_C241_U1308 : INVD1 port map( A => mult_21_C241_n1536, Z => 
                           mult_21_C241_n1541);
   mult_21_C241_U1307 : ADHALFDL port map( A => mult_21_C241_n1252, B => 
                           mult_21_C241_n1092, CO => mult_21_C241_n768, S => 
                           mult_21_C241_n769);
   mult_21_C241_U1306 : INVD1 port map( A => mult_21_C241_n1534, Z => 
                           mult_21_C241_n1542);
   mult_21_C241_U1305 : ADHALFDL port map( A => mult_21_C241_n1331, B => 
                           mult_21_C241_n1361, CO => mult_21_C241_n774, S => 
                           mult_21_C241_n775);
   mult_21_C241_U1304 : INVD1 port map( A => mult_21_C241_n1535, Z => 
                           mult_21_C241_n1544);
   mult_21_C241_U1303 : NOR2D1 port map( A1 => mult_21_C241_n1537, A2 => 
                           mult_21_C241_n30, Z => mult_21_C241_n1093);
   mult_21_C241_U1302 : ADHALFDL port map( A => mult_21_C241_n1336, B => 
                           mult_21_C241_n1095, CO => mult_21_C241_n792, S => 
                           mult_21_C241_n793);
   mult_21_C241_U1301 : INVD1 port map( A => mult_21_C241_n1533, Z => 
                           mult_21_C241_n1545);
   mult_21_C241_U1300 : ADHALFDL port map( A => mult_21_C241_n1335, B => 
                           mult_21_C241_n1365, CO => mult_21_C241_n790, S => 
                           mult_21_C241_n791);
   mult_21_C241_U1299 : EXOR2D1 port map( A1 => mult_21_C241_n329, A2 => 
                           mult_21_C241_n344, Z => mult_21_C241_n155);
   mult_21_C241_U1298 : EXOR2D1 port map( A1 => mult_21_C241_n178, A2 => 
                           mult_21_C241_n155, Z => N3264);
   mult_21_C241_U1297 : NOR2D1 port map( A1 => mult_21_C241_n303, A2 => 
                           mult_21_C241_n305, Z => mult_21_C241_n302);
   mult_21_C241_U1296 : NAN2D1 port map( A1 => mult_21_C241_n1368, A2 => 
                           mult_21_C241_n1096, Z => mult_21_C241_n305);
   mult_21_C241_U1295 : NAN2D1 port map( A1 => mult_21_C241_n791, A2 => 
                           mult_21_C241_n792, Z => mult_21_C241_n296);
   mult_21_C241_U1294 : NAN2D1 port map( A1 => mult_21_C241_n783, A2 => 
                           mult_21_C241_n786, Z => mult_21_C241_n288);
   mult_21_C241_U1293 : NOR2D1 port map( A1 => mult_21_C241_n791, A2 => 
                           mult_21_C241_n792, Z => mult_21_C241_n295);
   mult_21_C241_U1292 : NOR2D1 port map( A1 => mult_21_C241_n783, A2 => 
                           mult_21_C241_n786, Z => mult_21_C241_n287);
   mult_21_C241_U1291 : NAN2D1 port map( A1 => mult_21_C241_n777, A2 => 
                           mult_21_C241_n782, Z => mult_21_C241_n284);
   mult_21_C241_U1290 : NAN2D1 port map( A1 => mult_21_C241_n793, A2 => 
                           mult_21_C241_n1366, Z => mult_21_C241_n301);
   mult_21_C241_U1289 : NAN2D1 port map( A1 => mult_21_C241_n787, A2 => 
                           mult_21_C241_n789, Z => mult_21_C241_n293);
   mult_21_C241_U1288 : NOR2D1 port map( A1 => mult_21_C241_n777, A2 => 
                           mult_21_C241_n782, Z => mult_21_C241_n283);
   mult_21_C241_U1287 : OR2D1 port map( A1 => mult_21_C241_n793, A2 => 
                           mult_21_C241_n1366, Z => mult_21_C241_n1532);
   mult_21_C241_U1286 : OR2D1 port map( A1 => mult_21_C241_n787, A2 => 
                           mult_21_C241_n789, Z => mult_21_C241_n1531);
   mult_21_C241_U1285 : NAN2D1 port map( A1 => mult_21_C241_n1532, A2 => 
                           mult_21_C241_n301, Z => mult_21_C241_n176);
   mult_21_C241_U1284 : INVD1 port map( A => mult_21_C241_n295, Z => 
                           mult_21_C241_n326);
   mult_21_C241_U1283 : NAN2D1 port map( A1 => mult_21_C241_n326, A2 => 
                           mult_21_C241_n296, Z => mult_21_C241_n175);
   mult_21_C241_U1282 : NAN2D1 port map( A1 => mult_21_C241_n1531, A2 => 
                           mult_21_C241_n293, Z => mult_21_C241_n174);
   mult_21_C241_U1281 : INVD1 port map( A => mult_21_C241_n287, Z => 
                           mult_21_C241_n324);
   mult_21_C241_U1280 : NAN2D1 port map( A1 => mult_21_C241_n324, A2 => 
                           mult_21_C241_n288, Z => mult_21_C241_n173);
   mult_21_C241_U1279 : INVD1 port map( A => mult_21_C241_n283, Z => 
                           mult_21_C241_n323);
   mult_21_C241_U1278 : NAN2D1 port map( A1 => mult_21_C241_n323, A2 => 
                           mult_21_C241_n284, Z => mult_21_C241_n172);
   mult_21_C241_U1277 : INVD1 port map( A => mult_21_C241_n280, Z => 
                           mult_21_C241_n322);
   mult_21_C241_U1276 : NAN2D1 port map( A1 => mult_21_C241_n322, A2 => 
                           mult_21_C241_n281, Z => mult_21_C241_n171);
   mult_21_C241_U1275 : NAN2D1 port map( A1 => mult_21_C241_n697, A2 => 
                           mult_21_C241_n710, Z => mult_21_C241_n240);
   mult_21_C241_U1274 : NAN2D1 port map( A1 => mult_21_C241_n711, A2 => 
                           mult_21_C241_n722, Z => mult_21_C241_n248);
   mult_21_C241_U1273 : NAN2D1 port map( A1 => mult_21_C241_n633, A2 => 
                           mult_21_C241_n650, Z => mult_21_C241_n221);
   mult_21_C241_U1272 : NOR2D1 port map( A1 => mult_21_C241_n697, A2 => 
                           mult_21_C241_n710, Z => mult_21_C241_n239);
   mult_21_C241_U1271 : NAN2D1 port map( A1 => mult_21_C241_n735, A2 => 
                           mult_21_C241_n744, Z => mult_21_C241_n259);
   mult_21_C241_U1270 : NOR2D1 port map( A1 => mult_21_C241_n615, A2 => 
                           mult_21_C241_n632, Z => mult_21_C241_n208);
   mult_21_C241_U1269 : NAN2D1 port map( A1 => mult_21_C241_n771, A2 => 
                           mult_21_C241_n776, Z => mult_21_C241_n281);
   mult_21_C241_U1268 : OR2D1 port map( A1 => mult_21_C241_n711, A2 => 
                           mult_21_C241_n722, Z => mult_21_C241_n1530);
   mult_21_C241_U1267 : NAN2D1 port map( A1 => mult_21_C241_n615, A2 => 
                           mult_21_C241_n632, Z => mult_21_C241_n209);
   mult_21_C241_U1266 : OR2D1 port map( A1 => mult_21_C241_n723, A2 => 
                           mult_21_C241_n734, Z => mult_21_C241_n1529);
   mult_21_C241_U1265 : NAN2D1 port map( A1 => mult_21_C241_n745, A2 => 
                           mult_21_C241_n754, Z => mult_21_C241_n262);
   mult_21_C241_U1264 : OR2D1 port map( A1 => mult_21_C241_n633, A2 => 
                           mult_21_C241_n650, Z => mult_21_C241_n1528);
   mult_21_C241_U1263 : NAN2D1 port map( A1 => mult_21_C241_n595, A2 => 
                           mult_21_C241_n614, Z => mult_21_C241_n206);
   mult_21_C241_U1262 : OR2D1 port map( A1 => mult_21_C241_n763, A2 => 
                           mult_21_C241_n770, Z => mult_21_C241_n1527);
   mult_21_C241_U1261 : NAN2D1 port map( A1 => mult_21_C241_n651, A2 => 
                           mult_21_C241_n666, Z => mult_21_C241_n226);
   mult_21_C241_U1260 : NAN2D1 port map( A1 => mult_21_C241_n723, A2 => 
                           mult_21_C241_n734, Z => mult_21_C241_n253);
   mult_21_C241_U1259 : NAN2D1 port map( A1 => mult_21_C241_n575, A2 => 
                           mult_21_C241_n594, Z => mult_21_C241_n199);
   mult_21_C241_U1258 : OR2D1 port map( A1 => mult_21_C241_n575, A2 => 
                           mult_21_C241_n594, Z => mult_21_C241_n1526);
   mult_21_C241_U1257 : NAN2D1 port map( A1 => mult_21_C241_n763, A2 => 
                           mult_21_C241_n770, Z => mult_21_C241_n275);
   mult_21_C241_U1256 : NOR2D1 port map( A1 => mult_21_C241_n735, A2 => 
                           mult_21_C241_n744, Z => mult_21_C241_n258);
   mult_21_C241_U1255 : NOR2D1 port map( A1 => mult_21_C241_n745, A2 => 
                           mult_21_C241_n754, Z => mult_21_C241_n261);
   mult_21_C241_U1254 : NOR2D1 port map( A1 => mult_21_C241_n771, A2 => 
                           mult_21_C241_n776, Z => mult_21_C241_n280);
   mult_21_C241_U1253 : OR2D1 port map( A1 => mult_21_C241_n595, A2 => 
                           mult_21_C241_n614, Z => mult_21_C241_n1525);
   mult_21_C241_U1252 : OA21M20D1 port map( A1 => mult_21_C241_n1532, A2 => 
                           mult_21_C241_n302, B => mult_21_C241_n301, Z => 
                           mult_21_C241_n297);
   mult_21_C241_U1251 : NOR2D1 port map( A1 => mult_21_C241_n651, A2 => 
                           mult_21_C241_n666, Z => mult_21_C241_n225);
   mult_21_C241_U1250 : OA21M20D1 port map( A1 => mult_21_C241_n1531, A2 => 
                           mult_21_C241_n294, B => mult_21_C241_n293, Z => 
                           mult_21_C241_n289);
   mult_21_C241_U1249 : NOR2D1 port map( A1 => mult_21_C241_n280, A2 => 
                           mult_21_C241_n283, Z => mult_21_C241_n278);
   mult_21_C241_U1248 : NAN2D1 port map( A1 => mult_21_C241_n755, A2 => 
                           mult_21_C241_n762, Z => mult_21_C241_n270);
   mult_21_C241_U1247 : OR2D1 port map( A1 => mult_21_C241_n755, A2 => 
                           mult_21_C241_n762, Z => mult_21_C241_n1524);
   mult_21_C241_U1246 : INVD1 port map( A => mult_21_C241_n286, Z => 
                           mult_21_C241_n285);
   mult_21_C241_U1245 : NAN2D1 port map( A1 => mult_21_C241_n1527, A2 => 
                           mult_21_C241_n275, Z => mult_21_C241_n170);
   mult_21_C241_U1244 : NAN2D1 port map( A1 => mult_21_C241_n1524, A2 => 
                           mult_21_C241_n270, Z => mult_21_C241_n169);
   mult_21_C241_U1243 : INVD1 port map( A => mult_21_C241_n277, Z => 
                           mult_21_C241_n276);
   mult_21_C241_U1242 : INVD1 port map( A => mult_21_C241_n261, Z => 
                           mult_21_C241_n319);
   mult_21_C241_U1241 : NAN2D1 port map( A1 => mult_21_C241_n319, A2 => 
                           mult_21_C241_n262, Z => mult_21_C241_n168);
   mult_21_C241_U1240 : INVD1 port map( A => mult_21_C241_n258, Z => 
                           mult_21_C241_n318);
   mult_21_C241_U1239 : NAN2D1 port map( A1 => mult_21_C241_n318, A2 => 
                           mult_21_C241_n259, Z => mult_21_C241_n167);
   mult_21_C241_U1238 : NAN2D1 port map( A1 => mult_21_C241_n1529, A2 => 
                           mult_21_C241_n253, Z => mult_21_C241_n166);
   mult_21_C241_U1237 : INVD1 port map( A => mult_21_C241_n239, Z => 
                           mult_21_C241_n315);
   mult_21_C241_U1236 : NAN2D1 port map( A1 => mult_21_C241_n315, A2 => 
                           mult_21_C241_n240, Z => mult_21_C241_n164);
   mult_21_C241_U1235 : NAN2D1 port map( A1 => mult_21_C241_n1530, A2 => 
                           mult_21_C241_n248, Z => mult_21_C241_n165);
   mult_21_C241_U1234 : INVD1 port map( A => mult_21_C241_n236, Z => 
                           mult_21_C241_n314);
   mult_21_C241_U1233 : NAN2D1 port map( A1 => mult_21_C241_n314, A2 => 
                           mult_21_C241_n237, Z => mult_21_C241_n163);
   mult_21_C241_U1232 : NAN2D1 port map( A1 => mult_21_C241_n1528, A2 => 
                           mult_21_C241_n221, Z => mult_21_C241_n160);
   mult_21_C241_U1231 : INVD1 port map( A => mult_21_C241_n225, Z => 
                           mult_21_C241_n312);
   mult_21_C241_U1230 : NAN2D1 port map( A1 => mult_21_C241_n312, A2 => 
                           mult_21_C241_n226, Z => mult_21_C241_n161);
   mult_21_C241_U1229 : NAN2D1 port map( A1 => mult_21_C241_n310, A2 => 
                           mult_21_C241_n209, Z => mult_21_C241_n159);
   mult_21_C241_U1228 : NAN2D1 port map( A1 => mult_21_C241_n1525, A2 => 
                           mult_21_C241_n206, Z => mult_21_C241_n158);
   mult_21_C241_U1227 : NAN2D1 port map( A1 => mult_21_C241_n1526, A2 => 
                           mult_21_C241_n199, Z => mult_21_C241_n157);
   mult_21_C241_U1226 : NAN2D1 port map( A1 => mult_21_C241_n1523, A2 => 
                           mult_21_C241_n194, Z => mult_21_C241_n156);
   mult_21_C241_U1225 : NAN2D1 port map( A1 => mult_21_C241_n683, A2 => 
                           mult_21_C241_n696, Z => mult_21_C241_n237);
   mult_21_C241_U1224 : NOR2D1 port map( A1 => mult_21_C241_n667, A2 => 
                           mult_21_C241_n682, Z => mult_21_C241_n230);
   mult_21_C241_U1223 : INVD1 port map( A => mult_21_C241_n208, Z => 
                           mult_21_C241_n310);
   mult_21_C241_U1222 : NAN2D1 port map( A1 => mult_21_C241_n553, A2 => 
                           mult_21_C241_n574, Z => mult_21_C241_n194);
   mult_21_C241_U1221 : NOR2D1 port map( A1 => mult_21_C241_n683, A2 => 
                           mult_21_C241_n696, Z => mult_21_C241_n236);
   mult_21_C241_U1220 : NAN2D1 port map( A1 => mult_21_C241_n1525, A2 => 
                           mult_21_C241_n310, Z => mult_21_C241_n201);
   mult_21_C241_U1219 : NOR2D1 port map( A1 => mult_21_C241_n225, A2 => 
                           mult_21_C241_n230, Z => mult_21_C241_n223);
   mult_21_C241_U1218 : NAN2D1 port map( A1 => mult_21_C241_n667, A2 => 
                           mult_21_C241_n682, Z => mult_21_C241_n231);
   mult_21_C241_U1217 : INVD1 port map( A => mult_21_C241_n253, Z => 
                           mult_21_C241_n251);
   mult_21_C241_U1216 : INVD1 port map( A => mult_21_C241_n199, Z => 
                           mult_21_C241_n197);
   mult_21_C241_U1215 : NAN2D1 port map( A1 => mult_21_C241_n1523, A2 => 
                           mult_21_C241_n1526, Z => mult_21_C241_n189);
   mult_21_C241_U1214 : OR2D1 port map( A1 => mult_21_C241_n553, A2 => 
                           mult_21_C241_n574, Z => mult_21_C241_n1523);
   mult_21_C241_U1213 : INVD1 port map( A => mult_21_C241_n275, Z => 
                           mult_21_C241_n273);
   mult_21_C241_U1212 : INVD1 port map( A => mult_21_C241_n206, Z => 
                           mult_21_C241_n204);
   mult_21_C241_U1211 : INVD1 port map( A => mult_21_C241_n209, Z => 
                           mult_21_C241_n211);
   mult_21_C241_U1210 : NOR2D1 port map( A1 => mult_21_C241_n189, A2 => 
                           mult_21_C241_n201, Z => mult_21_C241_n187);
   mult_21_C241_U1209 : NOR2D1 port map( A1 => mult_21_C241_n236, A2 => 
                           mult_21_C241_n239, Z => mult_21_C241_n234);
   mult_21_C241_U1208 : NOR2D1 port map( A1 => mult_21_C241_n258, A2 => 
                           mult_21_C241_n261, Z => mult_21_C241_n256);
   mult_21_C241_U1207 : INVD1 port map( A => mult_21_C241_n270, Z => 
                           mult_21_C241_n268);
   mult_21_C241_U1206 : NAN2D1 port map( A1 => mult_21_C241_n1524, A2 => 
                           mult_21_C241_n1527, Z => mult_21_C241_n265);
   mult_21_C241_U1205 : INVD1 port map( A => mult_21_C241_n248, Z => 
                           mult_21_C241_n246);
   mult_21_C241_U1204 : NAN2D1 port map( A1 => mult_21_C241_n1530, A2 => 
                           mult_21_C241_n1529, Z => mult_21_C241_n243);
   mult_21_C241_U1203 : INVD1 port map( A => mult_21_C241_n221, Z => 
                           mult_21_C241_n219);
   mult_21_C241_U1202 : NAN2D1 port map( A1 => mult_21_C241_n223, A2 => 
                           mult_21_C241_n1528, Z => mult_21_C241_n216);
   mult_21_C241_U1201 : INVD1 port map( A => mult_21_C241_n264, Z => 
                           mult_21_C241_n263);
   mult_21_C241_U1200 : INVD1 port map( A => mult_21_C241_n231, Z => 
                           mult_21_C241_n229);
   mult_21_C241_U1199 : INVD1 port map( A => mult_21_C241_n230, Z => 
                           mult_21_C241_n313);
   mult_21_C241_U1198 : INVD1 port map( A => mult_21_C241_n255, Z => 
                           mult_21_C241_n254);
   mult_21_C241_U1197 : INVD1 port map( A => mult_21_C241_n242, Z => 
                           mult_21_C241_n241);
   mult_21_C241_U1196 : NAN2D1 port map( A1 => mult_21_C241_n313, A2 => 
                           mult_21_C241_n231, Z => mult_21_C241_n162);
   mult_21_C241_U1195 : INVD1 port map( A => mult_21_C241_n233, Z => 
                           mult_21_C241_n232);
   mult_21_C241_U1194 : INVD1 port map( A => mult_21_C241_n215, Z => 
                           mult_21_C241_n214);
   mult_21_C241_U1193 : OA21M20D1 port map( A1 => mult_21_C241_n1523, A2 => 
                           mult_21_C241_n197, B => mult_21_C241_n194, Z => 
                           mult_21_C241_n190);
   mult_21_C241_U1192 : OR2D1 port map( A1 => mult_21_C241_n1368, A2 => 
                           mult_21_C241_n1096, Z => mult_21_C241_n1522);
   mult_21_C241_U1191 : AO21D1 port map( A1 => mult_21_C241_n215, A2 => 
                           mult_21_C241_n187, B => mult_21_C241_n188, Z => 
                           mult_21_C241_n1521);
   mult_21_C241_U1190 : AND2D1 port map( A1 => mult_21_C241_n1522, A2 => 
                           mult_21_C241_n305, Z => N3233);
   mult_21_C241_U1189 : OAI21D1 port map( A1 => N2920, A2 => N2921, B => 
                           mult_21_C241_n1077, Z => mult_21_C241_n1519);
   mult_21_C241_U1188 : OAI21D1 port map( A1 => N2916, A2 => N2917, B => 
                           mult_21_C241_n1079, Z => mult_21_C241_n1518);
   mult_21_C241_U1187 : OAI21D1 port map( A1 => N2914, A2 => N2915, B => 
                           mult_21_C241_n1080, Z => mult_21_C241_n1517);
   mult_21_C241_U1186 : ADHALFDL port map( A => mult_21_C241_n1278, B => 
                           mult_21_C241_n1093, CO => mult_21_C241_n780, S => 
                           mult_21_C241_n781);
   mult_21_C241_U1135 : EXNOR2D1 port map( A1 => N2936, A2 => N2937, Z => 
                           mult_21_C241_n93);
   mult_21_C241_U1131 : EXNOR2D1 port map( A1 => N2938, A2 => N2939, Z => 
                           mult_21_C241_n98);
   mult_21_C241_U1129 : OAI21D1 port map( A1 => N2938, A2 => N2939, B => 
                           mult_21_C241_n1068, Z => mult_21_C241_n94);
   mult_21_C241_U1127 : EXNOR2D1 port map( A1 => N2940, A2 => N2941, Z => 
                           mult_21_C241_n103);
   mult_21_C241_U1125 : OAI21D1 port map( A1 => N2940, A2 => N2941, B => 
                           mult_21_C241_n1067, Z => mult_21_C241_n99);
   mult_21_C241_U1123 : EXNOR2D1 port map( A1 => N2942, A2 => N2943, Z => 
                           mult_21_C241_n106);
   mult_21_C241_U1121 : OAI21D1 port map( A1 => N2942, A2 => N2943, B => 
                           mult_21_C241_n1066, Z => mult_21_C241_n104);
   mult_21_C241_U1120 : NAN2M1D1 port map( A1 => mult_21_C241_n8, A2 => 
                           mult_21_C241_n1548, Z => mult_21_C241_n1065);
   mult_21_C241_U1119 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1065, Z => 
                           mult_21_C241_n1368);
   mult_21_C241_U1118 : MUXB2DL port map( A0 => N3074, A1 => mult_21_C241_n1548
                           , SL => mult_21_C241_n8, Z => mult_21_C241_n1064);
   mult_21_C241_U1117 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1064, Z => 
                           mult_21_C241_n1367);
   mult_21_C241_U1116 : MUXB2DL port map( A0 => N3075, A1 => N3074, SL => 
                           mult_21_C241_n8, Z => mult_21_C241_n1063);
   mult_21_C241_U1115 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1063, Z => 
                           mult_21_C241_n1366);
   mult_21_C241_U1114 : MUXB2DL port map( A0 => N3076, A1 => mult_21_C241_n1546
                           , SL => mult_21_C241_n8, Z => mult_21_C241_n1062);
   mult_21_C241_U1113 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1062, Z => 
                           mult_21_C241_n1365);
   mult_21_C241_U1112 : MUXB2DL port map( A0 => N3077, A1 => N3076, SL => 
                           mult_21_C241_n8, Z => mult_21_C241_n1061);
   mult_21_C241_U1111 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1061, Z => 
                           mult_21_C241_n1364);
   mult_21_C241_U1110 : MUXB2DL port map( A0 => N3078, A1 => N3077, SL => 
                           mult_21_C241_n8, Z => mult_21_C241_n1060);
   mult_21_C241_U1109 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1060, Z => 
                           mult_21_C241_n1363);
   mult_21_C241_U1108 : MUXB2DL port map( A0 => N3079, A1 => N3078, SL => 
                           mult_21_C241_n8, Z => mult_21_C241_n1059);
   mult_21_C241_U1107 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1059, Z => 
                           mult_21_C241_n1362);
   mult_21_C241_U1106 : MUXB2DL port map( A0 => N3080, A1 => N3079, SL => 
                           mult_21_C241_n8, Z => mult_21_C241_n1058);
   mult_21_C241_U1105 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1058, Z => 
                           mult_21_C241_n1361);
   mult_21_C241_U1104 : MUXB2DL port map( A0 => N3081, A1 => N3080, SL => 
                           mult_21_C241_n8, Z => mult_21_C241_n1057);
   mult_21_C241_U1103 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1057, Z => 
                           mult_21_C241_n1360);
   mult_21_C241_U1102 : MUXB2DL port map( A0 => mult_21_C241_n1538, A1 => N3081
                           , SL => mult_21_C241_n8, Z => mult_21_C241_n1056);
   mult_21_C241_U1101 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1056, Z => 
                           mult_21_C241_n1359);
   mult_21_C241_U1100 : MUXB2DL port map( A0 => mult_21_C241_n1539, A1 => 
                           mult_21_C241_n1538, SL => mult_21_C241_n8, Z => 
                           mult_21_C241_n1055);
   mult_21_C241_U1099 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1055, Z => 
                           mult_21_C241_n1358);
   mult_21_C241_U1098 : MUXB2DL port map( A0 => mult_21_C241_n1540, A1 => 
                           mult_21_C241_n1539, SL => mult_21_C241_n8, Z => 
                           mult_21_C241_n1054);
   mult_21_C241_U1097 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1054, Z => 
                           mult_21_C241_n1357);
   mult_21_C241_U1096 : MUXB2DL port map( A0 => N3085, A1 => mult_21_C241_n1540
                           , SL => mult_21_C241_n8, Z => mult_21_C241_n1053);
   mult_21_C241_U1095 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1053, Z => 
                           mult_21_C241_n1356);
   mult_21_C241_U1094 : MUXB2DL port map( A0 => N3086, A1 => N3085, SL => 
                           mult_21_C241_n8, Z => mult_21_C241_n1052);
   mult_21_C241_U1093 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1052, Z => 
                           mult_21_C241_n1355);
   mult_21_C241_U1092 : MUXB2DL port map( A0 => N3087, A1 => N3086, SL => 
                           mult_21_C241_n8, Z => mult_21_C241_n1051);
   mult_21_C241_U1091 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1051, Z => 
                           mult_21_C241_n1354);
   mult_21_C241_U1090 : MUXB2DL port map( A0 => N3088, A1 => N3087, SL => 
                           mult_21_C241_n8, Z => mult_21_C241_n1050);
   mult_21_C241_U1089 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1050, Z => 
                           mult_21_C241_n1353);
   mult_21_C241_U1088 : MUXB2DL port map( A0 => N3089, A1 => N3088, SL => 
                           mult_21_C241_n8, Z => mult_21_C241_n1049);
   mult_21_C241_U1087 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1049, Z => 
                           mult_21_C241_n1352);
   mult_21_C241_U1086 : MUXB2DL port map( A0 => N3090, A1 => N3089, SL => 
                           mult_21_C241_n8, Z => mult_21_C241_n1048);
   mult_21_C241_U1085 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1048, Z => 
                           mult_21_C241_n1351);
   mult_21_C241_U1084 : MUXB2DL port map( A0 => N3091, A1 => N3090, SL => 
                           mult_21_C241_n8, Z => mult_21_C241_n1047);
   mult_21_C241_U1083 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1047, Z => 
                           mult_21_C241_n1350);
   mult_21_C241_U1082 : MUXB2DL port map( A0 => N3092, A1 => N3091, SL => 
                           mult_21_C241_n8, Z => mult_21_C241_n1046);
   mult_21_C241_U1081 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1046, Z => 
                           mult_21_C241_n1349);
   mult_21_C241_U1080 : MUXB2DL port map( A0 => N3093, A1 => N3092, SL => 
                           mult_21_C241_n8, Z => mult_21_C241_n1045);
   mult_21_C241_U1079 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1045, Z => 
                           mult_21_C241_n1348);
   mult_21_C241_U1078 : MUXB2DL port map( A0 => N3094, A1 => N3093, SL => 
                           mult_21_C241_n8, Z => mult_21_C241_n1044);
   mult_21_C241_U1077 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1044, Z => 
                           mult_21_C241_n1347);
   mult_21_C241_U1076 : MUXB2DL port map( A0 => N3095, A1 => N3094, SL => 
                           mult_21_C241_n8, Z => mult_21_C241_n1043);
   mult_21_C241_U1075 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1043, Z => 
                           mult_21_C241_n1346);
   mult_21_C241_U1074 : MUXB2DL port map( A0 => N3096, A1 => N3095, SL => 
                           mult_21_C241_n8, Z => mult_21_C241_n1042);
   mult_21_C241_U1073 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1042, Z => 
                           mult_21_C241_n1345);
   mult_21_C241_U1072 : MUXB2DL port map( A0 => N3097, A1 => N3096, SL => 
                           mult_21_C241_n8, Z => mult_21_C241_n1041);
   mult_21_C241_U1071 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1041, Z => 
                           mult_21_C241_n1344);
   mult_21_C241_U1070 : MUXB2DL port map( A0 => N3098, A1 => N3097, SL => 
                           mult_21_C241_n8, Z => mult_21_C241_n1040);
   mult_21_C241_U1069 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1040, Z => 
                           mult_21_C241_n1343);
   mult_21_C241_U1068 : MUXB2DL port map( A0 => N3099, A1 => N3098, SL => 
                           mult_21_C241_n8, Z => mult_21_C241_n1039);
   mult_21_C241_U1067 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1039, Z => 
                           mult_21_C241_n1342);
   mult_21_C241_U1066 : MUXB2DL port map( A0 => N3100, A1 => N3099, SL => 
                           mult_21_C241_n8, Z => mult_21_C241_n1038);
   mult_21_C241_U1065 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1038, Z => 
                           mult_21_C241_n1341);
   mult_21_C241_U1064 : MUXB2DL port map( A0 => N3101, A1 => N3100, SL => 
                           mult_21_C241_n8, Z => mult_21_C241_n1037);
   mult_21_C241_U1063 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1037, Z => 
                           mult_21_C241_n1340);
   mult_21_C241_U1062 : MUXB2DL port map( A0 => N3102, A1 => N3101, SL => 
                           mult_21_C241_n8, Z => mult_21_C241_n1036);
   mult_21_C241_U1061 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1036, Z => 
                           mult_21_C241_n1339);
   mult_21_C241_U1060 : MUXB2DL port map( A0 => N3103, A1 => N3102, SL => 
                           mult_21_C241_n8, Z => mult_21_C241_n1035);
   mult_21_C241_U1059 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1035, Z => 
                           mult_21_C241_n1338);
   mult_21_C241_U1058 : MUXB2DL port map( A0 => N3104, A1 => N3103, SL => 
                           mult_21_C241_n8, Z => mult_21_C241_n1034);
   mult_21_C241_U1057 : MUXB2DL port map( A0 => mult_21_C241_n3, A1 => 
                           mult_21_C241_n6, SL => mult_21_C241_n1034, Z => 
                           mult_21_C241_n1337);
   mult_21_C241_U1056 : NOR2M1D1 port map( A1 => mult_21_C241_n3, A2 => 
                           mult_21_C241_n6, Z => mult_21_C241_n1096);
   mult_21_C241_U1055 : NAN2M1D1 port map( A1 => mult_21_C241_n1545, A2 => 
                           N3073, Z => mult_21_C241_n1033);
   mult_21_C241_U1054 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1033, Z => 
                           mult_21_C241_n1336);
   mult_21_C241_U1053 : MUXB2DL port map( A0 => N3074, A1 => mult_21_C241_n1548
                           , SL => mult_21_C241_n1545, Z => mult_21_C241_n1032)
                           ;
   mult_21_C241_U1052 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1032, Z => 
                           mult_21_C241_n1335);
   mult_21_C241_U1051 : MUXB2DL port map( A0 => N3075, A1 => N3074, SL => 
                           mult_21_C241_n1545, Z => mult_21_C241_n1031);
   mult_21_C241_U1050 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1031, Z => 
                           mult_21_C241_n1334);
   mult_21_C241_U1049 : MUXB2DL port map( A0 => N3076, A1 => mult_21_C241_n1546
                           , SL => mult_21_C241_n1545, Z => mult_21_C241_n1030)
                           ;
   mult_21_C241_U1048 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1030, Z => 
                           mult_21_C241_n1333);
   mult_21_C241_U1047 : MUXB2DL port map( A0 => N3077, A1 => N3076, SL => 
                           mult_21_C241_n1545, Z => mult_21_C241_n1029);
   mult_21_C241_U1046 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1029, Z => 
                           mult_21_C241_n1332);
   mult_21_C241_U1045 : MUXB2DL port map( A0 => N3078, A1 => N3077, SL => 
                           mult_21_C241_n1545, Z => mult_21_C241_n1028);
   mult_21_C241_U1044 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1028, Z => 
                           mult_21_C241_n1331);
   mult_21_C241_U1043 : MUXB2DL port map( A0 => N3079, A1 => N3078, SL => 
                           mult_21_C241_n1545, Z => mult_21_C241_n1027);
   mult_21_C241_U1042 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1027, Z => 
                           mult_21_C241_n1330);
   mult_21_C241_U1041 : MUXB2DL port map( A0 => N3080, A1 => N3079, SL => 
                           mult_21_C241_n1545, Z => mult_21_C241_n1026);
   mult_21_C241_U1040 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1026, Z => 
                           mult_21_C241_n1329);
   mult_21_C241_U1039 : MUXB2DL port map( A0 => N3081, A1 => N3080, SL => 
                           mult_21_C241_n1545, Z => mult_21_C241_n1025);
   mult_21_C241_U1038 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1025, Z => 
                           mult_21_C241_n1328);
   mult_21_C241_U1037 : MUXB2DL port map( A0 => mult_21_C241_n1538, A1 => N3081
                           , SL => mult_21_C241_n1545, Z => mult_21_C241_n1024)
                           ;
   mult_21_C241_U1036 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1024, Z => 
                           mult_21_C241_n1327);
   mult_21_C241_U1035 : MUXB2DL port map( A0 => mult_21_C241_n1539, A1 => 
                           mult_21_C241_n1538, SL => mult_21_C241_n1545, Z => 
                           mult_21_C241_n1023);
   mult_21_C241_U1034 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1023, Z => 
                           mult_21_C241_n1326);
   mult_21_C241_U1033 : MUXB2DL port map( A0 => mult_21_C241_n1540, A1 => 
                           mult_21_C241_n1539, SL => mult_21_C241_n1545, Z => 
                           mult_21_C241_n1022);
   mult_21_C241_U1032 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1022, Z => 
                           mult_21_C241_n1325);
   mult_21_C241_U1031 : MUXB2DL port map( A0 => N3085, A1 => mult_21_C241_n1540
                           , SL => mult_21_C241_n1545, Z => mult_21_C241_n1021)
                           ;
   mult_21_C241_U1030 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1021, Z => 
                           mult_21_C241_n1324);
   mult_21_C241_U1029 : MUXB2DL port map( A0 => N3086, A1 => N3085, SL => 
                           mult_21_C241_n1545, Z => mult_21_C241_n1020);
   mult_21_C241_U1028 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1020, Z => 
                           mult_21_C241_n1323);
   mult_21_C241_U1027 : MUXB2DL port map( A0 => N3087, A1 => N3086, SL => 
                           mult_21_C241_n1545, Z => mult_21_C241_n1019);
   mult_21_C241_U1026 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1019, Z => 
                           mult_21_C241_n1322);
   mult_21_C241_U1025 : MUXB2DL port map( A0 => N3088, A1 => N3087, SL => 
                           mult_21_C241_n1545, Z => mult_21_C241_n1018);
   mult_21_C241_U1024 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1018, Z => 
                           mult_21_C241_n1321);
   mult_21_C241_U1023 : MUXB2DL port map( A0 => N3089, A1 => N3088, SL => 
                           mult_21_C241_n1545, Z => mult_21_C241_n1017);
   mult_21_C241_U1022 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1017, Z => 
                           mult_21_C241_n1320);
   mult_21_C241_U1021 : MUXB2DL port map( A0 => N3090, A1 => N3089, SL => 
                           mult_21_C241_n1545, Z => mult_21_C241_n1016);
   mult_21_C241_U1020 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1016, Z => 
                           mult_21_C241_n1319);
   mult_21_C241_U1019 : MUXB2DL port map( A0 => N3091, A1 => N3090, SL => 
                           mult_21_C241_n1545, Z => mult_21_C241_n1015);
   mult_21_C241_U1018 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1015, Z => 
                           mult_21_C241_n1318);
   mult_21_C241_U1017 : MUXB2DL port map( A0 => N3092, A1 => N3091, SL => 
                           mult_21_C241_n1545, Z => mult_21_C241_n1014);
   mult_21_C241_U1016 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1014, Z => 
                           mult_21_C241_n1317);
   mult_21_C241_U1015 : MUXB2DL port map( A0 => N3093, A1 => N3092, SL => 
                           mult_21_C241_n1545, Z => mult_21_C241_n1013);
   mult_21_C241_U1014 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1013, Z => 
                           mult_21_C241_n1316);
   mult_21_C241_U1013 : MUXB2DL port map( A0 => N3094, A1 => N3093, SL => 
                           mult_21_C241_n1545, Z => mult_21_C241_n1012);
   mult_21_C241_U1012 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1012, Z => 
                           mult_21_C241_n1315);
   mult_21_C241_U1011 : MUXB2DL port map( A0 => N3095, A1 => N3094, SL => 
                           mult_21_C241_n1545, Z => mult_21_C241_n1011);
   mult_21_C241_U1010 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1011, Z => 
                           mult_21_C241_n1314);
   mult_21_C241_U1009 : MUXB2DL port map( A0 => N3096, A1 => N3095, SL => 
                           mult_21_C241_n1545, Z => mult_21_C241_n1010);
   mult_21_C241_U1008 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1010, Z => 
                           mult_21_C241_n1313);
   mult_21_C241_U1007 : MUXB2DL port map( A0 => N3097, A1 => N3096, SL => 
                           mult_21_C241_n1545, Z => mult_21_C241_n1009);
   mult_21_C241_U1006 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1009, Z => 
                           mult_21_C241_n1312);
   mult_21_C241_U1005 : MUXB2DL port map( A0 => N3098, A1 => N3097, SL => 
                           mult_21_C241_n1545, Z => mult_21_C241_n1008);
   mult_21_C241_U1004 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1008, Z => 
                           mult_21_C241_n1311);
   mult_21_C241_U1003 : MUXB2DL port map( A0 => N3099, A1 => N3098, SL => 
                           mult_21_C241_n1545, Z => mult_21_C241_n1007);
   mult_21_C241_U1002 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1007, Z => 
                           mult_21_C241_n1310);
   mult_21_C241_U1001 : MUXB2DL port map( A0 => N3100, A1 => N3099, SL => 
                           mult_21_C241_n1545, Z => mult_21_C241_n1006);
   mult_21_C241_U1000 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1006, Z => 
                           mult_21_C241_n1309);
   mult_21_C241_U999 : MUXB2DL port map( A0 => N3101, A1 => N3100, SL => 
                           mult_21_C241_n1545, Z => mult_21_C241_n1005);
   mult_21_C241_U998 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1005, Z => 
                           mult_21_C241_n1308);
   mult_21_C241_U997 : MUXB2DL port map( A0 => N3102, A1 => N3101, SL => 
                           mult_21_C241_n1545, Z => mult_21_C241_n1004);
   mult_21_C241_U996 : MUXB2DL port map( A0 => mult_21_C241_n1517, A1 => 
                           mult_21_C241_n14, SL => mult_21_C241_n1004, Z => 
                           mult_21_C241_n1307);
   mult_21_C241_U995 : NOR2M1D1 port map( A1 => mult_21_C241_n1517, A2 => 
                           mult_21_C241_n14, Z => mult_21_C241_n1095);
   mult_21_C241_U994 : NAN2M1D1 port map( A1 => mult_21_C241_n1544, A2 => N3073
                           , Z => mult_21_C241_n1003);
   mult_21_C241_U993 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n1003, Z => 
                           mult_21_C241_n1306);
   mult_21_C241_U992 : MUXB2DL port map( A0 => N3074, A1 => mult_21_C241_n1548,
                           SL => mult_21_C241_n1544, Z => mult_21_C241_n1002);
   mult_21_C241_U991 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n1002, Z => 
                           mult_21_C241_n1305);
   mult_21_C241_U990 : MUXB2DL port map( A0 => N3075, A1 => N3074, SL => 
                           mult_21_C241_n1544, Z => mult_21_C241_n1001);
   mult_21_C241_U989 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n1001, Z => 
                           mult_21_C241_n1304);
   mult_21_C241_U988 : MUXB2DL port map( A0 => N3076, A1 => mult_21_C241_n1546,
                           SL => mult_21_C241_n1544, Z => mult_21_C241_n1000);
   mult_21_C241_U987 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n1000, Z => 
                           mult_21_C241_n1303);
   mult_21_C241_U986 : MUXB2DL port map( A0 => N3077, A1 => N3076, SL => 
                           mult_21_C241_n1544, Z => mult_21_C241_n999);
   mult_21_C241_U985 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n999, Z => 
                           mult_21_C241_n1302);
   mult_21_C241_U984 : MUXB2DL port map( A0 => N3078, A1 => N3077, SL => 
                           mult_21_C241_n1544, Z => mult_21_C241_n998);
   mult_21_C241_U983 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n998, Z => 
                           mult_21_C241_n1301);
   mult_21_C241_U982 : MUXB2DL port map( A0 => N3079, A1 => N3078, SL => 
                           mult_21_C241_n1544, Z => mult_21_C241_n997);
   mult_21_C241_U981 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n997, Z => 
                           mult_21_C241_n1300);
   mult_21_C241_U980 : MUXB2DL port map( A0 => N3080, A1 => N3079, SL => 
                           mult_21_C241_n1544, Z => mult_21_C241_n996);
   mult_21_C241_U979 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n996, Z => 
                           mult_21_C241_n1299);
   mult_21_C241_U978 : MUXB2DL port map( A0 => N3081, A1 => N3080, SL => 
                           mult_21_C241_n1544, Z => mult_21_C241_n995);
   mult_21_C241_U977 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n995, Z => 
                           mult_21_C241_n1298);
   mult_21_C241_U976 : MUXB2DL port map( A0 => mult_21_C241_n1538, A1 => N3081,
                           SL => mult_21_C241_n1544, Z => mult_21_C241_n994);
   mult_21_C241_U975 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n994, Z => 
                           mult_21_C241_n1297);
   mult_21_C241_U974 : MUXB2DL port map( A0 => mult_21_C241_n1539, A1 => 
                           mult_21_C241_n1538, SL => mult_21_C241_n1544, Z => 
                           mult_21_C241_n993);
   mult_21_C241_U973 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n993, Z => 
                           mult_21_C241_n1296);
   mult_21_C241_U972 : MUXB2DL port map( A0 => mult_21_C241_n1540, A1 => 
                           mult_21_C241_n1539, SL => mult_21_C241_n1544, Z => 
                           mult_21_C241_n992);
   mult_21_C241_U971 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n992, Z => 
                           mult_21_C241_n1295);
   mult_21_C241_U970 : MUXB2DL port map( A0 => N3085, A1 => mult_21_C241_n1540,
                           SL => mult_21_C241_n1544, Z => mult_21_C241_n991);
   mult_21_C241_U969 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n991, Z => 
                           mult_21_C241_n1294);
   mult_21_C241_U968 : MUXB2DL port map( A0 => N3086, A1 => N3085, SL => 
                           mult_21_C241_n1544, Z => mult_21_C241_n990);
   mult_21_C241_U967 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n990, Z => 
                           mult_21_C241_n1293);
   mult_21_C241_U966 : MUXB2DL port map( A0 => N3087, A1 => N3086, SL => 
                           mult_21_C241_n1544, Z => mult_21_C241_n989);
   mult_21_C241_U965 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n989, Z => 
                           mult_21_C241_n1292);
   mult_21_C241_U964 : MUXB2DL port map( A0 => N3088, A1 => N3087, SL => 
                           mult_21_C241_n1544, Z => mult_21_C241_n988);
   mult_21_C241_U963 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n988, Z => 
                           mult_21_C241_n1291);
   mult_21_C241_U962 : MUXB2DL port map( A0 => N3089, A1 => N3088, SL => 
                           mult_21_C241_n1544, Z => mult_21_C241_n987);
   mult_21_C241_U961 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n987, Z => 
                           mult_21_C241_n1290);
   mult_21_C241_U960 : MUXB2DL port map( A0 => N3090, A1 => N3089, SL => 
                           mult_21_C241_n1544, Z => mult_21_C241_n986);
   mult_21_C241_U959 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n986, Z => 
                           mult_21_C241_n1289);
   mult_21_C241_U958 : MUXB2DL port map( A0 => N3091, A1 => N3090, SL => 
                           mult_21_C241_n1544, Z => mult_21_C241_n985);
   mult_21_C241_U957 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n985, Z => 
                           mult_21_C241_n1288);
   mult_21_C241_U956 : MUXB2DL port map( A0 => N3092, A1 => N3091, SL => 
                           mult_21_C241_n1544, Z => mult_21_C241_n984);
   mult_21_C241_U955 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n984, Z => 
                           mult_21_C241_n1287);
   mult_21_C241_U954 : MUXB2DL port map( A0 => N3093, A1 => N3092, SL => 
                           mult_21_C241_n1544, Z => mult_21_C241_n983);
   mult_21_C241_U953 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n983, Z => 
                           mult_21_C241_n1286);
   mult_21_C241_U952 : MUXB2DL port map( A0 => N3094, A1 => N3093, SL => 
                           mult_21_C241_n1544, Z => mult_21_C241_n982);
   mult_21_C241_U951 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n982, Z => 
                           mult_21_C241_n1285);
   mult_21_C241_U950 : MUXB2DL port map( A0 => N3095, A1 => N3094, SL => 
                           mult_21_C241_n1544, Z => mult_21_C241_n981);
   mult_21_C241_U949 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n981, Z => 
                           mult_21_C241_n1284);
   mult_21_C241_U948 : MUXB2DL port map( A0 => N3096, A1 => N3095, SL => 
                           mult_21_C241_n1544, Z => mult_21_C241_n980);
   mult_21_C241_U947 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n980, Z => 
                           mult_21_C241_n1283);
   mult_21_C241_U946 : MUXB2DL port map( A0 => N3097, A1 => N3096, SL => 
                           mult_21_C241_n1544, Z => mult_21_C241_n979);
   mult_21_C241_U945 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n979, Z => 
                           mult_21_C241_n1282);
   mult_21_C241_U944 : MUXB2DL port map( A0 => N3098, A1 => N3097, SL => 
                           mult_21_C241_n1544, Z => mult_21_C241_n978);
   mult_21_C241_U943 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n978, Z => 
                           mult_21_C241_n1281);
   mult_21_C241_U942 : MUXB2DL port map( A0 => N3099, A1 => N3098, SL => 
                           mult_21_C241_n1544, Z => mult_21_C241_n977);
   mult_21_C241_U941 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n977, Z => 
                           mult_21_C241_n1280);
   mult_21_C241_U940 : MUXB2DL port map( A0 => N3100, A1 => N3099, SL => 
                           mult_21_C241_n1544, Z => mult_21_C241_n976);
   mult_21_C241_U939 : MUXB2DL port map( A0 => mult_21_C241_n1518, A1 => 
                           mult_21_C241_n22, SL => mult_21_C241_n976, Z => 
                           mult_21_C241_n1279);
   mult_21_C241_U938 : NOR2M1D1 port map( A1 => mult_21_C241_n1518, A2 => 
                           mult_21_C241_n22, Z => mult_21_C241_n1094);
   mult_21_C241_U937 : NAN2M1D1 port map( A1 => mult_21_C241_n1542, A2 => N3073
                           , Z => mult_21_C241_n975);
   mult_21_C241_U936 : MUXB2DL port map( A0 => mult_21_C241_n1543, A1 => 
                           mult_21_C241_n30, SL => mult_21_C241_n975, Z => 
                           mult_21_C241_n1278);
   mult_21_C241_U935 : MUXB2DL port map( A0 => N3074, A1 => N3073, SL => 
                           mult_21_C241_n1542, Z => mult_21_C241_n974);
   mult_21_C241_U934 : MUXB2DL port map( A0 => mult_21_C241_n1543, A1 => 
                           mult_21_C241_n30, SL => mult_21_C241_n974, Z => 
                           mult_21_C241_n1277);
   mult_21_C241_U933 : MUXB2DL port map( A0 => N3075, A1 => N3074, SL => 
                           mult_21_C241_n1542, Z => mult_21_C241_n973);
   mult_21_C241_U932 : MUXB2DL port map( A0 => mult_21_C241_n1543, A1 => 
                           mult_21_C241_n30, SL => mult_21_C241_n973, Z => 
                           mult_21_C241_n1276);
   mult_21_C241_U931 : MUXB2DL port map( A0 => N3076, A1 => N3075, SL => 
                           mult_21_C241_n1542, Z => mult_21_C241_n972);
   mult_21_C241_U930 : MUXB2DL port map( A0 => mult_21_C241_n1543, A1 => 
                           mult_21_C241_n30, SL => mult_21_C241_n972, Z => 
                           mult_21_C241_n1275);
   mult_21_C241_U929 : MUXB2DL port map( A0 => N3077, A1 => N3076, SL => 
                           mult_21_C241_n1542, Z => mult_21_C241_n971);
   mult_21_C241_U928 : MUXB2DL port map( A0 => mult_21_C241_n1543, A1 => 
                           mult_21_C241_n30, SL => mult_21_C241_n971, Z => 
                           mult_21_C241_n1274);
   mult_21_C241_U927 : MUXB2DL port map( A0 => N3078, A1 => N3077, SL => 
                           mult_21_C241_n1542, Z => mult_21_C241_n970);
   mult_21_C241_U926 : MUXB2DL port map( A0 => mult_21_C241_n1543, A1 => 
                           mult_21_C241_n30, SL => mult_21_C241_n970, Z => 
                           mult_21_C241_n1273);
   mult_21_C241_U925 : MUXB2DL port map( A0 => N3079, A1 => N3078, SL => 
                           mult_21_C241_n1542, Z => mult_21_C241_n969);
   mult_21_C241_U924 : MUXB2DL port map( A0 => mult_21_C241_n1543, A1 => 
                           mult_21_C241_n30, SL => mult_21_C241_n969, Z => 
                           mult_21_C241_n1272);
   mult_21_C241_U923 : MUXB2DL port map( A0 => N3080, A1 => N3079, SL => 
                           mult_21_C241_n1542, Z => mult_21_C241_n968);
   mult_21_C241_U922 : MUXB2DL port map( A0 => mult_21_C241_n1543, A1 => 
                           mult_21_C241_n30, SL => mult_21_C241_n968, Z => 
                           mult_21_C241_n1271);
   mult_21_C241_U921 : MUXB2DL port map( A0 => N3081, A1 => N3080, SL => 
                           mult_21_C241_n1542, Z => mult_21_C241_n967);
   mult_21_C241_U920 : MUXB2DL port map( A0 => mult_21_C241_n1543, A1 => 
                           mult_21_C241_n30, SL => mult_21_C241_n967, Z => 
                           mult_21_C241_n1270);
   mult_21_C241_U919 : MUXB2DL port map( A0 => mult_21_C241_n1538, A1 => N3081,
                           SL => mult_21_C241_n1542, Z => mult_21_C241_n966);
   mult_21_C241_U918 : MUXB2DL port map( A0 => mult_21_C241_n1543, A1 => 
                           mult_21_C241_n30, SL => mult_21_C241_n966, Z => 
                           mult_21_C241_n1269);
   mult_21_C241_U917 : MUXB2DL port map( A0 => mult_21_C241_n1539, A1 => 
                           mult_21_C241_n1538, SL => mult_21_C241_n1542, Z => 
                           mult_21_C241_n965);
   mult_21_C241_U916 : MUXB2DL port map( A0 => mult_21_C241_n1543, A1 => 
                           mult_21_C241_n30, SL => mult_21_C241_n965, Z => 
                           mult_21_C241_n1268);
   mult_21_C241_U915 : MUXB2DL port map( A0 => mult_21_C241_n1540, A1 => 
                           mult_21_C241_n1539, SL => mult_21_C241_n1542, Z => 
                           mult_21_C241_n964);
   mult_21_C241_U914 : MUXB2DL port map( A0 => mult_21_C241_n1543, A1 => 
                           mult_21_C241_n30, SL => mult_21_C241_n964, Z => 
                           mult_21_C241_n1267);
   mult_21_C241_U913 : MUXB2DL port map( A0 => N3085, A1 => mult_21_C241_n1540,
                           SL => mult_21_C241_n1542, Z => mult_21_C241_n963);
   mult_21_C241_U912 : MUXB2DL port map( A0 => mult_21_C241_n1543, A1 => 
                           mult_21_C241_n30, SL => mult_21_C241_n963, Z => 
                           mult_21_C241_n1266);
   mult_21_C241_U911 : MUXB2DL port map( A0 => N3086, A1 => N3085, SL => 
                           mult_21_C241_n1542, Z => mult_21_C241_n962);
   mult_21_C241_U910 : MUXB2DL port map( A0 => mult_21_C241_n1543, A1 => 
                           mult_21_C241_n30, SL => mult_21_C241_n962, Z => 
                           mult_21_C241_n1265);
   mult_21_C241_U909 : MUXB2DL port map( A0 => N3087, A1 => N3086, SL => 
                           mult_21_C241_n1542, Z => mult_21_C241_n961);
   mult_21_C241_U908 : MUXB2DL port map( A0 => mult_21_C241_n1543, A1 => 
                           mult_21_C241_n30, SL => mult_21_C241_n961, Z => 
                           mult_21_C241_n1264);
   mult_21_C241_U907 : MUXB2DL port map( A0 => N3088, A1 => N3087, SL => 
                           mult_21_C241_n1542, Z => mult_21_C241_n960);
   mult_21_C241_U906 : MUXB2DL port map( A0 => mult_21_C241_n1543, A1 => 
                           mult_21_C241_n30, SL => mult_21_C241_n960, Z => 
                           mult_21_C241_n1263);
   mult_21_C241_U905 : MUXB2DL port map( A0 => N3089, A1 => N3088, SL => 
                           mult_21_C241_n1542, Z => mult_21_C241_n959);
   mult_21_C241_U904 : MUXB2DL port map( A0 => mult_21_C241_n1543, A1 => 
                           mult_21_C241_n30, SL => mult_21_C241_n959, Z => 
                           mult_21_C241_n1262);
   mult_21_C241_U903 : MUXB2DL port map( A0 => N3090, A1 => N3089, SL => 
                           mult_21_C241_n1542, Z => mult_21_C241_n958);
   mult_21_C241_U902 : MUXB2DL port map( A0 => mult_21_C241_n1543, A1 => 
                           mult_21_C241_n30, SL => mult_21_C241_n958, Z => 
                           mult_21_C241_n1261);
   mult_21_C241_U901 : MUXB2DL port map( A0 => N3091, A1 => N3090, SL => 
                           mult_21_C241_n1542, Z => mult_21_C241_n957);
   mult_21_C241_U900 : MUXB2DL port map( A0 => mult_21_C241_n1543, A1 => 
                           mult_21_C241_n30, SL => mult_21_C241_n957, Z => 
                           mult_21_C241_n1260);
   mult_21_C241_U899 : MUXB2DL port map( A0 => N3092, A1 => N3091, SL => 
                           mult_21_C241_n1542, Z => mult_21_C241_n956);
   mult_21_C241_U898 : MUXB2DL port map( A0 => mult_21_C241_n1543, A1 => 
                           mult_21_C241_n30, SL => mult_21_C241_n956, Z => 
                           mult_21_C241_n1259);
   mult_21_C241_U897 : MUXB2DL port map( A0 => N3093, A1 => N3092, SL => 
                           mult_21_C241_n1542, Z => mult_21_C241_n955);
   mult_21_C241_U896 : MUXB2DL port map( A0 => mult_21_C241_n1543, A1 => 
                           mult_21_C241_n30, SL => mult_21_C241_n955, Z => 
                           mult_21_C241_n1258);
   mult_21_C241_U895 : MUXB2DL port map( A0 => N3094, A1 => N3093, SL => 
                           mult_21_C241_n1542, Z => mult_21_C241_n954);
   mult_21_C241_U894 : MUXB2DL port map( A0 => mult_21_C241_n1543, A1 => 
                           mult_21_C241_n30, SL => mult_21_C241_n954, Z => 
                           mult_21_C241_n1257);
   mult_21_C241_U893 : MUXB2DL port map( A0 => N3095, A1 => N3094, SL => 
                           mult_21_C241_n1542, Z => mult_21_C241_n953);
   mult_21_C241_U892 : MUXB2DL port map( A0 => mult_21_C241_n1543, A1 => 
                           mult_21_C241_n30, SL => mult_21_C241_n953, Z => 
                           mult_21_C241_n1256);
   mult_21_C241_U891 : MUXB2DL port map( A0 => N3096, A1 => N3095, SL => 
                           mult_21_C241_n1542, Z => mult_21_C241_n952);
   mult_21_C241_U890 : MUXB2DL port map( A0 => mult_21_C241_n1543, A1 => 
                           mult_21_C241_n30, SL => mult_21_C241_n952, Z => 
                           mult_21_C241_n1255);
   mult_21_C241_U889 : MUXB2DL port map( A0 => N3097, A1 => N3096, SL => 
                           mult_21_C241_n1542, Z => mult_21_C241_n951);
   mult_21_C241_U888 : MUXB2DL port map( A0 => mult_21_C241_n1543, A1 => 
                           mult_21_C241_n30, SL => mult_21_C241_n951, Z => 
                           mult_21_C241_n1254);
   mult_21_C241_U887 : MUXB2DL port map( A0 => N3098, A1 => N3097, SL => 
                           mult_21_C241_n1542, Z => mult_21_C241_n950);
   mult_21_C241_U886 : MUXB2DL port map( A0 => mult_21_C241_n1543, A1 => 
                           mult_21_C241_n30, SL => mult_21_C241_n950, Z => 
                           mult_21_C241_n1253);
   mult_21_C241_U884 : NAN2M1D1 port map( A1 => mult_21_C241_n1541, A2 => N3073
                           , Z => mult_21_C241_n949);
   mult_21_C241_U883 : MUXB2DL port map( A0 => mult_21_C241_n1519, A1 => 
                           mult_21_C241_n38, SL => mult_21_C241_n949, Z => 
                           mult_21_C241_n1252);
   mult_21_C241_U882 : MUXB2DL port map( A0 => N3074, A1 => N3073, SL => 
                           mult_21_C241_n1541, Z => mult_21_C241_n948);
   mult_21_C241_U881 : MUXB2DL port map( A0 => mult_21_C241_n1519, A1 => 
                           mult_21_C241_n38, SL => mult_21_C241_n948, Z => 
                           mult_21_C241_n1251);
   mult_21_C241_U880 : MUXB2DL port map( A0 => N3075, A1 => N3074, SL => 
                           mult_21_C241_n1541, Z => mult_21_C241_n947);
   mult_21_C241_U879 : MUXB2DL port map( A0 => mult_21_C241_n1519, A1 => 
                           mult_21_C241_n38, SL => mult_21_C241_n947, Z => 
                           mult_21_C241_n1250);
   mult_21_C241_U878 : MUXB2DL port map( A0 => N3076, A1 => N3075, SL => 
                           mult_21_C241_n1541, Z => mult_21_C241_n946);
   mult_21_C241_U877 : MUXB2DL port map( A0 => mult_21_C241_n1519, A1 => 
                           mult_21_C241_n38, SL => mult_21_C241_n946, Z => 
                           mult_21_C241_n1249);
   mult_21_C241_U876 : MUXB2DL port map( A0 => N3077, A1 => N3076, SL => 
                           mult_21_C241_n1541, Z => mult_21_C241_n945);
   mult_21_C241_U875 : MUXB2DL port map( A0 => mult_21_C241_n1519, A1 => 
                           mult_21_C241_n38, SL => mult_21_C241_n945, Z => 
                           mult_21_C241_n1248);
   mult_21_C241_U874 : MUXB2DL port map( A0 => N3078, A1 => N3077, SL => 
                           mult_21_C241_n1541, Z => mult_21_C241_n944);
   mult_21_C241_U873 : MUXB2DL port map( A0 => mult_21_C241_n1519, A1 => 
                           mult_21_C241_n38, SL => mult_21_C241_n944, Z => 
                           mult_21_C241_n1247);
   mult_21_C241_U872 : MUXB2DL port map( A0 => N3079, A1 => N3078, SL => 
                           mult_21_C241_n1541, Z => mult_21_C241_n943);
   mult_21_C241_U871 : MUXB2DL port map( A0 => mult_21_C241_n1519, A1 => 
                           mult_21_C241_n38, SL => mult_21_C241_n943, Z => 
                           mult_21_C241_n1246);
   mult_21_C241_U870 : MUXB2DL port map( A0 => N3080, A1 => N3079, SL => 
                           mult_21_C241_n1541, Z => mult_21_C241_n942);
   mult_21_C241_U869 : MUXB2DL port map( A0 => mult_21_C241_n1519, A1 => 
                           mult_21_C241_n38, SL => mult_21_C241_n942, Z => 
                           mult_21_C241_n1245);
   mult_21_C241_U868 : MUXB2DL port map( A0 => N3081, A1 => N3080, SL => 
                           mult_21_C241_n1541, Z => mult_21_C241_n941);
   mult_21_C241_U867 : MUXB2DL port map( A0 => mult_21_C241_n1519, A1 => 
                           mult_21_C241_n38, SL => mult_21_C241_n941, Z => 
                           mult_21_C241_n1244);
   mult_21_C241_U866 : MUXB2DL port map( A0 => mult_21_C241_n1538, A1 => N3081,
                           SL => mult_21_C241_n1541, Z => mult_21_C241_n940);
   mult_21_C241_U865 : MUXB2DL port map( A0 => mult_21_C241_n1519, A1 => 
                           mult_21_C241_n38, SL => mult_21_C241_n940, Z => 
                           mult_21_C241_n1243);
   mult_21_C241_U864 : MUXB2DL port map( A0 => mult_21_C241_n1539, A1 => 
                           mult_21_C241_n1538, SL => mult_21_C241_n1541, Z => 
                           mult_21_C241_n939);
   mult_21_C241_U863 : MUXB2DL port map( A0 => mult_21_C241_n1519, A1 => 
                           mult_21_C241_n38, SL => mult_21_C241_n939, Z => 
                           mult_21_C241_n1242);
   mult_21_C241_U862 : MUXB2DL port map( A0 => mult_21_C241_n1540, A1 => 
                           mult_21_C241_n1539, SL => mult_21_C241_n1541, Z => 
                           mult_21_C241_n938);
   mult_21_C241_U861 : MUXB2DL port map( A0 => mult_21_C241_n1519, A1 => 
                           mult_21_C241_n38, SL => mult_21_C241_n938, Z => 
                           mult_21_C241_n1241);
   mult_21_C241_U860 : MUXB2DL port map( A0 => N3085, A1 => mult_21_C241_n1540,
                           SL => mult_21_C241_n1541, Z => mult_21_C241_n937);
   mult_21_C241_U859 : MUXB2DL port map( A0 => mult_21_C241_n1519, A1 => 
                           mult_21_C241_n38, SL => mult_21_C241_n937, Z => 
                           mult_21_C241_n1240);
   mult_21_C241_U858 : MUXB2DL port map( A0 => N3086, A1 => N3085, SL => 
                           mult_21_C241_n1541, Z => mult_21_C241_n936);
   mult_21_C241_U857 : MUXB2DL port map( A0 => mult_21_C241_n1519, A1 => 
                           mult_21_C241_n38, SL => mult_21_C241_n936, Z => 
                           mult_21_C241_n1239);
   mult_21_C241_U856 : MUXB2DL port map( A0 => N3087, A1 => N3086, SL => 
                           mult_21_C241_n1541, Z => mult_21_C241_n935);
   mult_21_C241_U855 : MUXB2DL port map( A0 => mult_21_C241_n1519, A1 => 
                           mult_21_C241_n38, SL => mult_21_C241_n935, Z => 
                           mult_21_C241_n1238);
   mult_21_C241_U854 : MUXB2DL port map( A0 => N3088, A1 => N3087, SL => 
                           mult_21_C241_n1541, Z => mult_21_C241_n934);
   mult_21_C241_U853 : MUXB2DL port map( A0 => mult_21_C241_n1519, A1 => 
                           mult_21_C241_n38, SL => mult_21_C241_n934, Z => 
                           mult_21_C241_n1237);
   mult_21_C241_U852 : MUXB2DL port map( A0 => N3089, A1 => N3088, SL => 
                           mult_21_C241_n1541, Z => mult_21_C241_n933);
   mult_21_C241_U851 : MUXB2DL port map( A0 => mult_21_C241_n1519, A1 => 
                           mult_21_C241_n38, SL => mult_21_C241_n933, Z => 
                           mult_21_C241_n1236);
   mult_21_C241_U850 : MUXB2DL port map( A0 => N3090, A1 => N3089, SL => 
                           mult_21_C241_n1541, Z => mult_21_C241_n932);
   mult_21_C241_U849 : MUXB2DL port map( A0 => mult_21_C241_n1519, A1 => 
                           mult_21_C241_n38, SL => mult_21_C241_n932, Z => 
                           mult_21_C241_n1235);
   mult_21_C241_U848 : MUXB2DL port map( A0 => N3091, A1 => N3090, SL => 
                           mult_21_C241_n1541, Z => mult_21_C241_n931);
   mult_21_C241_U847 : MUXB2DL port map( A0 => mult_21_C241_n1519, A1 => 
                           mult_21_C241_n38, SL => mult_21_C241_n931, Z => 
                           mult_21_C241_n1234);
   mult_21_C241_U846 : MUXB2DL port map( A0 => N3092, A1 => N3091, SL => 
                           mult_21_C241_n1541, Z => mult_21_C241_n930);
   mult_21_C241_U845 : MUXB2DL port map( A0 => mult_21_C241_n1519, A1 => 
                           mult_21_C241_n38, SL => mult_21_C241_n930, Z => 
                           mult_21_C241_n1233);
   mult_21_C241_U844 : MUXB2DL port map( A0 => N3093, A1 => N3092, SL => 
                           mult_21_C241_n1541, Z => mult_21_C241_n929);
   mult_21_C241_U843 : MUXB2DL port map( A0 => mult_21_C241_n1519, A1 => 
                           mult_21_C241_n38, SL => mult_21_C241_n929, Z => 
                           mult_21_C241_n1232);
   mult_21_C241_U842 : MUXB2DL port map( A0 => N3094, A1 => N3093, SL => 
                           mult_21_C241_n1541, Z => mult_21_C241_n928);
   mult_21_C241_U841 : MUXB2DL port map( A0 => mult_21_C241_n1519, A1 => 
                           mult_21_C241_n38, SL => mult_21_C241_n928, Z => 
                           mult_21_C241_n1231);
   mult_21_C241_U840 : MUXB2DL port map( A0 => N3095, A1 => N3094, SL => 
                           mult_21_C241_n1541, Z => mult_21_C241_n927);
   mult_21_C241_U839 : MUXB2DL port map( A0 => mult_21_C241_n1519, A1 => 
                           mult_21_C241_n38, SL => mult_21_C241_n927, Z => 
                           mult_21_C241_n1230);
   mult_21_C241_U838 : MUXB2DL port map( A0 => N3096, A1 => N3095, SL => 
                           mult_21_C241_n1541, Z => mult_21_C241_n926);
   mult_21_C241_U837 : MUXB2DL port map( A0 => mult_21_C241_n1519, A1 => 
                           mult_21_C241_n38, SL => mult_21_C241_n926, Z => 
                           mult_21_C241_n1229);
   mult_21_C241_U836 : NOR2M1D1 port map( A1 => mult_21_C241_n1519, A2 => 
                           mult_21_C241_n38, Z => mult_21_C241_n1092);
   mult_21_C241_U835 : NAN2M1D1 port map( A1 => mult_21_C241_n48, A2 => N3073, 
                           Z => mult_21_C241_n925);
   mult_21_C241_U834 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n45, SL => mult_21_C241_n925, Z => 
                           mult_21_C241_n1228);
   mult_21_C241_U833 : MUXB2DL port map( A0 => N3074, A1 => N3073, SL => 
                           mult_21_C241_n48, Z => mult_21_C241_n924);
   mult_21_C241_U832 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n45, SL => mult_21_C241_n924, Z => 
                           mult_21_C241_n1227);
   mult_21_C241_U831 : MUXB2DL port map( A0 => N3075, A1 => N3074, SL => 
                           mult_21_C241_n48, Z => mult_21_C241_n923);
   mult_21_C241_U830 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n45, SL => mult_21_C241_n923, Z => 
                           mult_21_C241_n1226);
   mult_21_C241_U829 : MUXB2DL port map( A0 => N3076, A1 => N3075, SL => 
                           mult_21_C241_n48, Z => mult_21_C241_n922);
   mult_21_C241_U828 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n45, SL => mult_21_C241_n922, Z => 
                           mult_21_C241_n1225);
   mult_21_C241_U827 : MUXB2DL port map( A0 => N3077, A1 => N3076, SL => 
                           mult_21_C241_n48, Z => mult_21_C241_n921);
   mult_21_C241_U826 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n45, SL => mult_21_C241_n921, Z => 
                           mult_21_C241_n1224);
   mult_21_C241_U825 : MUXB2DL port map( A0 => N3078, A1 => N3077, SL => 
                           mult_21_C241_n48, Z => mult_21_C241_n920);
   mult_21_C241_U824 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n45, SL => mult_21_C241_n920, Z => 
                           mult_21_C241_n1223);
   mult_21_C241_U823 : MUXB2DL port map( A0 => N3079, A1 => N3078, SL => 
                           mult_21_C241_n48, Z => mult_21_C241_n919);
   mult_21_C241_U822 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n45, SL => mult_21_C241_n919, Z => 
                           mult_21_C241_n1222);
   mult_21_C241_U821 : MUXB2DL port map( A0 => N3080, A1 => N3079, SL => 
                           mult_21_C241_n48, Z => mult_21_C241_n918);
   mult_21_C241_U820 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n45, SL => mult_21_C241_n918, Z => 
                           mult_21_C241_n1221);
   mult_21_C241_U819 : MUXB2DL port map( A0 => N3081, A1 => N3080, SL => 
                           mult_21_C241_n48, Z => mult_21_C241_n917);
   mult_21_C241_U818 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n45, SL => mult_21_C241_n917, Z => 
                           mult_21_C241_n1220);
   mult_21_C241_U817 : MUXB2DL port map( A0 => mult_21_C241_n1538, A1 => N3081,
                           SL => mult_21_C241_n48, Z => mult_21_C241_n916);
   mult_21_C241_U816 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n45, SL => mult_21_C241_n916, Z => 
                           mult_21_C241_n1219);
   mult_21_C241_U815 : MUXB2DL port map( A0 => mult_21_C241_n1539, A1 => 
                           mult_21_C241_n1538, SL => mult_21_C241_n48, Z => 
                           mult_21_C241_n915);
   mult_21_C241_U814 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n45, SL => mult_21_C241_n915, Z => 
                           mult_21_C241_n1218);
   mult_21_C241_U813 : MUXB2DL port map( A0 => mult_21_C241_n1540, A1 => 
                           mult_21_C241_n1539, SL => mult_21_C241_n48, Z => 
                           mult_21_C241_n914);
   mult_21_C241_U812 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n45, SL => mult_21_C241_n914, Z => 
                           mult_21_C241_n1217);
   mult_21_C241_U811 : MUXB2DL port map( A0 => N3085, A1 => mult_21_C241_n1540,
                           SL => mult_21_C241_n48, Z => mult_21_C241_n913);
   mult_21_C241_U810 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n45, SL => mult_21_C241_n913, Z => 
                           mult_21_C241_n1216);
   mult_21_C241_U809 : MUXB2DL port map( A0 => N3086, A1 => N3085, SL => 
                           mult_21_C241_n48, Z => mult_21_C241_n912);
   mult_21_C241_U808 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n45, SL => mult_21_C241_n912, Z => 
                           mult_21_C241_n1215);
   mult_21_C241_U807 : MUXB2DL port map( A0 => N3087, A1 => N3086, SL => 
                           mult_21_C241_n48, Z => mult_21_C241_n911);
   mult_21_C241_U806 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n45, SL => mult_21_C241_n911, Z => 
                           mult_21_C241_n1214);
   mult_21_C241_U805 : MUXB2DL port map( A0 => N3088, A1 => N3087, SL => 
                           mult_21_C241_n48, Z => mult_21_C241_n910);
   mult_21_C241_U804 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n45, SL => mult_21_C241_n910, Z => 
                           mult_21_C241_n1213);
   mult_21_C241_U803 : MUXB2DL port map( A0 => N3089, A1 => N3088, SL => 
                           mult_21_C241_n48, Z => mult_21_C241_n909);
   mult_21_C241_U802 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n45, SL => mult_21_C241_n909, Z => 
                           mult_21_C241_n1212);
   mult_21_C241_U801 : MUXB2DL port map( A0 => N3090, A1 => N3089, SL => 
                           mult_21_C241_n48, Z => mult_21_C241_n908);
   mult_21_C241_U800 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n45, SL => mult_21_C241_n908, Z => 
                           mult_21_C241_n1211);
   mult_21_C241_U799 : MUXB2DL port map( A0 => N3091, A1 => N3090, SL => 
                           mult_21_C241_n48, Z => mult_21_C241_n907);
   mult_21_C241_U798 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n45, SL => mult_21_C241_n907, Z => 
                           mult_21_C241_n1210);
   mult_21_C241_U797 : MUXB2DL port map( A0 => N3092, A1 => N3091, SL => 
                           mult_21_C241_n48, Z => mult_21_C241_n906);
   mult_21_C241_U796 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n45, SL => mult_21_C241_n906, Z => 
                           mult_21_C241_n1209);
   mult_21_C241_U795 : MUXB2DL port map( A0 => N3093, A1 => N3092, SL => 
                           mult_21_C241_n48, Z => mult_21_C241_n905);
   mult_21_C241_U794 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n45, SL => mult_21_C241_n905, Z => 
                           mult_21_C241_n1208);
   mult_21_C241_U793 : MUXB2DL port map( A0 => N3094, A1 => N3093, SL => 
                           mult_21_C241_n48, Z => mult_21_C241_n904);
   mult_21_C241_U792 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n45, SL => mult_21_C241_n904, Z => 
                           mult_21_C241_n1207);
   mult_21_C241_U791 : NOR2M1D1 port map( A1 => mult_21_C241_n42, A2 => 
                           mult_21_C241_n45, Z => mult_21_C241_n1091);
   mult_21_C241_U790 : NAN2M1D1 port map( A1 => mult_21_C241_n56, A2 => 
                           mult_21_C241_n1548, Z => mult_21_C241_n903);
   mult_21_C241_U789 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n53, SL => mult_21_C241_n903, Z => 
                           mult_21_C241_n1206);
   mult_21_C241_U788 : MUXB2DL port map( A0 => N3074, A1 => N3073, SL => 
                           mult_21_C241_n56, Z => mult_21_C241_n902);
   mult_21_C241_U787 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n53, SL => mult_21_C241_n902, Z => 
                           mult_21_C241_n1205);
   mult_21_C241_U786 : MUXB2DL port map( A0 => N3075, A1 => N3074, SL => 
                           mult_21_C241_n56, Z => mult_21_C241_n901);
   mult_21_C241_U785 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n53, SL => mult_21_C241_n901, Z => 
                           mult_21_C241_n1204);
   mult_21_C241_U784 : MUXB2DL port map( A0 => N3076, A1 => mult_21_C241_n1546,
                           SL => mult_21_C241_n56, Z => mult_21_C241_n900);
   mult_21_C241_U783 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n53, SL => mult_21_C241_n900, Z => 
                           mult_21_C241_n1203);
   mult_21_C241_U782 : MUXB2DL port map( A0 => N3077, A1 => N3076, SL => 
                           mult_21_C241_n56, Z => mult_21_C241_n899);
   mult_21_C241_U781 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n53, SL => mult_21_C241_n899, Z => 
                           mult_21_C241_n1202);
   mult_21_C241_U780 : MUXB2DL port map( A0 => N3078, A1 => N3077, SL => 
                           mult_21_C241_n56, Z => mult_21_C241_n898);
   mult_21_C241_U779 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n53, SL => mult_21_C241_n898, Z => 
                           mult_21_C241_n1201);
   mult_21_C241_U778 : MUXB2DL port map( A0 => N3079, A1 => N3078, SL => 
                           mult_21_C241_n56, Z => mult_21_C241_n897);
   mult_21_C241_U777 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n53, SL => mult_21_C241_n897, Z => 
                           mult_21_C241_n1200);
   mult_21_C241_U776 : MUXB2DL port map( A0 => N3080, A1 => N3079, SL => 
                           mult_21_C241_n56, Z => mult_21_C241_n896);
   mult_21_C241_U775 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n53, SL => mult_21_C241_n896, Z => 
                           mult_21_C241_n1199);
   mult_21_C241_U774 : MUXB2DL port map( A0 => N3081, A1 => N3080, SL => 
                           mult_21_C241_n56, Z => mult_21_C241_n895);
   mult_21_C241_U773 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n53, SL => mult_21_C241_n895, Z => 
                           mult_21_C241_n1198);
   mult_21_C241_U772 : MUXB2DL port map( A0 => mult_21_C241_n1538, A1 => N3081,
                           SL => mult_21_C241_n56, Z => mult_21_C241_n894);
   mult_21_C241_U771 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n53, SL => mult_21_C241_n894, Z => 
                           mult_21_C241_n1197);
   mult_21_C241_U770 : MUXB2DL port map( A0 => mult_21_C241_n1539, A1 => 
                           mult_21_C241_n1538, SL => mult_21_C241_n56, Z => 
                           mult_21_C241_n893);
   mult_21_C241_U769 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n53, SL => mult_21_C241_n893, Z => 
                           mult_21_C241_n1196);
   mult_21_C241_U768 : MUXB2DL port map( A0 => mult_21_C241_n1540, A1 => 
                           mult_21_C241_n1539, SL => mult_21_C241_n56, Z => 
                           mult_21_C241_n892);
   mult_21_C241_U767 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n53, SL => mult_21_C241_n892, Z => 
                           mult_21_C241_n1195);
   mult_21_C241_U766 : MUXB2DL port map( A0 => N3085, A1 => mult_21_C241_n1540,
                           SL => mult_21_C241_n56, Z => mult_21_C241_n891);
   mult_21_C241_U765 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n53, SL => mult_21_C241_n891, Z => 
                           mult_21_C241_n1194);
   mult_21_C241_U764 : MUXB2DL port map( A0 => N3086, A1 => N3085, SL => 
                           mult_21_C241_n56, Z => mult_21_C241_n890);
   mult_21_C241_U763 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n53, SL => mult_21_C241_n890, Z => 
                           mult_21_C241_n1193);
   mult_21_C241_U762 : MUXB2DL port map( A0 => N3087, A1 => N3086, SL => 
                           mult_21_C241_n56, Z => mult_21_C241_n889);
   mult_21_C241_U761 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n53, SL => mult_21_C241_n889, Z => 
                           mult_21_C241_n1192);
   mult_21_C241_U760 : MUXB2DL port map( A0 => N3088, A1 => N3087, SL => 
                           mult_21_C241_n56, Z => mult_21_C241_n888);
   mult_21_C241_U759 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n53, SL => mult_21_C241_n888, Z => 
                           mult_21_C241_n1191);
   mult_21_C241_U758 : MUXB2DL port map( A0 => N3089, A1 => N3088, SL => 
                           mult_21_C241_n56, Z => mult_21_C241_n887);
   mult_21_C241_U757 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n53, SL => mult_21_C241_n887, Z => 
                           mult_21_C241_n1190);
   mult_21_C241_U756 : MUXB2DL port map( A0 => N3090, A1 => N3089, SL => 
                           mult_21_C241_n56, Z => mult_21_C241_n886);
   mult_21_C241_U755 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n53, SL => mult_21_C241_n886, Z => 
                           mult_21_C241_n1189);
   mult_21_C241_U754 : MUXB2DL port map( A0 => N3091, A1 => N3090, SL => 
                           mult_21_C241_n56, Z => mult_21_C241_n885);
   mult_21_C241_U753 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n53, SL => mult_21_C241_n885, Z => 
                           mult_21_C241_n1188);
   mult_21_C241_U752 : MUXB2DL port map( A0 => N3092, A1 => N3091, SL => 
                           mult_21_C241_n56, Z => mult_21_C241_n884);
   mult_21_C241_U751 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n53, SL => mult_21_C241_n884, Z => 
                           mult_21_C241_n1187);
   mult_21_C241_U750 : NOR2M1D1 port map( A1 => mult_21_C241_n50, A2 => 
                           mult_21_C241_n53, Z => mult_21_C241_n1090);
   mult_21_C241_U749 : NAN2M1D1 port map( A1 => mult_21_C241_n63, A2 => N3073, 
                           Z => mult_21_C241_n883);
   mult_21_C241_U748 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n61, SL => mult_21_C241_n883, Z => 
                           mult_21_C241_n1186);
   mult_21_C241_U747 : MUXB2DL port map( A0 => N3074, A1 => mult_21_C241_n1548,
                           SL => mult_21_C241_n63, Z => mult_21_C241_n882);
   mult_21_C241_U746 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n61, SL => mult_21_C241_n882, Z => 
                           mult_21_C241_n1185);
   mult_21_C241_U745 : MUXB2DL port map( A0 => mult_21_C241_n1546, A1 => N3074,
                           SL => mult_21_C241_n63, Z => mult_21_C241_n881);
   mult_21_C241_U744 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n61, SL => mult_21_C241_n881, Z => 
                           mult_21_C241_n1184);
   mult_21_C241_U743 : MUXB2DL port map( A0 => N3076, A1 => mult_21_C241_n1546,
                           SL => mult_21_C241_n63, Z => mult_21_C241_n880);
   mult_21_C241_U742 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n61, SL => mult_21_C241_n880, Z => 
                           mult_21_C241_n1183);
   mult_21_C241_U741 : MUXB2DL port map( A0 => N3077, A1 => N3076, SL => 
                           mult_21_C241_n63, Z => mult_21_C241_n879);
   mult_21_C241_U740 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n61, SL => mult_21_C241_n879, Z => 
                           mult_21_C241_n1182);
   mult_21_C241_U739 : MUXB2DL port map( A0 => N3078, A1 => N3077, SL => 
                           mult_21_C241_n63, Z => mult_21_C241_n878);
   mult_21_C241_U738 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n61, SL => mult_21_C241_n878, Z => 
                           mult_21_C241_n1181);
   mult_21_C241_U737 : MUXB2DL port map( A0 => N3079, A1 => N3078, SL => 
                           mult_21_C241_n63, Z => mult_21_C241_n877);
   mult_21_C241_U736 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n61, SL => mult_21_C241_n877, Z => 
                           mult_21_C241_n1180);
   mult_21_C241_U735 : MUXB2DL port map( A0 => N3080, A1 => N3079, SL => 
                           mult_21_C241_n63, Z => mult_21_C241_n876);
   mult_21_C241_U734 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n61, SL => mult_21_C241_n876, Z => 
                           mult_21_C241_n1179);
   mult_21_C241_U733 : MUXB2DL port map( A0 => N3081, A1 => N3080, SL => 
                           mult_21_C241_n63, Z => mult_21_C241_n875);
   mult_21_C241_U732 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n61, SL => mult_21_C241_n875, Z => 
                           mult_21_C241_n1178);
   mult_21_C241_U731 : MUXB2DL port map( A0 => mult_21_C241_n1538, A1 => N3081,
                           SL => mult_21_C241_n63, Z => mult_21_C241_n874);
   mult_21_C241_U730 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n61, SL => mult_21_C241_n874, Z => 
                           mult_21_C241_n1177);
   mult_21_C241_U729 : MUXB2DL port map( A0 => mult_21_C241_n1539, A1 => 
                           mult_21_C241_n1538, SL => mult_21_C241_n63, Z => 
                           mult_21_C241_n873);
   mult_21_C241_U728 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n61, SL => mult_21_C241_n873, Z => 
                           mult_21_C241_n1176);
   mult_21_C241_U727 : MUXB2DL port map( A0 => mult_21_C241_n1540, A1 => 
                           mult_21_C241_n1539, SL => mult_21_C241_n63, Z => 
                           mult_21_C241_n872);
   mult_21_C241_U726 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n61, SL => mult_21_C241_n872, Z => 
                           mult_21_C241_n1175);
   mult_21_C241_U725 : MUXB2DL port map( A0 => N3085, A1 => mult_21_C241_n1540,
                           SL => mult_21_C241_n63, Z => mult_21_C241_n871);
   mult_21_C241_U724 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n61, SL => mult_21_C241_n871, Z => 
                           mult_21_C241_n1174);
   mult_21_C241_U723 : MUXB2DL port map( A0 => N3086, A1 => N3085, SL => 
                           mult_21_C241_n63, Z => mult_21_C241_n870);
   mult_21_C241_U722 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n61, SL => mult_21_C241_n870, Z => 
                           mult_21_C241_n1173);
   mult_21_C241_U721 : MUXB2DL port map( A0 => N3087, A1 => N3086, SL => 
                           mult_21_C241_n63, Z => mult_21_C241_n869);
   mult_21_C241_U720 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n61, SL => mult_21_C241_n869, Z => 
                           mult_21_C241_n1172);
   mult_21_C241_U719 : MUXB2DL port map( A0 => N3088, A1 => N3087, SL => 
                           mult_21_C241_n63, Z => mult_21_C241_n868);
   mult_21_C241_U718 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n61, SL => mult_21_C241_n868, Z => 
                           mult_21_C241_n1171);
   mult_21_C241_U717 : MUXB2DL port map( A0 => N3089, A1 => N3088, SL => 
                           mult_21_C241_n63, Z => mult_21_C241_n867);
   mult_21_C241_U716 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n61, SL => mult_21_C241_n867, Z => 
                           mult_21_C241_n1170);
   mult_21_C241_U715 : MUXB2DL port map( A0 => N3090, A1 => N3089, SL => 
                           mult_21_C241_n63, Z => mult_21_C241_n866);
   mult_21_C241_U714 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n61, SL => mult_21_C241_n866, Z => 
                           mult_21_C241_n1169);
   mult_21_C241_U713 : NOR2M1D1 port map( A1 => mult_21_C241_n58, A2 => 
                           mult_21_C241_n61, Z => mult_21_C241_n1089);
   mult_21_C241_U712 : NAN2M1D1 port map( A1 => mult_21_C241_n71, A2 => N3073, 
                           Z => mult_21_C241_n865);
   mult_21_C241_U711 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n69, SL => mult_21_C241_n865, Z => 
                           mult_21_C241_n1168);
   mult_21_C241_U710 : MUXB2DL port map( A0 => N3074, A1 => mult_21_C241_n1548,
                           SL => mult_21_C241_n71, Z => mult_21_C241_n864);
   mult_21_C241_U709 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n69, SL => mult_21_C241_n864, Z => 
                           mult_21_C241_n1167);
   mult_21_C241_U708 : MUXB2DL port map( A0 => N3075, A1 => N3074, SL => 
                           mult_21_C241_n71, Z => mult_21_C241_n863);
   mult_21_C241_U707 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n69, SL => mult_21_C241_n863, Z => 
                           mult_21_C241_n1166);
   mult_21_C241_U706 : MUXB2DL port map( A0 => N3076, A1 => mult_21_C241_n1546,
                           SL => mult_21_C241_n71, Z => mult_21_C241_n862);
   mult_21_C241_U705 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n69, SL => mult_21_C241_n862, Z => 
                           mult_21_C241_n1165);
   mult_21_C241_U704 : MUXB2DL port map( A0 => N3077, A1 => N3076, SL => 
                           mult_21_C241_n71, Z => mult_21_C241_n861);
   mult_21_C241_U703 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n69, SL => mult_21_C241_n861, Z => 
                           mult_21_C241_n1164);
   mult_21_C241_U702 : MUXB2DL port map( A0 => N3078, A1 => N3077, SL => 
                           mult_21_C241_n71, Z => mult_21_C241_n860);
   mult_21_C241_U701 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n69, SL => mult_21_C241_n860, Z => 
                           mult_21_C241_n1163);
   mult_21_C241_U700 : MUXB2DL port map( A0 => N3079, A1 => N3078, SL => 
                           mult_21_C241_n71, Z => mult_21_C241_n859);
   mult_21_C241_U699 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n69, SL => mult_21_C241_n859, Z => 
                           mult_21_C241_n1162);
   mult_21_C241_U698 : MUXB2DL port map( A0 => N3080, A1 => N3079, SL => 
                           mult_21_C241_n71, Z => mult_21_C241_n858);
   mult_21_C241_U697 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n69, SL => mult_21_C241_n858, Z => 
                           mult_21_C241_n1161);
   mult_21_C241_U696 : MUXB2DL port map( A0 => N3081, A1 => N3080, SL => 
                           mult_21_C241_n71, Z => mult_21_C241_n857);
   mult_21_C241_U695 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n69, SL => mult_21_C241_n857, Z => 
                           mult_21_C241_n1160);
   mult_21_C241_U694 : MUXB2DL port map( A0 => mult_21_C241_n1538, A1 => N3081,
                           SL => mult_21_C241_n71, Z => mult_21_C241_n856);
   mult_21_C241_U693 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n69, SL => mult_21_C241_n856, Z => 
                           mult_21_C241_n1159);
   mult_21_C241_U692 : MUXB2DL port map( A0 => mult_21_C241_n1539, A1 => 
                           mult_21_C241_n1538, SL => mult_21_C241_n71, Z => 
                           mult_21_C241_n855);
   mult_21_C241_U691 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n69, SL => mult_21_C241_n855, Z => 
                           mult_21_C241_n1158);
   mult_21_C241_U690 : MUXB2DL port map( A0 => mult_21_C241_n1540, A1 => 
                           mult_21_C241_n1539, SL => mult_21_C241_n71, Z => 
                           mult_21_C241_n854);
   mult_21_C241_U689 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n69, SL => mult_21_C241_n854, Z => 
                           mult_21_C241_n1157);
   mult_21_C241_U688 : MUXB2DL port map( A0 => N3085, A1 => mult_21_C241_n1540,
                           SL => mult_21_C241_n71, Z => mult_21_C241_n853);
   mult_21_C241_U687 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n69, SL => mult_21_C241_n853, Z => 
                           mult_21_C241_n1156);
   mult_21_C241_U686 : MUXB2DL port map( A0 => N3086, A1 => N3085, SL => 
                           mult_21_C241_n71, Z => mult_21_C241_n852);
   mult_21_C241_U685 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n69, SL => mult_21_C241_n852, Z => 
                           mult_21_C241_n1155);
   mult_21_C241_U684 : MUXB2DL port map( A0 => N3087, A1 => N3086, SL => 
                           mult_21_C241_n71, Z => mult_21_C241_n851);
   mult_21_C241_U683 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n69, SL => mult_21_C241_n851, Z => 
                           mult_21_C241_n1154);
   mult_21_C241_U682 : MUXB2DL port map( A0 => N3088, A1 => N3087, SL => 
                           mult_21_C241_n71, Z => mult_21_C241_n850);
   mult_21_C241_U681 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n69, SL => mult_21_C241_n850, Z => 
                           mult_21_C241_n1153);
   mult_21_C241_U680 : NOR2M1D1 port map( A1 => mult_21_C241_n66, A2 => 
                           mult_21_C241_n69, Z => mult_21_C241_n1088);
   mult_21_C241_U679 : NAN2M1D1 port map( A1 => mult_21_C241_n78, A2 => 
                           mult_21_C241_n1548, Z => mult_21_C241_n849);
   mult_21_C241_U678 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n76, SL => mult_21_C241_n849, Z => 
                           mult_21_C241_n1152);
   mult_21_C241_U677 : MUXB2DL port map( A0 => N3074, A1 => mult_21_C241_n1548,
                           SL => mult_21_C241_n78, Z => mult_21_C241_n848);
   mult_21_C241_U676 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n76, SL => mult_21_C241_n848, Z => 
                           mult_21_C241_n1151);
   mult_21_C241_U675 : MUXB2DL port map( A0 => mult_21_C241_n1546, A1 => N3074,
                           SL => mult_21_C241_n78, Z => mult_21_C241_n847);
   mult_21_C241_U674 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n76, SL => mult_21_C241_n847, Z => 
                           mult_21_C241_n1150);
   mult_21_C241_U673 : MUXB2DL port map( A0 => N3076, A1 => mult_21_C241_n1546,
                           SL => mult_21_C241_n78, Z => mult_21_C241_n846);
   mult_21_C241_U672 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n76, SL => mult_21_C241_n846, Z => 
                           mult_21_C241_n1149);
   mult_21_C241_U671 : MUXB2DL port map( A0 => N3077, A1 => N3076, SL => 
                           mult_21_C241_n78, Z => mult_21_C241_n845);
   mult_21_C241_U670 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n76, SL => mult_21_C241_n845, Z => 
                           mult_21_C241_n1148);
   mult_21_C241_U669 : MUXB2DL port map( A0 => N3078, A1 => N3077, SL => 
                           mult_21_C241_n78, Z => mult_21_C241_n844);
   mult_21_C241_U668 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n76, SL => mult_21_C241_n844, Z => 
                           mult_21_C241_n1147);
   mult_21_C241_U667 : MUXB2DL port map( A0 => N3079, A1 => N3078, SL => 
                           mult_21_C241_n78, Z => mult_21_C241_n843);
   mult_21_C241_U666 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n76, SL => mult_21_C241_n843, Z => 
                           mult_21_C241_n1146);
   mult_21_C241_U665 : MUXB2DL port map( A0 => N3080, A1 => N3079, SL => 
                           mult_21_C241_n78, Z => mult_21_C241_n842);
   mult_21_C241_U664 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n76, SL => mult_21_C241_n842, Z => 
                           mult_21_C241_n1145);
   mult_21_C241_U663 : MUXB2DL port map( A0 => N3081, A1 => N3080, SL => 
                           mult_21_C241_n78, Z => mult_21_C241_n841);
   mult_21_C241_U662 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n76, SL => mult_21_C241_n841, Z => 
                           mult_21_C241_n1144);
   mult_21_C241_U661 : MUXB2DL port map( A0 => mult_21_C241_n1538, A1 => N3081,
                           SL => mult_21_C241_n78, Z => mult_21_C241_n840);
   mult_21_C241_U660 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n76, SL => mult_21_C241_n840, Z => 
                           mult_21_C241_n1143);
   mult_21_C241_U659 : MUXB2DL port map( A0 => mult_21_C241_n1539, A1 => 
                           mult_21_C241_n1538, SL => mult_21_C241_n78, Z => 
                           mult_21_C241_n839);
   mult_21_C241_U658 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n76, SL => mult_21_C241_n839, Z => 
                           mult_21_C241_n1142);
   mult_21_C241_U657 : MUXB2DL port map( A0 => mult_21_C241_n1540, A1 => 
                           mult_21_C241_n1539, SL => mult_21_C241_n78, Z => 
                           mult_21_C241_n838);
   mult_21_C241_U656 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n76, SL => mult_21_C241_n838, Z => 
                           mult_21_C241_n1141);
   mult_21_C241_U655 : MUXB2DL port map( A0 => N3085, A1 => mult_21_C241_n1540,
                           SL => mult_21_C241_n78, Z => mult_21_C241_n837);
   mult_21_C241_U654 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n76, SL => mult_21_C241_n837, Z => 
                           mult_21_C241_n1140);
   mult_21_C241_U653 : MUXB2DL port map( A0 => N3086, A1 => N3085, SL => 
                           mult_21_C241_n78, Z => mult_21_C241_n836);
   mult_21_C241_U652 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n76, SL => mult_21_C241_n836, Z => 
                           mult_21_C241_n1139);
   mult_21_C241_U651 : NOR2M1D1 port map( A1 => mult_21_C241_n73, A2 => 
                           mult_21_C241_n76, Z => mult_21_C241_n1087);
   mult_21_C241_U650 : NAN2M1D1 port map( A1 => mult_21_C241_n83, A2 => N3073, 
                           Z => mult_21_C241_n835);
   mult_21_C241_U649 : MUXB2DL port map( A0 => mult_21_C241_n79, A1 => 
                           mult_21_C241_n81, SL => mult_21_C241_n835, Z => 
                           mult_21_C241_n1138);
   mult_21_C241_U648 : MUXB2DL port map( A0 => N3074, A1 => mult_21_C241_n1548,
                           SL => mult_21_C241_n83, Z => mult_21_C241_n834);
   mult_21_C241_U647 : MUXB2DL port map( A0 => mult_21_C241_n79, A1 => 
                           mult_21_C241_n81, SL => mult_21_C241_n834, Z => 
                           mult_21_C241_n1137);
   mult_21_C241_U646 : MUXB2DL port map( A0 => mult_21_C241_n1546, A1 => N3074,
                           SL => mult_21_C241_n83, Z => mult_21_C241_n833);
   mult_21_C241_U645 : MUXB2DL port map( A0 => mult_21_C241_n79, A1 => 
                           mult_21_C241_n81, SL => mult_21_C241_n833, Z => 
                           mult_21_C241_n1136);
   mult_21_C241_U644 : MUXB2DL port map( A0 => N3076, A1 => mult_21_C241_n1546,
                           SL => mult_21_C241_n83, Z => mult_21_C241_n832);
   mult_21_C241_U643 : MUXB2DL port map( A0 => mult_21_C241_n79, A1 => 
                           mult_21_C241_n81, SL => mult_21_C241_n832, Z => 
                           mult_21_C241_n1135);
   mult_21_C241_U642 : MUXB2DL port map( A0 => N3077, A1 => N3076, SL => 
                           mult_21_C241_n83, Z => mult_21_C241_n831);
   mult_21_C241_U641 : MUXB2DL port map( A0 => mult_21_C241_n79, A1 => 
                           mult_21_C241_n81, SL => mult_21_C241_n831, Z => 
                           mult_21_C241_n1134);
   mult_21_C241_U640 : MUXB2DL port map( A0 => N3078, A1 => N3077, SL => 
                           mult_21_C241_n83, Z => mult_21_C241_n830);
   mult_21_C241_U639 : MUXB2DL port map( A0 => mult_21_C241_n79, A1 => 
                           mult_21_C241_n81, SL => mult_21_C241_n830, Z => 
                           mult_21_C241_n1133);
   mult_21_C241_U638 : MUXB2DL port map( A0 => N3079, A1 => N3078, SL => 
                           mult_21_C241_n83, Z => mult_21_C241_n829);
   mult_21_C241_U637 : MUXB2DL port map( A0 => mult_21_C241_n79, A1 => 
                           mult_21_C241_n81, SL => mult_21_C241_n829, Z => 
                           mult_21_C241_n1132);
   mult_21_C241_U636 : MUXB2DL port map( A0 => N3080, A1 => N3079, SL => 
                           mult_21_C241_n83, Z => mult_21_C241_n828);
   mult_21_C241_U635 : MUXB2DL port map( A0 => mult_21_C241_n79, A1 => 
                           mult_21_C241_n81, SL => mult_21_C241_n828, Z => 
                           mult_21_C241_n1131);
   mult_21_C241_U634 : MUXB2DL port map( A0 => N3081, A1 => N3080, SL => 
                           mult_21_C241_n83, Z => mult_21_C241_n827);
   mult_21_C241_U633 : MUXB2DL port map( A0 => mult_21_C241_n79, A1 => 
                           mult_21_C241_n81, SL => mult_21_C241_n827, Z => 
                           mult_21_C241_n1130);
   mult_21_C241_U632 : MUXB2DL port map( A0 => mult_21_C241_n1538, A1 => N3081,
                           SL => mult_21_C241_n83, Z => mult_21_C241_n826);
   mult_21_C241_U631 : MUXB2DL port map( A0 => mult_21_C241_n79, A1 => 
                           mult_21_C241_n81, SL => mult_21_C241_n826, Z => 
                           mult_21_C241_n1129);
   mult_21_C241_U630 : MUXB2DL port map( A0 => mult_21_C241_n1539, A1 => 
                           mult_21_C241_n1538, SL => mult_21_C241_n83, Z => 
                           mult_21_C241_n825);
   mult_21_C241_U629 : MUXB2DL port map( A0 => mult_21_C241_n79, A1 => 
                           mult_21_C241_n81, SL => mult_21_C241_n825, Z => 
                           mult_21_C241_n1128);
   mult_21_C241_U628 : MUXB2DL port map( A0 => mult_21_C241_n1540, A1 => 
                           mult_21_C241_n1539, SL => mult_21_C241_n83, Z => 
                           mult_21_C241_n824);
   mult_21_C241_U627 : MUXB2DL port map( A0 => mult_21_C241_n79, A1 => 
                           mult_21_C241_n81, SL => mult_21_C241_n824, Z => 
                           mult_21_C241_n1127);
   mult_21_C241_U626 : NOR2M1D1 port map( A1 => mult_21_C241_n79, A2 => 
                           mult_21_C241_n81, Z => mult_21_C241_n1086);
   mult_21_C241_U625 : NAN2M1D1 port map( A1 => mult_21_C241_n88, A2 => 
                           mult_21_C241_n1548, Z => mult_21_C241_n823);
   mult_21_C241_U624 : MUXB2DL port map( A0 => mult_21_C241_n84, A1 => 
                           mult_21_C241_n86, SL => mult_21_C241_n823, Z => 
                           mult_21_C241_n1126);
   mult_21_C241_U623 : MUXB2DL port map( A0 => N3074, A1 => mult_21_C241_n1548,
                           SL => mult_21_C241_n88, Z => mult_21_C241_n822);
   mult_21_C241_U622 : MUXB2DL port map( A0 => mult_21_C241_n84, A1 => 
                           mult_21_C241_n86, SL => mult_21_C241_n822, Z => 
                           mult_21_C241_n1125);
   mult_21_C241_U621 : MUXB2DL port map( A0 => N3075, A1 => N3074, SL => 
                           mult_21_C241_n88, Z => mult_21_C241_n821);
   mult_21_C241_U620 : MUXB2DL port map( A0 => mult_21_C241_n84, A1 => 
                           mult_21_C241_n86, SL => mult_21_C241_n821, Z => 
                           mult_21_C241_n1124);
   mult_21_C241_U619 : MUXB2DL port map( A0 => N3076, A1 => mult_21_C241_n1546,
                           SL => mult_21_C241_n88, Z => mult_21_C241_n820);
   mult_21_C241_U618 : MUXB2DL port map( A0 => mult_21_C241_n84, A1 => 
                           mult_21_C241_n86, SL => mult_21_C241_n820, Z => 
                           mult_21_C241_n1123);
   mult_21_C241_U617 : MUXB2DL port map( A0 => N3077, A1 => N3076, SL => 
                           mult_21_C241_n88, Z => mult_21_C241_n819);
   mult_21_C241_U616 : MUXB2DL port map( A0 => mult_21_C241_n84, A1 => 
                           mult_21_C241_n86, SL => mult_21_C241_n819, Z => 
                           mult_21_C241_n1122);
   mult_21_C241_U615 : MUXB2DL port map( A0 => N3078, A1 => N3077, SL => 
                           mult_21_C241_n88, Z => mult_21_C241_n818);
   mult_21_C241_U614 : MUXB2DL port map( A0 => mult_21_C241_n84, A1 => 
                           mult_21_C241_n86, SL => mult_21_C241_n818, Z => 
                           mult_21_C241_n1121);
   mult_21_C241_U613 : MUXB2DL port map( A0 => N3079, A1 => N3078, SL => 
                           mult_21_C241_n88, Z => mult_21_C241_n817);
   mult_21_C241_U612 : MUXB2DL port map( A0 => mult_21_C241_n84, A1 => 
                           mult_21_C241_n86, SL => mult_21_C241_n817, Z => 
                           mult_21_C241_n1120);
   mult_21_C241_U611 : MUXB2DL port map( A0 => N3080, A1 => N3079, SL => 
                           mult_21_C241_n88, Z => mult_21_C241_n816);
   mult_21_C241_U610 : MUXB2DL port map( A0 => mult_21_C241_n84, A1 => 
                           mult_21_C241_n86, SL => mult_21_C241_n816, Z => 
                           mult_21_C241_n1119);
   mult_21_C241_U609 : MUXB2DL port map( A0 => N3081, A1 => N3080, SL => 
                           mult_21_C241_n88, Z => mult_21_C241_n815);
   mult_21_C241_U608 : MUXB2DL port map( A0 => mult_21_C241_n84, A1 => 
                           mult_21_C241_n86, SL => mult_21_C241_n815, Z => 
                           mult_21_C241_n1118);
   mult_21_C241_U607 : MUXB2DL port map( A0 => mult_21_C241_n1538, A1 => N3081,
                           SL => mult_21_C241_n88, Z => mult_21_C241_n814);
   mult_21_C241_U606 : MUXB2DL port map( A0 => mult_21_C241_n84, A1 => 
                           mult_21_C241_n86, SL => mult_21_C241_n814, Z => 
                           mult_21_C241_n1117);
   mult_21_C241_U605 : NOR2M1D1 port map( A1 => mult_21_C241_n84, A2 => 
                           mult_21_C241_n86, Z => mult_21_C241_n1085);
   mult_21_C241_U604 : NAN2M1D1 port map( A1 => mult_21_C241_n93, A2 => 
                           mult_21_C241_n1548, Z => mult_21_C241_n813);
   mult_21_C241_U603 : MUXB2DL port map( A0 => mult_21_C241_n89, A1 => 
                           mult_21_C241_n91, SL => mult_21_C241_n813, Z => 
                           mult_21_C241_n1116);
   mult_21_C241_U602 : MUXB2DL port map( A0 => N3074, A1 => mult_21_C241_n1548,
                           SL => mult_21_C241_n93, Z => mult_21_C241_n812);
   mult_21_C241_U601 : MUXB2DL port map( A0 => mult_21_C241_n89, A1 => 
                           mult_21_C241_n91, SL => mult_21_C241_n812, Z => 
                           mult_21_C241_n1115);
   mult_21_C241_U600 : MUXB2DL port map( A0 => N3075, A1 => N3074, SL => 
                           mult_21_C241_n93, Z => mult_21_C241_n811);
   mult_21_C241_U599 : MUXB2DL port map( A0 => mult_21_C241_n89, A1 => 
                           mult_21_C241_n91, SL => mult_21_C241_n811, Z => 
                           mult_21_C241_n1114);
   mult_21_C241_U598 : MUXB2DL port map( A0 => N3076, A1 => mult_21_C241_n1546,
                           SL => mult_21_C241_n93, Z => mult_21_C241_n810);
   mult_21_C241_U597 : MUXB2DL port map( A0 => mult_21_C241_n89, A1 => 
                           mult_21_C241_n91, SL => mult_21_C241_n810, Z => 
                           mult_21_C241_n1113);
   mult_21_C241_U596 : MUXB2DL port map( A0 => N3077, A1 => N3076, SL => 
                           mult_21_C241_n93, Z => mult_21_C241_n809);
   mult_21_C241_U595 : MUXB2DL port map( A0 => mult_21_C241_n89, A1 => 
                           mult_21_C241_n91, SL => mult_21_C241_n809, Z => 
                           mult_21_C241_n1112);
   mult_21_C241_U594 : MUXB2DL port map( A0 => N3078, A1 => N3077, SL => 
                           mult_21_C241_n93, Z => mult_21_C241_n808);
   mult_21_C241_U593 : MUXB2DL port map( A0 => mult_21_C241_n89, A1 => 
                           mult_21_C241_n91, SL => mult_21_C241_n808, Z => 
                           mult_21_C241_n1111);
   mult_21_C241_U592 : MUXB2DL port map( A0 => N3079, A1 => N3078, SL => 
                           mult_21_C241_n93, Z => mult_21_C241_n807);
   mult_21_C241_U591 : MUXB2DL port map( A0 => mult_21_C241_n89, A1 => 
                           mult_21_C241_n91, SL => mult_21_C241_n807, Z => 
                           mult_21_C241_n1110);
   mult_21_C241_U590 : MUXB2DL port map( A0 => N3080, A1 => N3079, SL => 
                           mult_21_C241_n93, Z => mult_21_C241_n806);
   mult_21_C241_U589 : MUXB2DL port map( A0 => mult_21_C241_n89, A1 => 
                           mult_21_C241_n91, SL => mult_21_C241_n806, Z => 
                           mult_21_C241_n1109);
   mult_21_C241_U588 : NOR2M1D1 port map( A1 => mult_21_C241_n89, A2 => 
                           mult_21_C241_n91, Z => mult_21_C241_n1084);
   mult_21_C241_U587 : NAN2M1D1 port map( A1 => mult_21_C241_n98, A2 => N3073, 
                           Z => mult_21_C241_n805);
   mult_21_C241_U586 : MUXB2DL port map( A0 => mult_21_C241_n94, A1 => 
                           mult_21_C241_n96, SL => mult_21_C241_n805, Z => 
                           mult_21_C241_n1108);
   mult_21_C241_U585 : MUXB2DL port map( A0 => N3074, A1 => mult_21_C241_n1548,
                           SL => mult_21_C241_n98, Z => mult_21_C241_n804);
   mult_21_C241_U584 : MUXB2DL port map( A0 => mult_21_C241_n94, A1 => 
                           mult_21_C241_n96, SL => mult_21_C241_n804, Z => 
                           mult_21_C241_n1107);
   mult_21_C241_U583 : MUXB2DL port map( A0 => N3075, A1 => N3074, SL => 
                           mult_21_C241_n98, Z => mult_21_C241_n803);
   mult_21_C241_U582 : MUXB2DL port map( A0 => mult_21_C241_n94, A1 => 
                           mult_21_C241_n96, SL => mult_21_C241_n803, Z => 
                           mult_21_C241_n1106);
   mult_21_C241_U581 : MUXB2DL port map( A0 => N3076, A1 => mult_21_C241_n1546,
                           SL => mult_21_C241_n98, Z => mult_21_C241_n802);
   mult_21_C241_U580 : MUXB2DL port map( A0 => mult_21_C241_n94, A1 => 
                           mult_21_C241_n96, SL => mult_21_C241_n802, Z => 
                           mult_21_C241_n1105);
   mult_21_C241_U579 : MUXB2DL port map( A0 => N3077, A1 => N3076, SL => 
                           mult_21_C241_n98, Z => mult_21_C241_n801);
   mult_21_C241_U578 : MUXB2DL port map( A0 => mult_21_C241_n94, A1 => 
                           mult_21_C241_n96, SL => mult_21_C241_n801, Z => 
                           mult_21_C241_n1104);
   mult_21_C241_U577 : MUXB2DL port map( A0 => N3078, A1 => N3077, SL => 
                           mult_21_C241_n98, Z => mult_21_C241_n800);
   mult_21_C241_U576 : MUXB2DL port map( A0 => mult_21_C241_n94, A1 => 
                           mult_21_C241_n96, SL => mult_21_C241_n800, Z => 
                           mult_21_C241_n1103);
   mult_21_C241_U575 : NOR2M1D1 port map( A1 => mult_21_C241_n94, A2 => 
                           mult_21_C241_n96, Z => mult_21_C241_n1083);
   mult_21_C241_U574 : NAN2M1D1 port map( A1 => mult_21_C241_n103, A2 => N3073,
                           Z => mult_21_C241_n799);
   mult_21_C241_U573 : MUXB2DL port map( A0 => mult_21_C241_n99, A1 => 
                           mult_21_C241_n101, SL => mult_21_C241_n799, Z => 
                           mult_21_C241_n1102);
   mult_21_C241_U572 : MUXB2DL port map( A0 => N3074, A1 => mult_21_C241_n1548,
                           SL => mult_21_C241_n103, Z => mult_21_C241_n798);
   mult_21_C241_U571 : MUXB2DL port map( A0 => mult_21_C241_n99, A1 => 
                           mult_21_C241_n101, SL => mult_21_C241_n798, Z => 
                           mult_21_C241_n1101);
   mult_21_C241_U570 : MUXB2DL port map( A0 => N3075, A1 => N3074, SL => 
                           mult_21_C241_n103, Z => mult_21_C241_n797);
   mult_21_C241_U569 : MUXB2DL port map( A0 => mult_21_C241_n99, A1 => 
                           mult_21_C241_n101, SL => mult_21_C241_n797, Z => 
                           mult_21_C241_n1100);
   mult_21_C241_U568 : MUXB2DL port map( A0 => N3076, A1 => mult_21_C241_n1546,
                           SL => mult_21_C241_n103, Z => mult_21_C241_n796);
   mult_21_C241_U567 : MUXB2DL port map( A0 => mult_21_C241_n99, A1 => 
                           mult_21_C241_n101, SL => mult_21_C241_n796, Z => 
                           mult_21_C241_n1099);
   mult_21_C241_U566 : NOR2M1D1 port map( A1 => mult_21_C241_n99, A2 => 
                           mult_21_C241_n101, Z => mult_21_C241_n1082);
   mult_21_C241_U565 : NAN2M1D1 port map( A1 => mult_21_C241_n106, A2 => N3073,
                           Z => mult_21_C241_n795);
   mult_21_C241_U564 : MUXB2DL port map( A0 => mult_21_C241_n104, A1 => 
                           mult_21_C241_n105, SL => mult_21_C241_n795, Z => 
                           mult_21_C241_n1098);
   mult_21_C241_U563 : MUXB2DL port map( A0 => N3074, A1 => mult_21_C241_n1548,
                           SL => mult_21_C241_n106, Z => mult_21_C241_n794);
   mult_21_C241_U562 : MUXB2DL port map( A0 => mult_21_C241_n104, A1 => 
                           mult_21_C241_n105, SL => mult_21_C241_n794, Z => 
                           mult_21_C241_n1097);
   mult_21_C241_U561 : NOR2M1D1 port map( A1 => mult_21_C241_n104, A2 => 
                           mult_21_C241_n105, Z => mult_21_C241_n1081);
   mult_21_C241_U557 : ADFULD1 port map( A => mult_21_C241_n1334, B => 
                           mult_21_C241_n1364, CI => mult_21_C241_n790, CO => 
                           mult_21_C241_n786, S => mult_21_C241_n787);
   mult_21_C241_U555 : ADFULD1 port map( A => mult_21_C241_n788, B => 
                           mult_21_C241_n1305, CI => mult_21_C241_n785, CO => 
                           mult_21_C241_n782, S => mult_21_C241_n783);
   mult_21_C241_U553 : ADFULD1 port map( A => mult_21_C241_n1304, B => 
                           mult_21_C241_n1362, CI => mult_21_C241_n1332, CO => 
                           mult_21_C241_n778, S => mult_21_C241_n779);
   mult_21_C241_U552 : ADFULD1 port map( A => mult_21_C241_n781, B => 
                           mult_21_C241_n784, CI => mult_21_C241_n779, CO => 
                           mult_21_C241_n776, S => mult_21_C241_n777);
   mult_21_C241_U550 : ADFULD1 port map( A => mult_21_C241_n1277, B => 
                           mult_21_C241_n1303, CI => mult_21_C241_n780, CO => 
                           mult_21_C241_n772, S => mult_21_C241_n773);
   mult_21_C241_U549 : ADFULD1 port map( A => mult_21_C241_n778, B => 
                           mult_21_C241_n775, CI => mult_21_C241_n773, CO => 
                           mult_21_C241_n770, S => mult_21_C241_n771);
   mult_21_C241_U547 : ADFULD1 port map( A => mult_21_C241_n1276, B => 
                           mult_21_C241_n1360, CI => mult_21_C241_n1330, CO => 
                           mult_21_C241_n766, S => mult_21_C241_n767);
   mult_21_C241_U546 : ADFULD1 port map( A => mult_21_C241_n774, B => 
                           mult_21_C241_n1302, CI => mult_21_C241_n769, CO => 
                           mult_21_C241_n764, S => mult_21_C241_n765);
   mult_21_C241_U545 : ADFULD1 port map( A => mult_21_C241_n767, B => 
                           mult_21_C241_n772, CI => mult_21_C241_n765, CO => 
                           mult_21_C241_n762, S => mult_21_C241_n763);
   mult_21_C241_U543 : ADFULD1 port map( A => mult_21_C241_n1275, B => 
                           mult_21_C241_n1251, CI => mult_21_C241_n1301, CO => 
                           mult_21_C241_n758, S => mult_21_C241_n759);
   mult_21_C241_U542 : ADFULD1 port map( A => mult_21_C241_n761, B => 
                           mult_21_C241_n768, CI => mult_21_C241_n766, CO => 
                           mult_21_C241_n756, S => mult_21_C241_n757);
   mult_21_C241_U541 : ADFULD1 port map( A => mult_21_C241_n764, B => 
                           mult_21_C241_n759, CI => mult_21_C241_n757, CO => 
                           mult_21_C241_n754, S => mult_21_C241_n755);
   mult_21_C241_U539 : ADFULD1 port map( A => mult_21_C241_n1250, B => 
                           mult_21_C241_n1358, CI => mult_21_C241_n1328, CO => 
                           mult_21_C241_n750, S => mult_21_C241_n751);
   mult_21_C241_U538 : ADFULD1 port map( A => mult_21_C241_n1274, B => 
                           mult_21_C241_n1300, CI => mult_21_C241_n760, CO => 
                           mult_21_C241_n748, S => mult_21_C241_n749);
   mult_21_C241_U537 : ADFULD1 port map( A => mult_21_C241_n758, B => 
                           mult_21_C241_n753, CI => mult_21_C241_n751, CO => 
                           mult_21_C241_n746, S => mult_21_C241_n747);
   mult_21_C241_U536 : ADFULD1 port map( A => mult_21_C241_n756, B => 
                           mult_21_C241_n749, CI => mult_21_C241_n747, CO => 
                           mult_21_C241_n744, S => mult_21_C241_n745);
   mult_21_C241_U534 : ADFULD1 port map( A => mult_21_C241_n1273, B => 
                           mult_21_C241_n1249, CI => mult_21_C241_n1227, CO => 
                           mult_21_C241_n740, S => mult_21_C241_n741);
   mult_21_C241_U533 : ADFULD1 port map( A => mult_21_C241_n752, B => 
                           mult_21_C241_n1299, CI => mult_21_C241_n743, CO => 
                           mult_21_C241_n738, S => mult_21_C241_n739);
   mult_21_C241_U532 : ADFULD1 port map( A => mult_21_C241_n748, B => 
                           mult_21_C241_n750, CI => mult_21_C241_n741, CO => 
                           mult_21_C241_n736, S => mult_21_C241_n737);
   mult_21_C241_U531 : ADFULD1 port map( A => mult_21_C241_n746, B => 
                           mult_21_C241_n739, CI => mult_21_C241_n737, CO => 
                           mult_21_C241_n734, S => mult_21_C241_n735);
   mult_21_C241_U529 : ADFULD1 port map( A => mult_21_C241_n1248, B => 
                           mult_21_C241_n1356, CI => mult_21_C241_n1326, CO => 
                           mult_21_C241_n730, S => mult_21_C241_n731);
   mult_21_C241_U528 : ADFULD1 port map( A => mult_21_C241_n1272, B => 
                           mult_21_C241_n1298, CI => mult_21_C241_n1226, CO => 
                           mult_21_C241_n728, S => mult_21_C241_n729);
   mult_21_C241_U527 : ADFULD1 port map( A => mult_21_C241_n733, B => 
                           mult_21_C241_n742, CI => mult_21_C241_n740, CO => 
                           mult_21_C241_n726, S => mult_21_C241_n727);
   mult_21_C241_U526 : ADFULD1 port map( A => mult_21_C241_n729, B => 
                           mult_21_C241_n731, CI => mult_21_C241_n738, CO => 
                           mult_21_C241_n724, S => mult_21_C241_n725);
   mult_21_C241_U525 : ADFULD1 port map( A => mult_21_C241_n736, B => 
                           mult_21_C241_n727, CI => mult_21_C241_n725, CO => 
                           mult_21_C241_n722, S => mult_21_C241_n723);
   mult_21_C241_U523 : ADFULD1 port map( A => mult_21_C241_n1271, B => 
                           mult_21_C241_n1297, CI => mult_21_C241_n1225, CO => 
                           mult_21_C241_n718, S => mult_21_C241_n719);
   mult_21_C241_U522 : ADFULD1 port map( A => mult_21_C241_n1205, B => 
                           mult_21_C241_n1247, CI => mult_21_C241_n732, CO => 
                           mult_21_C241_n716, S => mult_21_C241_n717);
   mult_21_C241_U521 : ADFULD1 port map( A => mult_21_C241_n730, B => 
                           mult_21_C241_n721, CI => mult_21_C241_n728, CO => 
                           mult_21_C241_n714, S => mult_21_C241_n715);
   mult_21_C241_U520 : ADFULD1 port map( A => mult_21_C241_n717, B => 
                           mult_21_C241_n719, CI => mult_21_C241_n726, CO => 
                           mult_21_C241_n712, S => mult_21_C241_n713);
   mult_21_C241_U519 : ADFULD1 port map( A => mult_21_C241_n724, B => 
                           mult_21_C241_n715, CI => mult_21_C241_n713, CO => 
                           mult_21_C241_n710, S => mult_21_C241_n711);
   mult_21_C241_U517 : ADFULD1 port map( A => mult_21_C241_n1204, B => 
                           mult_21_C241_n1354, CI => mult_21_C241_n1324, CO => 
                           mult_21_C241_n706, S => mult_21_C241_n707);
   mult_21_C241_U516 : ADFULD1 port map( A => mult_21_C241_n1246, B => 
                           mult_21_C241_n1296, CI => mult_21_C241_n1224, CO => 
                           mult_21_C241_n704, S => mult_21_C241_n705);
   mult_21_C241_U515 : ADFULD1 port map( A => mult_21_C241_n720, B => 
                           mult_21_C241_n1270, CI => mult_21_C241_n709, CO => 
                           mult_21_C241_n702, S => mult_21_C241_n703);
   mult_21_C241_U514 : ADFULD1 port map( A => mult_21_C241_n716, B => 
                           mult_21_C241_n718, CI => mult_21_C241_n707, CO => 
                           mult_21_C241_n700, S => mult_21_C241_n701);
   mult_21_C241_U513 : ADFULD1 port map( A => mult_21_C241_n703, B => 
                           mult_21_C241_n705, CI => mult_21_C241_n714, CO => 
                           mult_21_C241_n698, S => mult_21_C241_n699);
   mult_21_C241_U512 : ADFULD1 port map( A => mult_21_C241_n712, B => 
                           mult_21_C241_n701, CI => mult_21_C241_n699, CO => 
                           mult_21_C241_n696, S => mult_21_C241_n697);
   mult_21_C241_U510 : ADFULD1 port map( A => mult_21_C241_n1295, B => 
                           mult_21_C241_n1269, CI => mult_21_C241_n1223, CO => 
                           mult_21_C241_n692, S => mult_21_C241_n693);
   mult_21_C241_U509 : ADFULD1 port map( A => mult_21_C241_n1185, B => 
                           mult_21_C241_n1245, CI => mult_21_C241_n1203, CO => 
                           mult_21_C241_n690, S => mult_21_C241_n691);
   mult_21_C241_U508 : ADFULD1 port map( A => mult_21_C241_n695, B => 
                           mult_21_C241_n708, CI => mult_21_C241_n706, CO => 
                           mult_21_C241_n688, S => mult_21_C241_n689);
   mult_21_C241_U507 : ADFULD1 port map( A => mult_21_C241_n691, B => 
                           mult_21_C241_n704, CI => mult_21_C241_n693, CO => 
                           mult_21_C241_n686, S => mult_21_C241_n687);
   mult_21_C241_U506 : ADFULD1 port map( A => mult_21_C241_n700, B => 
                           mult_21_C241_n702, CI => mult_21_C241_n689, CO => 
                           mult_21_C241_n684, S => mult_21_C241_n685);
   mult_21_C241_U505 : ADFULD1 port map( A => mult_21_C241_n698, B => 
                           mult_21_C241_n687, CI => mult_21_C241_n685, CO => 
                           mult_21_C241_n682, S => mult_21_C241_n683);
   mult_21_C241_U503 : ADFULD1 port map( A => mult_21_C241_n1202, B => 
                           mult_21_C241_n1352, CI => mult_21_C241_n1322, CO => 
                           mult_21_C241_n678, S => mult_21_C241_n679);
   mult_21_C241_U502 : ADFULD1 port map( A => mult_21_C241_n1184, B => 
                           mult_21_C241_n1268, CI => mult_21_C241_n1222, CO => 
                           mult_21_C241_n676, S => mult_21_C241_n677);
   mult_21_C241_U501 : ADFULD1 port map( A => mult_21_C241_n1244, B => 
                           mult_21_C241_n1294, CI => mult_21_C241_n694, CO => 
                           mult_21_C241_n674, S => mult_21_C241_n675);
   mult_21_C241_U500 : ADFULD1 port map( A => mult_21_C241_n692, B => 
                           mult_21_C241_n681, CI => mult_21_C241_n690, CO => 
                           mult_21_C241_n672, S => mult_21_C241_n673);
   mult_21_C241_U499 : ADFULD1 port map( A => mult_21_C241_n677, B => 
                           mult_21_C241_n679, CI => mult_21_C241_n675, CO => 
                           mult_21_C241_n670, S => mult_21_C241_n671);
   mult_21_C241_U498 : ADFULD1 port map( A => mult_21_C241_n686, B => 
                           mult_21_C241_n688, CI => mult_21_C241_n673, CO => 
                           mult_21_C241_n668, S => mult_21_C241_n669);
   mult_21_C241_U497 : ADFULD1 port map( A => mult_21_C241_n684, B => 
                           mult_21_C241_n671, CI => mult_21_C241_n669, CO => 
                           mult_21_C241_n666, S => mult_21_C241_n667);
   mult_21_C241_U495 : ADFULD1 port map( A => mult_21_C241_n1293, B => 
                           mult_21_C241_n1201, CI => mult_21_C241_n1221, CO => 
                           mult_21_C241_n662, S => mult_21_C241_n663);
   mult_21_C241_U494 : ADFULD1 port map( A => mult_21_C241_n1183, B => 
                           mult_21_C241_n1167, CI => mult_21_C241_n1243, CO => 
                           mult_21_C241_n660, S => mult_21_C241_n661);
   mult_21_C241_U493 : ADFULD1 port map( A => mult_21_C241_n680, B => 
                           mult_21_C241_n1267, CI => mult_21_C241_n665, CO => 
                           mult_21_C241_n658, S => mult_21_C241_n659);
   mult_21_C241_U492 : ADFULD1 port map( A => mult_21_C241_n676, B => 
                           mult_21_C241_n678, CI => mult_21_C241_n674, CO => 
                           mult_21_C241_n656, S => mult_21_C241_n657);
   mult_21_C241_U491 : ADFULD1 port map( A => mult_21_C241_n663, B => 
                           mult_21_C241_n661, CI => mult_21_C241_n672, CO => 
                           mult_21_C241_n654, S => mult_21_C241_n655);
   mult_21_C241_U490 : ADFULD1 port map( A => mult_21_C241_n670, B => 
                           mult_21_C241_n659, CI => mult_21_C241_n657, CO => 
                           mult_21_C241_n652, S => mult_21_C241_n653);
   mult_21_C241_U489 : ADFULD1 port map( A => mult_21_C241_n668, B => 
                           mult_21_C241_n655, CI => mult_21_C241_n653, CO => 
                           mult_21_C241_n650, S => mult_21_C241_n651);
   mult_21_C241_U487 : ADFULD1 port map( A => mult_21_C241_n1200, B => 
                           mult_21_C241_n1350, CI => mult_21_C241_n1320, CO => 
                           mult_21_C241_n646, S => mult_21_C241_n647);
   mult_21_C241_U486 : ADFULD1 port map( A => mult_21_C241_n1166, B => 
                           mult_21_C241_n1266, CI => mult_21_C241_n1220, CO => 
                           mult_21_C241_n644, S => mult_21_C241_n645);
   mult_21_C241_U485 : ADFULD1 port map( A => mult_21_C241_n1182, B => 
                           mult_21_C241_n1292, CI => mult_21_C241_n1242, CO => 
                           mult_21_C241_n642, S => mult_21_C241_n643);
   mult_21_C241_U484 : ADFULD1 port map( A => mult_21_C241_n649, B => 
                           mult_21_C241_n664, CI => mult_21_C241_n662, CO => 
                           mult_21_C241_n640, S => mult_21_C241_n641);
   mult_21_C241_U483 : ADFULD1 port map( A => mult_21_C241_n647, B => 
                           mult_21_C241_n660, CI => mult_21_C241_n643, CO => 
                           mult_21_C241_n638, S => mult_21_C241_n639);
   mult_21_C241_U482 : ADFULD1 port map( A => mult_21_C241_n658, B => 
                           mult_21_C241_n645, CI => mult_21_C241_n656, CO => 
                           mult_21_C241_n636, S => mult_21_C241_n637);
   mult_21_C241_U481 : ADFULD1 port map( A => mult_21_C241_n639, B => 
                           mult_21_C241_n641, CI => mult_21_C241_n654, CO => 
                           mult_21_C241_n634, S => mult_21_C241_n635);
   mult_21_C241_U480 : ADFULD1 port map( A => mult_21_C241_n652, B => 
                           mult_21_C241_n637, CI => mult_21_C241_n635, CO => 
                           mult_21_C241_n632, S => mult_21_C241_n633);
   mult_21_C241_U478 : ADFULD1 port map( A => mult_21_C241_n1151, B => 
                           mult_21_C241_n1199, CI => mult_21_C241_n1219, CO => 
                           mult_21_C241_n628, S => mult_21_C241_n629);
   mult_21_C241_U477 : ADFULD1 port map( A => mult_21_C241_n1291, B => 
                           mult_21_C241_n1181, CI => mult_21_C241_n1165, CO => 
                           mult_21_C241_n626, S => mult_21_C241_n627);
   mult_21_C241_U476 : ADFULD1 port map( A => mult_21_C241_n1241, B => 
                           mult_21_C241_n1265, CI => mult_21_C241_n648, CO => 
                           mult_21_C241_n624, S => mult_21_C241_n625);
   mult_21_C241_U475 : ADFULD1 port map( A => mult_21_C241_n646, B => 
                           mult_21_C241_n631, CI => mult_21_C241_n642, CO => 
                           mult_21_C241_n622, S => mult_21_C241_n623);
   mult_21_C241_U474 : ADFULD1 port map( A => mult_21_C241_n627, B => 
                           mult_21_C241_n644, CI => mult_21_C241_n629, CO => 
                           mult_21_C241_n620, S => mult_21_C241_n621);
   mult_21_C241_U473 : ADFULD1 port map( A => mult_21_C241_n640, B => 
                           mult_21_C241_n625, CI => mult_21_C241_n638, CO => 
                           mult_21_C241_n618, S => mult_21_C241_n619);
   mult_21_C241_U472 : ADFULD1 port map( A => mult_21_C241_n621, B => 
                           mult_21_C241_n623, CI => mult_21_C241_n636, CO => 
                           mult_21_C241_n616, S => mult_21_C241_n617);
   mult_21_C241_U471 : ADFULD1 port map( A => mult_21_C241_n634, B => 
                           mult_21_C241_n619, CI => mult_21_C241_n617, CO => 
                           mult_21_C241_n614, S => mult_21_C241_n615);
   mult_21_C241_U469 : ADFULD1 port map( A => mult_21_C241_n1164, B => 
                           mult_21_C241_n1348, CI => mult_21_C241_n1318, CO => 
                           mult_21_C241_n610, S => mult_21_C241_n611);
   mult_21_C241_U468 : ADFULD1 port map( A => mult_21_C241_n1290, B => 
                           mult_21_C241_n1198, CI => mult_21_C241_n1218, CO => 
                           mult_21_C241_n608, S => mult_21_C241_n609);
   mult_21_C241_U467 : ADFULD1 port map( A => mult_21_C241_n1150, B => 
                           mult_21_C241_n1264, CI => mult_21_C241_n1180, CO => 
                           mult_21_C241_n606, S => mult_21_C241_n607);
   mult_21_C241_U466 : ADFULD1 port map( A => mult_21_C241_n630, B => 
                           mult_21_C241_n1240, CI => mult_21_C241_n613, CO => 
                           mult_21_C241_n604, S => mult_21_C241_n605);
   mult_21_C241_U465 : ADFULD1 port map( A => mult_21_C241_n626, B => 
                           mult_21_C241_n628, CI => mult_21_C241_n624, CO => 
                           mult_21_C241_n602, S => mult_21_C241_n603);
   mult_21_C241_U464 : ADFULD1 port map( A => mult_21_C241_n609, B => 
                           mult_21_C241_n611, CI => mult_21_C241_n607, CO => 
                           mult_21_C241_n600, S => mult_21_C241_n601);
   mult_21_C241_U463 : ADFULD1 port map( A => mult_21_C241_n622, B => 
                           mult_21_C241_n605, CI => mult_21_C241_n620, CO => 
                           mult_21_C241_n598, S => mult_21_C241_n599);
   mult_21_C241_U462 : ADFULD1 port map( A => mult_21_C241_n601, B => 
                           mult_21_C241_n603, CI => mult_21_C241_n618, CO => 
                           mult_21_C241_n596, S => mult_21_C241_n597);
   mult_21_C241_U461 : ADFULD1 port map( A => mult_21_C241_n616, B => 
                           mult_21_C241_n599, CI => mult_21_C241_n597, CO => 
                           mult_21_C241_n594, S => mult_21_C241_n595);
   mult_21_C241_U459 : ADFULD1 port map( A => mult_21_C241_n1289, B => 
                           mult_21_C241_n1179, CI => mult_21_C241_n1217, CO => 
                           mult_21_C241_n590, S => mult_21_C241_n591);
   mult_21_C241_U458 : ADFULD1 port map( A => mult_21_C241_n1263, B => 
                           mult_21_C241_n1149, CI => mult_21_C241_n1137, CO => 
                           mult_21_C241_n588, S => mult_21_C241_n589);
   mult_21_C241_U457 : ADFULD1 port map( A => mult_21_C241_n1163, B => 
                           mult_21_C241_n1239, CI => mult_21_C241_n1197, CO => 
                           mult_21_C241_n586, S => mult_21_C241_n587);
   mult_21_C241_U456 : ADFULD1 port map( A => mult_21_C241_n593, B => 
                           mult_21_C241_n612, CI => mult_21_C241_n610, CO => 
                           mult_21_C241_n584, S => mult_21_C241_n585);
   mult_21_C241_U455 : ADFULD1 port map( A => mult_21_C241_n606, B => 
                           mult_21_C241_n608, CI => mult_21_C241_n587, CO => 
                           mult_21_C241_n582, S => mult_21_C241_n583);
   mult_21_C241_U454 : ADFULD1 port map( A => mult_21_C241_n591, B => 
                           mult_21_C241_n589, CI => mult_21_C241_n604, CO => 
                           mult_21_C241_n580, S => mult_21_C241_n581);
   mult_21_C241_U453 : ADFULD1 port map( A => mult_21_C241_n585, B => 
                           mult_21_C241_n602, CI => mult_21_C241_n600, CO => 
                           mult_21_C241_n578, S => mult_21_C241_n579);
   mult_21_C241_U452 : ADFULD1 port map( A => mult_21_C241_n581, B => 
                           mult_21_C241_n583, CI => mult_21_C241_n598, CO => 
                           mult_21_C241_n576, S => mult_21_C241_n577);
   mult_21_C241_U451 : ADFULD1 port map( A => mult_21_C241_n596, B => 
                           mult_21_C241_n579, CI => mult_21_C241_n577, CO => 
                           mult_21_C241_n574, S => mult_21_C241_n575);
   mult_21_C241_U449 : ADFULD1 port map( A => mult_21_C241_n1136, B => 
                           mult_21_C241_n1346, CI => mult_21_C241_n1316, CO => 
                           mult_21_C241_n570, S => mult_21_C241_n571);
   mult_21_C241_U448 : ADFULD1 port map( A => mult_21_C241_n1288, B => 
                           mult_21_C241_n1178, CI => mult_21_C241_n1216, CO => 
                           mult_21_C241_n568, S => mult_21_C241_n569);
   mult_21_C241_U447 : ADFULD1 port map( A => mult_21_C241_n1148, B => 
                           mult_21_C241_n1262, CI => mult_21_C241_n1162, CO => 
                           mult_21_C241_n566, S => mult_21_C241_n567);
   mult_21_C241_U446 : ADFULD1 port map( A => mult_21_C241_n1196, B => 
                           mult_21_C241_n1238, CI => mult_21_C241_n592, CO => 
                           mult_21_C241_n564, S => mult_21_C241_n565);
   mult_21_C241_U445 : ADFULD1 port map( A => mult_21_C241_n590, B => 
                           mult_21_C241_n573, CI => mult_21_C241_n588, CO => 
                           mult_21_C241_n562, S => mult_21_C241_n563);
   mult_21_C241_U444 : ADFULD1 port map( A => mult_21_C241_n571, B => 
                           mult_21_C241_n586, CI => mult_21_C241_n567, CO => 
                           mult_21_C241_n560, S => mult_21_C241_n561);
   mult_21_C241_U443 : ADFULD1 port map( A => mult_21_C241_n565, B => 
                           mult_21_C241_n569, CI => mult_21_C241_n584, CO => 
                           mult_21_C241_n558, S => mult_21_C241_n559);
   mult_21_C241_U442 : ADFULD1 port map( A => mult_21_C241_n563, B => 
                           mult_21_C241_n582, CI => mult_21_C241_n580, CO => 
                           mult_21_C241_n556, S => mult_21_C241_n557);
   mult_21_C241_U441 : ADFULD1 port map( A => mult_21_C241_n559, B => 
                           mult_21_C241_n561, CI => mult_21_C241_n578, CO => 
                           mult_21_C241_n554, S => mult_21_C241_n555);
   mult_21_C241_U440 : ADFULD1 port map( A => mult_21_C241_n576, B => 
                           mult_21_C241_n557, CI => mult_21_C241_n555, CO => 
                           mult_21_C241_n552, S => mult_21_C241_n553);
   mult_21_C241_U438 : ADFULD1 port map( A => mult_21_C241_n1125, B => 
                           mult_21_C241_n1177, CI => mult_21_C241_n1215, CO => 
                           mult_21_C241_n548, S => mult_21_C241_n549);
   mult_21_C241_U437 : ADFULD1 port map( A => mult_21_C241_n1287, B => 
                           mult_21_C241_n1161, CI => mult_21_C241_n1261, CO => 
                           mult_21_C241_n546, S => mult_21_C241_n547);
   mult_21_C241_U436 : ADFULD1 port map( A => mult_21_C241_n1135, B => 
                           mult_21_C241_n1237, CI => mult_21_C241_n1147, CO => 
                           mult_21_C241_n544, S => mult_21_C241_n545);
   mult_21_C241_U435 : ADFULD1 port map( A => mult_21_C241_n572, B => 
                           mult_21_C241_n1195, CI => mult_21_C241_n551, CO => 
                           mult_21_C241_n542, S => mult_21_C241_n543);
   mult_21_C241_U434 : ADFULD1 port map( A => mult_21_C241_n566, B => 
                           mult_21_C241_n570, CI => mult_21_C241_n568, CO => 
                           mult_21_C241_n540, S => mult_21_C241_n541);
   mult_21_C241_U433 : ADFULD1 port map( A => mult_21_C241_n549, B => 
                           mult_21_C241_n564, CI => mult_21_C241_n547, CO => 
                           mult_21_C241_n538, S => mult_21_C241_n539);
   mult_21_C241_U432 : ADFULD1 port map( A => mult_21_C241_n562, B => 
                           mult_21_C241_n545, CI => mult_21_C241_n543, CO => 
                           mult_21_C241_n536, S => mult_21_C241_n537);
   mult_21_C241_U431 : ADFULD1 port map( A => mult_21_C241_n541, B => 
                           mult_21_C241_n560, CI => mult_21_C241_n558, CO => 
                           mult_21_C241_n534, S => mult_21_C241_n535);
   mult_21_C241_U430 : ADFULD1 port map( A => mult_21_C241_n556, B => 
                           mult_21_C241_n539, CI => mult_21_C241_n537, CO => 
                           mult_21_C241_n532, S => mult_21_C241_n533);
   mult_21_C241_U429 : ADFULD1 port map( A => mult_21_C241_n554, B => 
                           mult_21_C241_n535, CI => mult_21_C241_n533, CO => 
                           mult_21_C241_n530, S => mult_21_C241_n531);
   mult_21_C241_U427 : ADFULD1 port map( A => mult_21_C241_n1146, B => 
                           mult_21_C241_n1344, CI => mult_21_C241_n1314, CO => 
                           mult_21_C241_n526, S => mult_21_C241_n527);
   mult_21_C241_U426 : ADFULD1 port map( A => mult_21_C241_n1124, B => 
                           mult_21_C241_n1176, CI => mult_21_C241_n1214, CO => 
                           mult_21_C241_n524, S => mult_21_C241_n525);
   mult_21_C241_U425 : ADFULD1 port map( A => mult_21_C241_n1134, B => 
                           mult_21_C241_n1286, CI => mult_21_C241_n1160, CO => 
                           mult_21_C241_n522, S => mult_21_C241_n523);
   mult_21_C241_U424 : ADFULD1 port map( A => mult_21_C241_n1194, B => 
                           mult_21_C241_n1260, CI => mult_21_C241_n1236, CO => 
                           mult_21_C241_n520, S => mult_21_C241_n521);
   mult_21_C241_U423 : ADFULD1 port map( A => mult_21_C241_n529, B => 
                           mult_21_C241_n550, CI => mult_21_C241_n548, CO => 
                           mult_21_C241_n518, S => mult_21_C241_n519);
   mult_21_C241_U422 : ADFULD1 port map( A => mult_21_C241_n544, B => 
                           mult_21_C241_n546, CI => mult_21_C241_n527, CO => 
                           mult_21_C241_n516, S => mult_21_C241_n517);
   mult_21_C241_U421 : ADFULD1 port map( A => mult_21_C241_n525, B => 
                           mult_21_C241_n521, CI => mult_21_C241_n523, CO => 
                           mult_21_C241_n514, S => mult_21_C241_n515);
   mult_21_C241_U420 : ADFULD1 port map( A => mult_21_C241_n540, B => 
                           mult_21_C241_n542, CI => mult_21_C241_n519, CO => 
                           mult_21_C241_n512, S => mult_21_C241_n513);
   mult_21_C241_U419 : ADFULD1 port map( A => mult_21_C241_n517, B => 
                           mult_21_C241_n538, CI => mult_21_C241_n515, CO => 
                           mult_21_C241_n510, S => mult_21_C241_n511);
   mult_21_C241_U418 : ADFULD1 port map( A => mult_21_C241_n513, B => 
                           mult_21_C241_n536, CI => mult_21_C241_n534, CO => 
                           mult_21_C241_n508, S => mult_21_C241_n509);
   mult_21_C241_U417 : ADFULD1 port map( A => mult_21_C241_n532, B => 
                           mult_21_C241_n511, CI => mult_21_C241_n509, CO => 
                           mult_21_C241_n506, S => mult_21_C241_n507);
   mult_21_C241_U415 : ADFULD1 port map( A => mult_21_C241_n1115, B => 
                           mult_21_C241_n1175, CI => mult_21_C241_n1213, CO => 
                           mult_21_C241_n502, S => mult_21_C241_n503);
   mult_21_C241_U414 : ADFULD1 port map( A => mult_21_C241_n1123, B => 
                           mult_21_C241_n1145, CI => mult_21_C241_n1133, CO => 
                           mult_21_C241_n500, S => mult_21_C241_n501);
   mult_21_C241_U413 : ADFULD1 port map( A => mult_21_C241_n1159, B => 
                           mult_21_C241_n1285, CI => mult_21_C241_n1193, CO => 
                           mult_21_C241_n498, S => mult_21_C241_n499);
   mult_21_C241_U412 : ADFULD1 port map( A => mult_21_C241_n1235, B => 
                           mult_21_C241_n1259, CI => mult_21_C241_n528, CO => 
                           mult_21_C241_n496, S => mult_21_C241_n497);
   mult_21_C241_U411 : ADFULD1 port map( A => mult_21_C241_n526, B => 
                           mult_21_C241_n505, CI => mult_21_C241_n520, CO => 
                           mult_21_C241_n494, S => mult_21_C241_n495);
   mult_21_C241_U410 : ADFULD1 port map( A => mult_21_C241_n522, B => 
                           mult_21_C241_n524, CI => mult_21_C241_n499, CO => 
                           mult_21_C241_n492, S => mult_21_C241_n493);
   mult_21_C241_U409 : ADFULD1 port map( A => mult_21_C241_n501, B => 
                           mult_21_C241_n503, CI => mult_21_C241_n497, CO => 
                           mult_21_C241_n490, S => mult_21_C241_n491);
   mult_21_C241_U408 : ADFULD1 port map( A => mult_21_C241_n516, B => 
                           mult_21_C241_n518, CI => mult_21_C241_n495, CO => 
                           mult_21_C241_n488, S => mult_21_C241_n489);
   mult_21_C241_U407 : ADFULD1 port map( A => mult_21_C241_n493, B => 
                           mult_21_C241_n514, CI => mult_21_C241_n491, CO => 
                           mult_21_C241_n486, S => mult_21_C241_n487);
   mult_21_C241_U406 : ADFULD1 port map( A => mult_21_C241_n510, B => 
                           mult_21_C241_n512, CI => mult_21_C241_n489, CO => 
                           mult_21_C241_n484, S => mult_21_C241_n485);
   mult_21_C241_U405 : ADFULD1 port map( A => mult_21_C241_n508, B => 
                           mult_21_C241_n487, CI => mult_21_C241_n485, CO => 
                           mult_21_C241_n482, S => mult_21_C241_n483);
   mult_21_C241_U403 : ADFULD1 port map( A => mult_21_C241_n1114, B => 
                           mult_21_C241_n1342, CI => mult_21_C241_n1312, CO => 
                           mult_21_C241_n478, S => mult_21_C241_n479);
   mult_21_C241_U402 : ADFULD1 port map( A => mult_21_C241_n1284, B => 
                           mult_21_C241_n1174, CI => mult_21_C241_n1212, CO => 
                           mult_21_C241_n476, S => mult_21_C241_n477);
   mult_21_C241_U401 : ADFULD1 port map( A => mult_21_C241_n1258, B => 
                           mult_21_C241_n1132, CI => mult_21_C241_n1122, CO => 
                           mult_21_C241_n474, S => mult_21_C241_n475);
   mult_21_C241_U400 : ADFULD1 port map( A => mult_21_C241_n1144, B => 
                           mult_21_C241_n1234, CI => mult_21_C241_n1158, CO => 
                           mult_21_C241_n472, S => mult_21_C241_n473);
   mult_21_C241_U399 : ADFULD1 port map( A => mult_21_C241_n504, B => 
                           mult_21_C241_n1192, CI => mult_21_C241_n481, CO => 
                           mult_21_C241_n470, S => mult_21_C241_n471);
   mult_21_C241_U398 : ADFULD1 port map( A => mult_21_C241_n498, B => 
                           mult_21_C241_n502, CI => mult_21_C241_n496, CO => 
                           mult_21_C241_n468, S => mult_21_C241_n469);
   mult_21_C241_U397 : ADFULD1 port map( A => mult_21_C241_n479, B => 
                           mult_21_C241_n500, CI => mult_21_C241_n473, CO => 
                           mult_21_C241_n466, S => mult_21_C241_n467);
   mult_21_C241_U396 : ADFULD1 port map( A => mult_21_C241_n475, B => 
                           mult_21_C241_n477, CI => mult_21_C241_n471, CO => 
                           mult_21_C241_n464, S => mult_21_C241_n465);
   mult_21_C241_U395 : ADFULD1 port map( A => mult_21_C241_n492, B => 
                           mult_21_C241_n494, CI => mult_21_C241_n490, CO => 
                           mult_21_C241_n462, S => mult_21_C241_n463);
   mult_21_C241_U394 : ADFULD1 port map( A => mult_21_C241_n467, B => 
                           mult_21_C241_n469, CI => mult_21_C241_n465, CO => 
                           mult_21_C241_n460, S => mult_21_C241_n461);
   mult_21_C241_U393 : ADFULD1 port map( A => mult_21_C241_n486, B => 
                           mult_21_C241_n488, CI => mult_21_C241_n463, CO => 
                           mult_21_C241_n458, S => mult_21_C241_n459);
   mult_21_C241_U392 : ADFULD1 port map( A => mult_21_C241_n484, B => 
                           mult_21_C241_n461, CI => mult_21_C241_n459, CO => 
                           mult_21_C241_n456, S => mult_21_C241_n457);
   mult_21_C241_U390 : ADFULD1 port map( A => mult_21_C241_n1107, B => 
                           mult_21_C241_n1157, CI => mult_21_C241_n1211, CO => 
                           mult_21_C241_n452, S => mult_21_C241_n453);
   mult_21_C241_U389 : ADFULD1 port map( A => mult_21_C241_n1283, B => 
                           mult_21_C241_n1143, CI => mult_21_C241_n1257, CO => 
                           mult_21_C241_n450, S => mult_21_C241_n451);
   mult_21_C241_U388 : ADFULD1 port map( A => mult_21_C241_n1113, B => 
                           mult_21_C241_n1233, CI => mult_21_C241_n1121, CO => 
                           mult_21_C241_n448, S => mult_21_C241_n449);
   mult_21_C241_U387 : ADFULD1 port map( A => mult_21_C241_n1131, B => 
                           mult_21_C241_n1191, CI => mult_21_C241_n1173, CO => 
                           mult_21_C241_n446, S => mult_21_C241_n447);
   mult_21_C241_U386 : ADFULD1 port map( A => mult_21_C241_n455, B => 
                           mult_21_C241_n480, CI => mult_21_C241_n478, CO => 
                           mult_21_C241_n444, S => mult_21_C241_n445);
   mult_21_C241_U385 : ADFULD1 port map( A => mult_21_C241_n474, B => 
                           mult_21_C241_n472, CI => mult_21_C241_n476, CO => 
                           mult_21_C241_n442, S => mult_21_C241_n443);
   mult_21_C241_U384 : ADFULD1 port map( A => mult_21_C241_n453, B => 
                           mult_21_C241_n447, CI => mult_21_C241_n470, CO => 
                           mult_21_C241_n440, S => mult_21_C241_n441);
   mult_21_C241_U383 : ADFULD1 port map( A => mult_21_C241_n449, B => 
                           mult_21_C241_n451, CI => mult_21_C241_n468, CO => 
                           mult_21_C241_n438, S => mult_21_C241_n439);
   mult_21_C241_U382 : ADFULD1 port map( A => mult_21_C241_n466, B => 
                           mult_21_C241_n445, CI => mult_21_C241_n443, CO => 
                           mult_21_C241_n436, S => mult_21_C241_n437);
   mult_21_C241_U381 : ADFULD1 port map( A => mult_21_C241_n441, B => 
                           mult_21_C241_n464, CI => mult_21_C241_n462, CO => 
                           mult_21_C241_n434, S => mult_21_C241_n435);
   mult_21_C241_U380 : ADFULD1 port map( A => mult_21_C241_n437, B => 
                           mult_21_C241_n439, CI => mult_21_C241_n460, CO => 
                           mult_21_C241_n432, S => mult_21_C241_n433);
   mult_21_C241_U379 : ADFULD1 port map( A => mult_21_C241_n458, B => 
                           mult_21_C241_n435, CI => mult_21_C241_n433, CO => 
                           mult_21_C241_n430, S => mult_21_C241_n431);
   mult_21_C241_U377 : ADFULD1 port map( A => mult_21_C241_n1106, B => 
                           mult_21_C241_n1340, CI => mult_21_C241_n1310, CO => 
                           mult_21_C241_n426, S => mult_21_C241_n427);
   mult_21_C241_U376 : ADFULD1 port map( A => mult_21_C241_n1282, B => 
                           mult_21_C241_n1156, CI => mult_21_C241_n1210, CO => 
                           mult_21_C241_n424, S => mult_21_C241_n425);
   mult_21_C241_U375 : ADFULD1 port map( A => mult_21_C241_n1112, B => 
                           mult_21_C241_n1130, CI => mult_21_C241_n1120, CO => 
                           mult_21_C241_n422, S => mult_21_C241_n423);
   mult_21_C241_U374 : ADFULD1 port map( A => mult_21_C241_n1142, B => 
                           mult_21_C241_n1256, CI => mult_21_C241_n1172, CO => 
                           mult_21_C241_n420, S => mult_21_C241_n421);
   mult_21_C241_U373 : ADFULD1 port map( A => mult_21_C241_n1232, B => 
                           mult_21_C241_n1190, CI => mult_21_C241_n454, CO => 
                           mult_21_C241_n418, S => mult_21_C241_n419);
   mult_21_C241_U372 : ADFULD1 port map( A => mult_21_C241_n452, B => 
                           mult_21_C241_n429, CI => mult_21_C241_n450, CO => 
                           mult_21_C241_n416, S => mult_21_C241_n417);
   mult_21_C241_U371 : ADFULD1 port map( A => mult_21_C241_n448, B => 
                           mult_21_C241_n446, CI => mult_21_C241_n427, CO => 
                           mult_21_C241_n414, S => mult_21_C241_n415);
   mult_21_C241_U370 : ADFULD1 port map( A => mult_21_C241_n421, B => 
                           mult_21_C241_n423, CI => mult_21_C241_n425, CO => 
                           mult_21_C241_n412, S => mult_21_C241_n413);
   mult_21_C241_U369 : ADFULD1 port map( A => mult_21_C241_n444, B => 
                           mult_21_C241_n419, CI => mult_21_C241_n442, CO => 
                           mult_21_C241_n410, S => mult_21_C241_n411);
   mult_21_C241_U368 : ADFULD1 port map( A => mult_21_C241_n440, B => 
                           mult_21_C241_n417, CI => mult_21_C241_n415, CO => 
                           mult_21_C241_n408, S => mult_21_C241_n409);
   mult_21_C241_U367 : ADFULD1 port map( A => mult_21_C241_n438, B => 
                           mult_21_C241_n413, CI => mult_21_C241_n411, CO => 
                           mult_21_C241_n406, S => mult_21_C241_n407);
   mult_21_C241_U366 : ADFULD1 port map( A => mult_21_C241_n409, B => 
                           mult_21_C241_n436, CI => mult_21_C241_n434, CO => 
                           mult_21_C241_n404, S => mult_21_C241_n405);
   mult_21_C241_U365 : ADFULD1 port map( A => mult_21_C241_n432, B => 
                           mult_21_C241_n407, CI => mult_21_C241_n405, CO => 
                           mult_21_C241_n402, S => mult_21_C241_n403);
   mult_21_C241_U363 : ADFULD1 port map( A => mult_21_C241_n1281, B => 
                           mult_21_C241_n1155, CI => mult_21_C241_n1209, CO => 
                           mult_21_C241_n398, S => mult_21_C241_n399);
   mult_21_C241_U362 : ADFULD1 port map( A => mult_21_C241_n1255, B => 
                           mult_21_C241_n1119, CI => mult_21_C241_n1101, CO => 
                           mult_21_C241_n396, S => mult_21_C241_n397);
   mult_21_C241_U361 : ADFULD1 port map( A => mult_21_C241_n1231, B => 
                           mult_21_C241_n1111, CI => mult_21_C241_n1105, CO => 
                           mult_21_C241_n394, S => mult_21_C241_n395);
   mult_21_C241_U360 : ADFULD1 port map( A => mult_21_C241_n1129, B => 
                           mult_21_C241_n1189, CI => mult_21_C241_n1141, CO => 
                           mult_21_C241_n392, S => mult_21_C241_n393);
   mult_21_C241_U359 : ADFULD1 port map( A => mult_21_C241_n428, B => 
                           mult_21_C241_n1171, CI => mult_21_C241_n401, CO => 
                           mult_21_C241_n390, S => mult_21_C241_n391);
   mult_21_C241_U358 : ADFULD1 port map( A => mult_21_C241_n424, B => 
                           mult_21_C241_n426, CI => mult_21_C241_n420, CO => 
                           mult_21_C241_n388, S => mult_21_C241_n389);
   mult_21_C241_U357 : ADFULD1 port map( A => mult_21_C241_n418, B => 
                           mult_21_C241_n422, CI => mult_21_C241_n393, CO => 
                           mult_21_C241_n386, S => mult_21_C241_n387);
   mult_21_C241_U356 : ADFULD1 port map( A => mult_21_C241_n395, B => 
                           mult_21_C241_n397, CI => mult_21_C241_n399, CO => 
                           mult_21_C241_n384, S => mult_21_C241_n385);
   mult_21_C241_U355 : ADFULD1 port map( A => mult_21_C241_n391, B => 
                           mult_21_C241_n416, CI => mult_21_C241_n414, CO => 
                           mult_21_C241_n382, S => mult_21_C241_n383);
   mult_21_C241_U354 : ADFULD1 port map( A => mult_21_C241_n412, B => 
                           mult_21_C241_n389, CI => mult_21_C241_n387, CO => 
                           mult_21_C241_n380, S => mult_21_C241_n381);
   mult_21_C241_U353 : ADFULD1 port map( A => mult_21_C241_n410, B => 
                           mult_21_C241_n385, CI => mult_21_C241_n383, CO => 
                           mult_21_C241_n378, S => mult_21_C241_n379);
   mult_21_C241_U352 : ADFULD1 port map( A => mult_21_C241_n381, B => 
                           mult_21_C241_n408, CI => mult_21_C241_n406, CO => 
                           mult_21_C241_n376, S => mult_21_C241_n377);
   mult_21_C241_U351 : ADFULD1 port map( A => mult_21_C241_n404, B => 
                           mult_21_C241_n379, CI => mult_21_C241_n377, CO => 
                           mult_21_C241_n374, S => mult_21_C241_n375);
   mult_21_C241_U349 : ADFULD1 port map( A => mult_21_C241_n1100, B => 
                           mult_21_C241_n1338, CI => mult_21_C241_n1308, CO => 
                           mult_21_C241_n370, S => mult_21_C241_n371);
   mult_21_C241_U348 : ADFULD1 port map( A => mult_21_C241_n1280, B => 
                           mult_21_C241_n1154, CI => mult_21_C241_n1208, CO => 
                           mult_21_C241_n368, S => mult_21_C241_n369);
   mult_21_C241_U347 : ADFULD1 port map( A => mult_21_C241_n1254, B => 
                           mult_21_C241_n1128, CI => mult_21_C241_n1230, CO => 
                           mult_21_C241_n366, S => mult_21_C241_n367);
   mult_21_C241_U346 : ADFULD1 port map( A => mult_21_C241_n1104, B => 
                           mult_21_C241_n1188, CI => mult_21_C241_n1110, CO => 
                           mult_21_C241_n364, S => mult_21_C241_n365);
   mult_21_C241_U345 : ADFULD1 port map( A => mult_21_C241_n1170, B => 
                           mult_21_C241_n1118, CI => mult_21_C241_n1140, CO => 
                           mult_21_C241_n362, S => mult_21_C241_n363);
   mult_21_C241_U344 : ADFULD1 port map( A => mult_21_C241_n373, B => 
                           mult_21_C241_n400, CI => mult_21_C241_n392, CO => 
                           mult_21_C241_n360, S => mult_21_C241_n361);
   mult_21_C241_U343 : ADFULD1 port map( A => mult_21_C241_n398, B => 
                           mult_21_C241_n394, CI => mult_21_C241_n396, CO => 
                           mult_21_C241_n358, S => mult_21_C241_n359);
   mult_21_C241_U342 : ADFULD1 port map( A => mult_21_C241_n369, B => 
                           mult_21_C241_n371, CI => mult_21_C241_n367, CO => 
                           mult_21_C241_n356, S => mult_21_C241_n357);
   mult_21_C241_U341 : ADFULD1 port map( A => mult_21_C241_n365, B => 
                           mult_21_C241_n363, CI => mult_21_C241_n390, CO => 
                           mult_21_C241_n354, S => mult_21_C241_n355);
   mult_21_C241_U340 : ADFULD1 port map( A => mult_21_C241_n361, B => 
                           mult_21_C241_n388, CI => mult_21_C241_n386, CO => 
                           mult_21_C241_n352, S => mult_21_C241_n353);
   mult_21_C241_U339 : ADFULD1 port map( A => mult_21_C241_n359, B => 
                           mult_21_C241_n384, CI => mult_21_C241_n357, CO => 
                           mult_21_C241_n350, S => mult_21_C241_n351);
   mult_21_C241_U338 : ADFULD1 port map( A => mult_21_C241_n382, B => 
                           mult_21_C241_n355, CI => mult_21_C241_n380, CO => 
                           mult_21_C241_n348, S => mult_21_C241_n349);
   mult_21_C241_U337 : ADFULD1 port map( A => mult_21_C241_n351, B => 
                           mult_21_C241_n353, CI => mult_21_C241_n378, CO => 
                           mult_21_C241_n346, S => mult_21_C241_n347);
   mult_21_C241_U336 : ADFULD1 port map( A => mult_21_C241_n376, B => 
                           mult_21_C241_n349, CI => mult_21_C241_n347, CO => 
                           mult_21_C241_n344, S => mult_21_C241_n345);
   mult_21_C241_U334 : EXOR3D1 port map( A1 => mult_21_C241_n1097, A2 => 
                           mult_21_C241_n1279, A3 => mult_21_C241_n1207, Z => 
                           mult_21_C241_n342);
   mult_21_C241_U333 : EXOR3D1 port map( A1 => mult_21_C241_n1253, A2 => 
                           mult_21_C241_n1127, A3 => mult_21_C241_n1099, Z => 
                           mult_21_C241_n341);
   mult_21_C241_U332 : EXOR3D1 port map( A1 => mult_21_C241_n1103, A2 => 
                           mult_21_C241_n1117, A3 => mult_21_C241_n1109, Z => 
                           mult_21_C241_n340);
   mult_21_C241_U331 : EXOR3D1 port map( A1 => mult_21_C241_n1139, A2 => 
                           mult_21_C241_n1229, A3 => mult_21_C241_n1153, Z => 
                           mult_21_C241_n339);
   mult_21_C241_U330 : EXOR3D1 port map( A1 => mult_21_C241_n1187, A2 => 
                           mult_21_C241_n1169, A3 => mult_21_C241_n372, Z => 
                           mult_21_C241_n338);
   mult_21_C241_U329 : EXOR3D1 port map( A1 => mult_21_C241_n368, A2 => 
                           mult_21_C241_n370, A3 => mult_21_C241_n364, Z => 
                           mult_21_C241_n337);
   mult_21_C241_U328 : EXOR3D1 port map( A1 => mult_21_C241_n366, A2 => 
                           mult_21_C241_n343, A3 => mult_21_C241_n362, Z => 
                           mult_21_C241_n336);
   mult_21_C241_U327 : EXOR3D1 port map( A1 => mult_21_C241_n342, A2 => 
                           mult_21_C241_n338, A3 => mult_21_C241_n341, Z => 
                           mult_21_C241_n335);
   mult_21_C241_U326 : EXOR3D1 port map( A1 => mult_21_C241_n339, A2 => 
                           mult_21_C241_n340, A3 => mult_21_C241_n360, Z => 
                           mult_21_C241_n334);
   mult_21_C241_U325 : EXOR3D1 port map( A1 => mult_21_C241_n337, A2 => 
                           mult_21_C241_n358, A3 => mult_21_C241_n336, Z => 
                           mult_21_C241_n333);
   mult_21_C241_U324 : EXOR3D1 port map( A1 => mult_21_C241_n354, A2 => 
                           mult_21_C241_n356, A3 => mult_21_C241_n335, Z => 
                           mult_21_C241_n332);
   mult_21_C241_U323 : EXOR3D1 port map( A1 => mult_21_C241_n352, A2 => 
                           mult_21_C241_n334, A3 => mult_21_C241_n333, Z => 
                           mult_21_C241_n331);
   mult_21_C241_U322 : EXOR3D1 port map( A1 => mult_21_C241_n332, A2 => 
                           mult_21_C241_n350, A3 => mult_21_C241_n348, Z => 
                           mult_21_C241_n330);
   mult_21_C241_U321 : EXOR3D1 port map( A1 => mult_21_C241_n346, A2 => 
                           mult_21_C241_n331, A3 => mult_21_C241_n330, Z => 
                           mult_21_C241_n329);
   mult_21_C241_U313 : EXOR2D1 port map( A1 => mult_21_C241_n303, A2 => 
                           mult_21_C241_n305, Z => N3234);
   mult_21_C241_U305 : EXNOR2D1 port map( A1 => mult_21_C241_n176, A2 => 
                           mult_21_C241_n302, Z => N3235);
   mult_21_C241_U300 : OAI21D1 port map( A1 => mult_21_C241_n297, A2 => 
                           mult_21_C241_n295, B => mult_21_C241_n296, Z => 
                           mult_21_C241_n294);
   mult_21_C241_U299 : EXOR2D1 port map( A1 => mult_21_C241_n297, A2 => 
                           mult_21_C241_n175, Z => N3236);
   mult_21_C241_U291 : EXNOR2D1 port map( A1 => mult_21_C241_n174, A2 => 
                           mult_21_C241_n294, Z => N3237);
   mult_21_C241_U286 : OAI21D1 port map( A1 => mult_21_C241_n289, A2 => 
                           mult_21_C241_n287, B => mult_21_C241_n288, Z => 
                           mult_21_C241_n286);
   mult_21_C241_U284 : EXOR2D1 port map( A1 => mult_21_C241_n173, A2 => 
                           mult_21_C241_n289, Z => N3238);
   mult_21_C241_U279 : OAI21D1 port map( A1 => mult_21_C241_n285, A2 => 
                           mult_21_C241_n283, B => mult_21_C241_n284, Z => 
                           mult_21_C241_n282);
   mult_21_C241_U278 : EXOR2D1 port map( A1 => mult_21_C241_n172, A2 => 
                           mult_21_C241_n285, Z => N3239);
   mult_21_C241_U273 : OAI21D1 port map( A1 => mult_21_C241_n280, A2 => 
                           mult_21_C241_n284, B => mult_21_C241_n281, Z => 
                           mult_21_C241_n279);
   mult_21_C241_U271 : AOI21D1 port map( A1 => mult_21_C241_n278, A2 => 
                           mult_21_C241_n286, B => mult_21_C241_n279, Z => 
                           mult_21_C241_n277);
   mult_21_C241_U269 : EXNOR2D1 port map( A1 => mult_21_C241_n282, A2 => 
                           mult_21_C241_n171, Z => N3240);
   mult_21_C241_U262 : AOI21D1 port map( A1 => mult_21_C241_n276, A2 => 
                           mult_21_C241_n1527, B => mult_21_C241_n273, Z => 
                           mult_21_C241_n271);
   mult_21_C241_U261 : EXNOR2D1 port map( A1 => mult_21_C241_n276, A2 => 
                           mult_21_C241_n170, Z => N3241);
   mult_21_C241_U254 : AOI21D1 port map( A1 => mult_21_C241_n1524, A2 => 
                           mult_21_C241_n273, B => mult_21_C241_n268, Z => 
                           mult_21_C241_n266);
   mult_21_C241_U252 : OAI21D1 port map( A1 => mult_21_C241_n265, A2 => 
                           mult_21_C241_n277, B => mult_21_C241_n266, Z => 
                           mult_21_C241_n264);
   mult_21_C241_U250 : EXOR2D1 port map( A1 => mult_21_C241_n271, A2 => 
                           mult_21_C241_n169, Z => N3242);
   mult_21_C241_U245 : OAI21D1 port map( A1 => mult_21_C241_n263, A2 => 
                           mult_21_C241_n261, B => mult_21_C241_n262, Z => 
                           mult_21_C241_n260);
   mult_21_C241_U244 : EXOR2D1 port map( A1 => mult_21_C241_n263, A2 => 
                           mult_21_C241_n168, Z => N3243);
   mult_21_C241_U239 : OAI21D1 port map( A1 => mult_21_C241_n258, A2 => 
                           mult_21_C241_n262, B => mult_21_C241_n259, Z => 
                           mult_21_C241_n257);
   mult_21_C241_U237 : AOI21D1 port map( A1 => mult_21_C241_n256, A2 => 
                           mult_21_C241_n264, B => mult_21_C241_n257, Z => 
                           mult_21_C241_n255);
   mult_21_C241_U235 : EXNOR2D1 port map( A1 => mult_21_C241_n260, A2 => 
                           mult_21_C241_n167, Z => N3244);
   mult_21_C241_U228 : AOI21D1 port map( A1 => mult_21_C241_n254, A2 => 
                           mult_21_C241_n1529, B => mult_21_C241_n251, Z => 
                           mult_21_C241_n249);
   mult_21_C241_U227 : EXNOR2D1 port map( A1 => mult_21_C241_n254, A2 => 
                           mult_21_C241_n166, Z => N3245);
   mult_21_C241_U220 : AOI21D1 port map( A1 => mult_21_C241_n1530, A2 => 
                           mult_21_C241_n251, B => mult_21_C241_n246, Z => 
                           mult_21_C241_n244);
   mult_21_C241_U218 : OAI21D1 port map( A1 => mult_21_C241_n255, A2 => 
                           mult_21_C241_n243, B => mult_21_C241_n244, Z => 
                           mult_21_C241_n242);
   mult_21_C241_U216 : EXOR2D1 port map( A1 => mult_21_C241_n249, A2 => 
                           mult_21_C241_n165, Z => N3246);
   mult_21_C241_U211 : OAI21D1 port map( A1 => mult_21_C241_n241, A2 => 
                           mult_21_C241_n239, B => mult_21_C241_n240, Z => 
                           mult_21_C241_n238);
   mult_21_C241_U210 : EXOR2D1 port map( A1 => mult_21_C241_n241, A2 => 
                           mult_21_C241_n164, Z => N3247);
   mult_21_C241_U205 : OAI21D1 port map( A1 => mult_21_C241_n236, A2 => 
                           mult_21_C241_n240, B => mult_21_C241_n237, Z => 
                           mult_21_C241_n235);
   mult_21_C241_U203 : AOI21D1 port map( A1 => mult_21_C241_n242, A2 => 
                           mult_21_C241_n234, B => mult_21_C241_n235, Z => 
                           mult_21_C241_n233);
   mult_21_C241_U201 : EXNOR2D1 port map( A1 => mult_21_C241_n238, A2 => 
                           mult_21_C241_n163, Z => N3248);
   mult_21_C241_U194 : AOI21D1 port map( A1 => mult_21_C241_n232, A2 => 
                           mult_21_C241_n313, B => mult_21_C241_n229, Z => 
                           mult_21_C241_n227);
   mult_21_C241_U193 : EXNOR2D1 port map( A1 => mult_21_C241_n232, A2 => 
                           mult_21_C241_n162, Z => N3249);
   mult_21_C241_U188 : OAI21D1 port map( A1 => mult_21_C241_n225, A2 => 
                           mult_21_C241_n231, B => mult_21_C241_n226, Z => 
                           mult_21_C241_n224);
   mult_21_C241_U186 : AOI21D1 port map( A1 => mult_21_C241_n232, A2 => 
                           mult_21_C241_n223, B => mult_21_C241_n224, Z => 
                           mult_21_C241_n222);
   mult_21_C241_U185 : EXOR2D1 port map( A1 => mult_21_C241_n227, A2 => 
                           mult_21_C241_n161, Z => N3250);
   mult_21_C241_U178 : AOI21D1 port map( A1 => mult_21_C241_n224, A2 => 
                           mult_21_C241_n1528, B => mult_21_C241_n219, Z => 
                           mult_21_C241_n217);
   mult_21_C241_U176 : OAI21D1 port map( A1 => mult_21_C241_n233, A2 => 
                           mult_21_C241_n216, B => mult_21_C241_n217, Z => 
                           mult_21_C241_n215);
   mult_21_C241_U174 : EXOR2D1 port map( A1 => mult_21_C241_n222, A2 => 
                           mult_21_C241_n160, Z => N3251);
   mult_21_C241_U165 : OAI21D1 port map( A1 => mult_21_C241_n214, A2 => 
                           mult_21_C241_n208, B => mult_21_C241_n209, Z => 
                           mult_21_C241_n207);
   mult_21_C241_U164 : EXOR2D1 port map( A1 => mult_21_C241_n214, A2 => 
                           mult_21_C241_n159, Z => N3252);
   mult_21_C241_U157 : AOI21D1 port map( A1 => mult_21_C241_n1525, A2 => 
                           mult_21_C241_n211, B => mult_21_C241_n204, Z => 
                           mult_21_C241_n202);
   mult_21_C241_U155 : OAI21D1 port map( A1 => mult_21_C241_n214, A2 => 
                           mult_21_C241_n201, B => mult_21_C241_n202, Z => 
                           mult_21_C241_n200);
   mult_21_C241_U154 : EXNOR2D1 port map( A1 => mult_21_C241_n207, A2 => 
                           mult_21_C241_n158, Z => N3253);
   mult_21_C241_U147 : AOI21D1 port map( A1 => mult_21_C241_n200, A2 => 
                           mult_21_C241_n1526, B => mult_21_C241_n197, Z => 
                           mult_21_C241_n195);
   mult_21_C241_U146 : EXNOR2D1 port map( A1 => mult_21_C241_n200, A2 => 
                           mult_21_C241_n157, Z => N3254);
   mult_21_C241_U137 : OAI21D1 port map( A1 => mult_21_C241_n202, A2 => 
                           mult_21_C241_n189, B => mult_21_C241_n190, Z => 
                           mult_21_C241_n188);
   mult_21_C241_U134 : EXOR2D1 port map( A1 => mult_21_C241_n195, A2 => 
                           mult_21_C241_n156, Z => N3255);
   mult_21_C241_U132 : ADFULD1 port map( A => mult_21_C241_n531, B => 
                           mult_21_C241_n552, CI => mult_21_C241_n1521, CO => 
                           mult_21_C241_n185, S => N3256);
   mult_21_C241_U131 : ADFULD1 port map( A => mult_21_C241_n507, B => 
                           mult_21_C241_n530, CI => mult_21_C241_n185, CO => 
                           mult_21_C241_n184, S => N3257);
   mult_21_C241_U130 : ADFULD1 port map( A => mult_21_C241_n483, B => 
                           mult_21_C241_n506, CI => mult_21_C241_n184, CO => 
                           mult_21_C241_n183, S => N3258);
   mult_21_C241_U129 : ADFULD1 port map( A => mult_21_C241_n457, B => 
                           mult_21_C241_n482, CI => mult_21_C241_n183, CO => 
                           mult_21_C241_n182, S => N3259);
   mult_21_C241_U128 : ADFULD1 port map( A => mult_21_C241_n431, B => 
                           mult_21_C241_n456, CI => mult_21_C241_n182, CO => 
                           mult_21_C241_n181, S => N3260);
   mult_21_C241_U127 : ADFULD1 port map( A => mult_21_C241_n403, B => 
                           mult_21_C241_n430, CI => mult_21_C241_n181, CO => 
                           mult_21_C241_n180, S => N3261);
   mult_21_C241_U126 : ADFULD1 port map( A => mult_21_C241_n375, B => 
                           mult_21_C241_n402, CI => mult_21_C241_n180, CO => 
                           mult_21_C241_n179, S => N3262);
   mult_21_C241_U125 : ADFULD1 port map( A => mult_21_C241_n345, B => 
                           mult_21_C241_n374, CI => mult_21_C241_n179, CO => 
                           mult_21_C241_n178, S => N3263);
   mult_21_C243_U1392 : INVD1 port map( A => N2976, Z => mult_21_C243_n1066);
   mult_21_C243_U1391 : INVD1 port map( A => N3108, Z => mult_21_C243_n1544);
   mult_21_C243_U1390 : INVD1 port map( A => N3106, Z => mult_21_C243_n1546);
   mult_21_C243_U1389 : AO21D1 port map( A1 => N2974, A2 => N2975, B => 
                           mult_21_C243_n1066, Z => mult_21_C243_n105);
   mult_21_C243_U1388 : INVD1 port map( A => N2974, Z => mult_21_C243_n1067);
   mult_21_C243_U1387 : AO21D1 port map( A1 => N2972, A2 => N2973, B => 
                           mult_21_C243_n1067, Z => mult_21_C243_n101);
   mult_21_C243_U1386 : EXOR2D1 port map( A1 => mult_21_C243_n1307, A2 => 
                           mult_21_C243_n1337, Z => mult_21_C243_n343);
   mult_21_C243_U1385 : INVD1 port map( A => N2972, Z => mult_21_C243_n1068);
   mult_21_C243_U1384 : AO21D1 port map( A1 => N2970, A2 => N2971, B => 
                           mult_21_C243_n1068, Z => mult_21_C243_n96);
   mult_21_C243_U1383 : ADHALFDL port map( A => mult_21_C243_n1309, B => 
                           mult_21_C243_n1339, CO => mult_21_C243_n400, S => 
                           mult_21_C243_n401);
   mult_21_C243_U1382 : AO21D1 port map( A1 => N2968, A2 => N2969, B => 
                           mult_21_C243_n1069, Z => mult_21_C243_n91);
   mult_21_C243_U1381 : INVD1 port map( A => N2970, Z => mult_21_C243_n1069);
   mult_21_C243_U1380 : ADHALFDL port map( A => mult_21_C243_n1311, B => 
                           mult_21_C243_n1341, CO => mult_21_C243_n454, S => 
                           mult_21_C243_n455);
   mult_21_C243_U1379 : OAI21D1 port map( A1 => N2968, A2 => N2969, B => 
                           mult_21_C243_n1069, Z => mult_21_C243_n89);
   mult_21_C243_U1378 : ADHALFDL port map( A => mult_21_C243_n1313, B => 
                           mult_21_C243_n1343, CO => mult_21_C243_n504, S => 
                           mult_21_C243_n505);
   mult_21_C243_U1377 : AO21D1 port map( A1 => N2966, A2 => N2967, B => 
                           mult_21_C243_n1070, Z => mult_21_C243_n86);
   mult_21_C243_U1376 : INVD1 port map( A => N2968, Z => mult_21_C243_n1070);
   mult_21_C243_U1375 : OAI21D1 port map( A1 => N2966, A2 => N2967, B => 
                           mult_21_C243_n1070, Z => mult_21_C243_n84);
   mult_21_C243_U1374 : AO21D1 port map( A1 => N2964, A2 => N2965, B => 
                           mult_21_C243_n1071, Z => mult_21_C243_n81);
   mult_21_C243_U1373 : INVD1 port map( A => N2966, Z => mult_21_C243_n1071);
   mult_21_C243_U1372 : OAI21D1 port map( A1 => N2964, A2 => N2965, B => 
                           mult_21_C243_n1071, Z => mult_21_C243_n79);
   mult_21_C243_U1371 : EXNOR2D1 port map( A1 => N2966, A2 => N2967, Z => 
                           mult_21_C243_n88);
   mult_21_C243_U1370 : AO21D1 port map( A1 => N2962, A2 => N2963, B => 
                           mult_21_C243_n1072, Z => mult_21_C243_n76);
   mult_21_C243_U1369 : OAI21D1 port map( A1 => N2954, A2 => N2955, B => 
                           mult_21_C243_n1076, Z => mult_21_C243_n42);
   mult_21_C243_U1368 : INVD1 port map( A => N2964, Z => mult_21_C243_n1072);
   mult_21_C243_U1367 : OAI21D1 port map( A1 => N2962, A2 => N2963, B => 
                           mult_21_C243_n1072, Z => mult_21_C243_n73);
   mult_21_C243_U1366 : INVD1 port map( A => N2956, Z => mult_21_C243_n1076);
   mult_21_C243_U1365 : AO21D1 port map( A1 => N2954, A2 => N2955, B => 
                           mult_21_C243_n1076, Z => mult_21_C243_n45);
   mult_21_C243_U1364 : OAI21D1 port map( A1 => N2960, A2 => N2961, B => 
                           mult_21_C243_n1073, Z => mult_21_C243_n66);
   mult_21_C243_U1363 : INVD1 port map( A => N2962, Z => mult_21_C243_n1073);
   mult_21_C243_U1362 : OAI21D1 port map( A1 => N2958, A2 => N2959, B => 
                           mult_21_C243_n1074, Z => mult_21_C243_n58);
   mult_21_C243_U1361 : INVD1 port map( A => N2960, Z => mult_21_C243_n1074);
   mult_21_C243_U1360 : AO21D1 port map( A1 => N2960, A2 => N2961, B => 
                           mult_21_C243_n1073, Z => mult_21_C243_n69);
   mult_21_C243_U1359 : AO21D1 port map( A1 => N2958, A2 => N2959, B => 
                           mult_21_C243_n1074, Z => mult_21_C243_n61);
   mult_21_C243_U1358 : OAI21D1 port map( A1 => N2956, A2 => N2957, B => 
                           mult_21_C243_n1075, Z => mult_21_C243_n50);
   mult_21_C243_U1357 : AO21D1 port map( A1 => N2952, A2 => N2953, B => 
                           mult_21_C243_n1077, Z => mult_21_C243_n38);
   mult_21_C243_U1356 : AO21D1 port map( A1 => N2948, A2 => N2949, B => 
                           mult_21_C243_n1079, Z => mult_21_C243_n22);
   mult_21_C243_U1355 : ADHALFDL port map( A => mult_21_C243_n1315, B => 
                           mult_21_C243_n1345, CO => mult_21_C243_n550, S => 
                           mult_21_C243_n551);
   mult_21_C243_U1354 : INVD1 port map( A => N2958, Z => mult_21_C243_n1075);
   mult_21_C243_U1353 : AO21D1 port map( A1 => N2956, A2 => N2957, B => 
                           mult_21_C243_n1075, Z => mult_21_C243_n53);
   mult_21_C243_U1352 : EXNOR2D1 port map( A1 => N2964, A2 => N2965, Z => 
                           mult_21_C243_n83);
   mult_21_C243_U1351 : INVD1 port map( A => N2945, Z => mult_21_C243_n8);
   mult_21_C243_U1350 : AO21D1 port map( A1 => N2950, A2 => N2951, B => 
                           mult_21_C243_n1078, Z => mult_21_C243_n30);
   mult_21_C243_U1349 : INVD1 port map( A => mult_21_C243_n1544, Z => 
                           mult_21_C243_n1543);
   mult_21_C243_U1348 : AO21D1 port map( A1 => N2946, A2 => N2947, B => 
                           mult_21_C243_n1080, Z => mult_21_C243_n14);
   mult_21_C243_U1347 : EXNOR2D1 port map( A1 => N2962, A2 => N2963, Z => 
                           mult_21_C243_n78);
   mult_21_C243_U1346 : INVD1 port map( A => mult_21_C243_n1546, Z => 
                           mult_21_C243_n1545);
   mult_21_C243_U1345 : EXNOR2D1 port map( A1 => N2954, A2 => N2955, Z => 
                           mult_21_C243_n48);
   mult_21_C243_U1344 : INVD1 port map( A => N2950, Z => mult_21_C243_n1079);
   mult_21_C243_U1343 : EXNOR2D1 port map( A1 => N2960, A2 => N2961, Z => 
                           mult_21_C243_n71);
   mult_21_C243_U1342 : EXNOR2D1 port map( A1 => N2958, A2 => N2959, Z => 
                           mult_21_C243_n63);
   mult_21_C243_U1341 : INVD1 port map( A => N2954, Z => mult_21_C243_n1077);
   mult_21_C243_U1340 : INVD1 port map( A => N2946, Z => mult_21_C243_n6);
   mult_21_C243_U1339 : NAN2D1 port map( A1 => N2945, A2 => mult_21_C243_n6, Z 
                           => mult_21_C243_n3);
   mult_21_C243_U1338 : INVD1 port map( A => N2952, Z => mult_21_C243_n1078);
   mult_21_C243_U1337 : EXNOR2D1 port map( A1 => N2956, A2 => N2957, Z => 
                           mult_21_C243_n56);
   mult_21_C243_U1336 : INVD1 port map( A => N2948, Z => mult_21_C243_n1080);
   mult_21_C243_U1335 : OA21D1 port map( A1 => N2950, A2 => N2951, B => 
                           mult_21_C243_n1078, Z => mult_21_C243_n1537);
   mult_21_C243_U1334 : ADHALFDL port map( A => mult_21_C243_n1325, B => 
                           mult_21_C243_n1355, CO => mult_21_C243_n720, S => 
                           mult_21_C243_n721);
   mult_21_C243_U1333 : ADHALFDL port map( A => mult_21_C243_n1321, B => 
                           mult_21_C243_n1351, CO => mult_21_C243_n664, S => 
                           mult_21_C243_n665);
   mult_21_C243_U1332 : ADHALFDL port map( A => mult_21_C243_n1319, B => 
                           mult_21_C243_n1349, CO => mult_21_C243_n630, S => 
                           mult_21_C243_n631);
   mult_21_C243_U1331 : ADHALFDL port map( A => mult_21_C243_n1327, B => 
                           mult_21_C243_n1357, CO => mult_21_C243_n742, S => 
                           mult_21_C243_n743);
   mult_21_C243_U1330 : ADHALFDL port map( A => mult_21_C243_n1317, B => 
                           mult_21_C243_n1347, CO => mult_21_C243_n592, S => 
                           mult_21_C243_n593);
   mult_21_C243_U1329 : EXOR2D1 port map( A1 => N2952, A2 => N2953, Z => 
                           mult_21_C243_n1536);
   mult_21_C243_U1328 : EXOR2D1 port map( A1 => N2948, A2 => N2949, Z => 
                           mult_21_C243_n1535);
   mult_21_C243_U1327 : EXOR2D1 port map( A1 => N2950, A2 => N2951, Z => 
                           mult_21_C243_n1534);
   mult_21_C243_U1326 : ADHALFDL port map( A => mult_21_C243_n1323, B => 
                           mult_21_C243_n1353, CO => mult_21_C243_n694, S => 
                           mult_21_C243_n695);
   mult_21_C243_U1325 : EXOR2D1 port map( A1 => N2946, A2 => N2947, Z => 
                           mult_21_C243_n1533);
   mult_21_C243_U1324 : ADHALFDL port map( A => mult_21_C243_n1329, B => 
                           mult_21_C243_n1359, CO => mult_21_C243_n760, S => 
                           mult_21_C243_n761);
   mult_21_C243_U1323 : ADHALFDL port map( A => mult_21_C243_n1098, B => 
                           mult_21_C243_n1081, CO => mult_21_C243_n372, S => 
                           mult_21_C243_n373);
   mult_21_C243_U1322 : ADHALFDL port map( A => mult_21_C243_n1102, B => 
                           mult_21_C243_n1082, CO => mult_21_C243_n428, S => 
                           mult_21_C243_n429);
   mult_21_C243_U1321 : ADHALFDL port map( A => mult_21_C243_n1108, B => 
                           mult_21_C243_n1083, CO => mult_21_C243_n480, S => 
                           mult_21_C243_n481);
   mult_21_C243_U1320 : ADHALFDL port map( A => mult_21_C243_n1116, B => 
                           mult_21_C243_n1084, CO => mult_21_C243_n528, S => 
                           mult_21_C243_n529);
   mult_21_C243_U1319 : ADHALFDL port map( A => mult_21_C243_n1126, B => 
                           mult_21_C243_n1085, CO => mult_21_C243_n572, S => 
                           mult_21_C243_n573);
   mult_21_C243_U1318 : INVD1 port map( A => mult_21_C243_n1367, Z => 
                           mult_21_C243_n303);
   mult_21_C243_U1317 : ADHALFDL port map( A => mult_21_C243_n1138, B => 
                           mult_21_C243_n1086, CO => mult_21_C243_n612, S => 
                           mult_21_C243_n613);
   mult_21_C243_U1316 : ADHALFDL port map( A => mult_21_C243_n1186, B => 
                           mult_21_C243_n1089, CO => mult_21_C243_n708, S => 
                           mult_21_C243_n709);
   mult_21_C243_U1315 : ADHALFDL port map( A => mult_21_C243_n1228, B => 
                           mult_21_C243_n1091, CO => mult_21_C243_n752, S => 
                           mult_21_C243_n753);
   mult_21_C243_U1314 : ADHALFDL port map( A => mult_21_C243_n1152, B => 
                           mult_21_C243_n1087, CO => mult_21_C243_n648, S => 
                           mult_21_C243_n649);
   mult_21_C243_U1313 : ADHALFDL port map( A => mult_21_C243_n1168, B => 
                           mult_21_C243_n1088, CO => mult_21_C243_n680, S => 
                           mult_21_C243_n681);
   mult_21_C243_U1312 : ADHALFDL port map( A => mult_21_C243_n1206, B => 
                           mult_21_C243_n1090, CO => mult_21_C243_n732, S => 
                           mult_21_C243_n733);
   mult_21_C243_U1311 : INVD1 port map( A => mult_21_C243_n1537, Z => 
                           mult_21_C243_n1540);
   mult_21_C243_U1310 : ADHALFDL port map( A => mult_21_C243_n1306, B => 
                           mult_21_C243_n1094, CO => mult_21_C243_n788, S => 
                           mult_21_C243_n789);
   mult_21_C243_U1309 : ADHALFDL port map( A => mult_21_C243_n1333, B => 
                           mult_21_C243_n1363, CO => mult_21_C243_n784, S => 
                           mult_21_C243_n785);
   mult_21_C243_U1308 : ADHALFDL port map( A => mult_21_C243_n1252, B => 
                           mult_21_C243_n1092, CO => mult_21_C243_n768, S => 
                           mult_21_C243_n769);
   mult_21_C243_U1307 : ADHALFDL port map( A => mult_21_C243_n1331, B => 
                           mult_21_C243_n1361, CO => mult_21_C243_n774, S => 
                           mult_21_C243_n775);
   mult_21_C243_U1306 : INVD1 port map( A => mult_21_C243_n1536, Z => 
                           mult_21_C243_n1538);
   mult_21_C243_U1305 : INVD1 port map( A => mult_21_C243_n1535, Z => 
                           mult_21_C243_n1541);
   mult_21_C243_U1304 : NOR2D1 port map( A1 => mult_21_C243_n1537, A2 => 
                           mult_21_C243_n30, Z => mult_21_C243_n1093);
   mult_21_C243_U1303 : INVD1 port map( A => mult_21_C243_n1534, Z => 
                           mult_21_C243_n1539);
   mult_21_C243_U1302 : ADHALFDL port map( A => mult_21_C243_n1336, B => 
                           mult_21_C243_n1095, CO => mult_21_C243_n792, S => 
                           mult_21_C243_n793);
   mult_21_C243_U1301 : ADHALFDL port map( A => mult_21_C243_n1335, B => 
                           mult_21_C243_n1365, CO => mult_21_C243_n790, S => 
                           mult_21_C243_n791);
   mult_21_C243_U1300 : EXOR2D1 port map( A1 => mult_21_C243_n329, A2 => 
                           mult_21_C243_n344, Z => mult_21_C243_n155);
   mult_21_C243_U1299 : EXOR2D1 port map( A1 => mult_21_C243_n178, A2 => 
                           mult_21_C243_n155, Z => N3296);
   mult_21_C243_U1298 : INVD1 port map( A => mult_21_C243_n1533, Z => 
                           mult_21_C243_n1542);
   mult_21_C243_U1297 : NOR2D1 port map( A1 => mult_21_C243_n303, A2 => 
                           mult_21_C243_n305, Z => mult_21_C243_n302);
   mult_21_C243_U1296 : NAN2D1 port map( A1 => mult_21_C243_n1368, A2 => 
                           mult_21_C243_n1096, Z => mult_21_C243_n305);
   mult_21_C243_U1295 : NAN2D1 port map( A1 => mult_21_C243_n791, A2 => 
                           mult_21_C243_n792, Z => mult_21_C243_n296);
   mult_21_C243_U1294 : NAN2D1 port map( A1 => mult_21_C243_n783, A2 => 
                           mult_21_C243_n786, Z => mult_21_C243_n288);
   mult_21_C243_U1293 : NOR2D1 port map( A1 => mult_21_C243_n791, A2 => 
                           mult_21_C243_n792, Z => mult_21_C243_n295);
   mult_21_C243_U1292 : NOR2D1 port map( A1 => mult_21_C243_n783, A2 => 
                           mult_21_C243_n786, Z => mult_21_C243_n287);
   mult_21_C243_U1291 : NAN2D1 port map( A1 => mult_21_C243_n777, A2 => 
                           mult_21_C243_n782, Z => mult_21_C243_n284);
   mult_21_C243_U1290 : NAN2D1 port map( A1 => mult_21_C243_n793, A2 => 
                           mult_21_C243_n1366, Z => mult_21_C243_n301);
   mult_21_C243_U1289 : NAN2D1 port map( A1 => mult_21_C243_n787, A2 => 
                           mult_21_C243_n789, Z => mult_21_C243_n293);
   mult_21_C243_U1288 : NOR2D1 port map( A1 => mult_21_C243_n777, A2 => 
                           mult_21_C243_n782, Z => mult_21_C243_n283);
   mult_21_C243_U1287 : OR2D1 port map( A1 => mult_21_C243_n793, A2 => 
                           mult_21_C243_n1366, Z => mult_21_C243_n1532);
   mult_21_C243_U1286 : OR2D1 port map( A1 => mult_21_C243_n787, A2 => 
                           mult_21_C243_n789, Z => mult_21_C243_n1531);
   mult_21_C243_U1285 : NAN2D1 port map( A1 => mult_21_C243_n1532, A2 => 
                           mult_21_C243_n301, Z => mult_21_C243_n176);
   mult_21_C243_U1284 : INVD1 port map( A => mult_21_C243_n295, Z => 
                           mult_21_C243_n326);
   mult_21_C243_U1283 : NAN2D1 port map( A1 => mult_21_C243_n326, A2 => 
                           mult_21_C243_n296, Z => mult_21_C243_n175);
   mult_21_C243_U1282 : NAN2D1 port map( A1 => mult_21_C243_n1531, A2 => 
                           mult_21_C243_n293, Z => mult_21_C243_n174);
   mult_21_C243_U1281 : INVD1 port map( A => mult_21_C243_n287, Z => 
                           mult_21_C243_n324);
   mult_21_C243_U1280 : NAN2D1 port map( A1 => mult_21_C243_n324, A2 => 
                           mult_21_C243_n288, Z => mult_21_C243_n173);
   mult_21_C243_U1279 : INVD1 port map( A => mult_21_C243_n283, Z => 
                           mult_21_C243_n323);
   mult_21_C243_U1278 : NAN2D1 port map( A1 => mult_21_C243_n323, A2 => 
                           mult_21_C243_n284, Z => mult_21_C243_n172);
   mult_21_C243_U1277 : INVD1 port map( A => mult_21_C243_n280, Z => 
                           mult_21_C243_n322);
   mult_21_C243_U1276 : NAN2D1 port map( A1 => mult_21_C243_n322, A2 => 
                           mult_21_C243_n281, Z => mult_21_C243_n171);
   mult_21_C243_U1275 : NAN2D1 port map( A1 => mult_21_C243_n697, A2 => 
                           mult_21_C243_n710, Z => mult_21_C243_n240);
   mult_21_C243_U1274 : NAN2D1 port map( A1 => mult_21_C243_n633, A2 => 
                           mult_21_C243_n650, Z => mult_21_C243_n221);
   mult_21_C243_U1273 : NAN2D1 port map( A1 => mult_21_C243_n711, A2 => 
                           mult_21_C243_n722, Z => mult_21_C243_n248);
   mult_21_C243_U1272 : NOR2D1 port map( A1 => mult_21_C243_n697, A2 => 
                           mult_21_C243_n710, Z => mult_21_C243_n239);
   mult_21_C243_U1271 : NOR2D1 port map( A1 => mult_21_C243_n615, A2 => 
                           mult_21_C243_n632, Z => mult_21_C243_n208);
   mult_21_C243_U1270 : NAN2D1 port map( A1 => mult_21_C243_n735, A2 => 
                           mult_21_C243_n744, Z => mult_21_C243_n259);
   mult_21_C243_U1269 : NAN2D1 port map( A1 => mult_21_C243_n771, A2 => 
                           mult_21_C243_n776, Z => mult_21_C243_n281);
   mult_21_C243_U1268 : NAN2D1 port map( A1 => mult_21_C243_n615, A2 => 
                           mult_21_C243_n632, Z => mult_21_C243_n209);
   mult_21_C243_U1267 : OR2D1 port map( A1 => mult_21_C243_n711, A2 => 
                           mult_21_C243_n722, Z => mult_21_C243_n1530);
   mult_21_C243_U1266 : NAN2D1 port map( A1 => mult_21_C243_n745, A2 => 
                           mult_21_C243_n754, Z => mult_21_C243_n262);
   mult_21_C243_U1265 : OR2D1 port map( A1 => mult_21_C243_n723, A2 => 
                           mult_21_C243_n734, Z => mult_21_C243_n1529);
   mult_21_C243_U1264 : OR2D1 port map( A1 => mult_21_C243_n633, A2 => 
                           mult_21_C243_n650, Z => mult_21_C243_n1528);
   mult_21_C243_U1263 : NAN2D1 port map( A1 => mult_21_C243_n595, A2 => 
                           mult_21_C243_n614, Z => mult_21_C243_n206);
   mult_21_C243_U1262 : OR2D1 port map( A1 => mult_21_C243_n763, A2 => 
                           mult_21_C243_n770, Z => mult_21_C243_n1527);
   mult_21_C243_U1261 : NAN2D1 port map( A1 => mult_21_C243_n651, A2 => 
                           mult_21_C243_n666, Z => mult_21_C243_n226);
   mult_21_C243_U1260 : NAN2D1 port map( A1 => mult_21_C243_n723, A2 => 
                           mult_21_C243_n734, Z => mult_21_C243_n253);
   mult_21_C243_U1259 : NAN2D1 port map( A1 => mult_21_C243_n575, A2 => 
                           mult_21_C243_n594, Z => mult_21_C243_n199);
   mult_21_C243_U1258 : OR2D1 port map( A1 => mult_21_C243_n575, A2 => 
                           mult_21_C243_n594, Z => mult_21_C243_n1526);
   mult_21_C243_U1257 : NAN2D1 port map( A1 => mult_21_C243_n763, A2 => 
                           mult_21_C243_n770, Z => mult_21_C243_n275);
   mult_21_C243_U1256 : NOR2D1 port map( A1 => mult_21_C243_n735, A2 => 
                           mult_21_C243_n744, Z => mult_21_C243_n258);
   mult_21_C243_U1255 : NOR2D1 port map( A1 => mult_21_C243_n745, A2 => 
                           mult_21_C243_n754, Z => mult_21_C243_n261);
   mult_21_C243_U1254 : NOR2D1 port map( A1 => mult_21_C243_n771, A2 => 
                           mult_21_C243_n776, Z => mult_21_C243_n280);
   mult_21_C243_U1253 : OR2D1 port map( A1 => mult_21_C243_n595, A2 => 
                           mult_21_C243_n614, Z => mult_21_C243_n1525);
   mult_21_C243_U1252 : OA21M20D1 port map( A1 => mult_21_C243_n1532, A2 => 
                           mult_21_C243_n302, B => mult_21_C243_n301, Z => 
                           mult_21_C243_n297);
   mult_21_C243_U1251 : NOR2D1 port map( A1 => mult_21_C243_n651, A2 => 
                           mult_21_C243_n666, Z => mult_21_C243_n225);
   mult_21_C243_U1250 : OA21M20D1 port map( A1 => mult_21_C243_n1531, A2 => 
                           mult_21_C243_n294, B => mult_21_C243_n293, Z => 
                           mult_21_C243_n289);
   mult_21_C243_U1249 : NOR2D1 port map( A1 => mult_21_C243_n280, A2 => 
                           mult_21_C243_n283, Z => mult_21_C243_n278);
   mult_21_C243_U1248 : NAN2D1 port map( A1 => mult_21_C243_n755, A2 => 
                           mult_21_C243_n762, Z => mult_21_C243_n270);
   mult_21_C243_U1247 : OR2D1 port map( A1 => mult_21_C243_n755, A2 => 
                           mult_21_C243_n762, Z => mult_21_C243_n1524);
   mult_21_C243_U1246 : INVD1 port map( A => mult_21_C243_n286, Z => 
                           mult_21_C243_n285);
   mult_21_C243_U1245 : NAN2D1 port map( A1 => mult_21_C243_n1527, A2 => 
                           mult_21_C243_n275, Z => mult_21_C243_n170);
   mult_21_C243_U1244 : NAN2D1 port map( A1 => mult_21_C243_n1524, A2 => 
                           mult_21_C243_n270, Z => mult_21_C243_n169);
   mult_21_C243_U1243 : INVD1 port map( A => mult_21_C243_n277, Z => 
                           mult_21_C243_n276);
   mult_21_C243_U1242 : INVD1 port map( A => mult_21_C243_n261, Z => 
                           mult_21_C243_n319);
   mult_21_C243_U1241 : NAN2D1 port map( A1 => mult_21_C243_n319, A2 => 
                           mult_21_C243_n262, Z => mult_21_C243_n168);
   mult_21_C243_U1240 : INVD1 port map( A => mult_21_C243_n258, Z => 
                           mult_21_C243_n318);
   mult_21_C243_U1239 : NAN2D1 port map( A1 => mult_21_C243_n318, A2 => 
                           mult_21_C243_n259, Z => mult_21_C243_n167);
   mult_21_C243_U1238 : NAN2D1 port map( A1 => mult_21_C243_n1529, A2 => 
                           mult_21_C243_n253, Z => mult_21_C243_n166);
   mult_21_C243_U1237 : INVD1 port map( A => mult_21_C243_n239, Z => 
                           mult_21_C243_n315);
   mult_21_C243_U1236 : NAN2D1 port map( A1 => mult_21_C243_n315, A2 => 
                           mult_21_C243_n240, Z => mult_21_C243_n164);
   mult_21_C243_U1235 : NAN2D1 port map( A1 => mult_21_C243_n1530, A2 => 
                           mult_21_C243_n248, Z => mult_21_C243_n165);
   mult_21_C243_U1234 : INVD1 port map( A => mult_21_C243_n236, Z => 
                           mult_21_C243_n314);
   mult_21_C243_U1233 : NAN2D1 port map( A1 => mult_21_C243_n314, A2 => 
                           mult_21_C243_n237, Z => mult_21_C243_n163);
   mult_21_C243_U1232 : NAN2D1 port map( A1 => mult_21_C243_n1528, A2 => 
                           mult_21_C243_n221, Z => mult_21_C243_n160);
   mult_21_C243_U1231 : INVD1 port map( A => mult_21_C243_n225, Z => 
                           mult_21_C243_n312);
   mult_21_C243_U1230 : NAN2D1 port map( A1 => mult_21_C243_n312, A2 => 
                           mult_21_C243_n226, Z => mult_21_C243_n161);
   mult_21_C243_U1229 : NAN2D1 port map( A1 => mult_21_C243_n310, A2 => 
                           mult_21_C243_n209, Z => mult_21_C243_n159);
   mult_21_C243_U1228 : NAN2D1 port map( A1 => mult_21_C243_n1525, A2 => 
                           mult_21_C243_n206, Z => mult_21_C243_n158);
   mult_21_C243_U1227 : NAN2D1 port map( A1 => mult_21_C243_n1526, A2 => 
                           mult_21_C243_n199, Z => mult_21_C243_n157);
   mult_21_C243_U1226 : NAN2D1 port map( A1 => mult_21_C243_n1523, A2 => 
                           mult_21_C243_n194, Z => mult_21_C243_n156);
   mult_21_C243_U1225 : NAN2D1 port map( A1 => mult_21_C243_n683, A2 => 
                           mult_21_C243_n696, Z => mult_21_C243_n237);
   mult_21_C243_U1224 : NOR2D1 port map( A1 => mult_21_C243_n667, A2 => 
                           mult_21_C243_n682, Z => mult_21_C243_n230);
   mult_21_C243_U1223 : INVD1 port map( A => mult_21_C243_n208, Z => 
                           mult_21_C243_n310);
   mult_21_C243_U1222 : NAN2D1 port map( A1 => mult_21_C243_n553, A2 => 
                           mult_21_C243_n574, Z => mult_21_C243_n194);
   mult_21_C243_U1221 : NOR2D1 port map( A1 => mult_21_C243_n683, A2 => 
                           mult_21_C243_n696, Z => mult_21_C243_n236);
   mult_21_C243_U1220 : NAN2D1 port map( A1 => mult_21_C243_n1525, A2 => 
                           mult_21_C243_n310, Z => mult_21_C243_n201);
   mult_21_C243_U1219 : NOR2D1 port map( A1 => mult_21_C243_n225, A2 => 
                           mult_21_C243_n230, Z => mult_21_C243_n223);
   mult_21_C243_U1218 : NAN2D1 port map( A1 => mult_21_C243_n667, A2 => 
                           mult_21_C243_n682, Z => mult_21_C243_n231);
   mult_21_C243_U1217 : INVD1 port map( A => mult_21_C243_n253, Z => 
                           mult_21_C243_n251);
   mult_21_C243_U1216 : INVD1 port map( A => mult_21_C243_n199, Z => 
                           mult_21_C243_n197);
   mult_21_C243_U1215 : NAN2D1 port map( A1 => mult_21_C243_n1523, A2 => 
                           mult_21_C243_n1526, Z => mult_21_C243_n189);
   mult_21_C243_U1214 : OR2D1 port map( A1 => mult_21_C243_n553, A2 => 
                           mult_21_C243_n574, Z => mult_21_C243_n1523);
   mult_21_C243_U1213 : INVD1 port map( A => mult_21_C243_n275, Z => 
                           mult_21_C243_n273);
   mult_21_C243_U1212 : INVD1 port map( A => mult_21_C243_n206, Z => 
                           mult_21_C243_n204);
   mult_21_C243_U1211 : INVD1 port map( A => mult_21_C243_n209, Z => 
                           mult_21_C243_n211);
   mult_21_C243_U1210 : NOR2D1 port map( A1 => mult_21_C243_n189, A2 => 
                           mult_21_C243_n201, Z => mult_21_C243_n187);
   mult_21_C243_U1209 : NOR2D1 port map( A1 => mult_21_C243_n236, A2 => 
                           mult_21_C243_n239, Z => mult_21_C243_n234);
   mult_21_C243_U1208 : NOR2D1 port map( A1 => mult_21_C243_n258, A2 => 
                           mult_21_C243_n261, Z => mult_21_C243_n256);
   mult_21_C243_U1207 : INVD1 port map( A => mult_21_C243_n270, Z => 
                           mult_21_C243_n268);
   mult_21_C243_U1206 : NAN2D1 port map( A1 => mult_21_C243_n1524, A2 => 
                           mult_21_C243_n1527, Z => mult_21_C243_n265);
   mult_21_C243_U1205 : INVD1 port map( A => mult_21_C243_n248, Z => 
                           mult_21_C243_n246);
   mult_21_C243_U1204 : NAN2D1 port map( A1 => mult_21_C243_n1530, A2 => 
                           mult_21_C243_n1529, Z => mult_21_C243_n243);
   mult_21_C243_U1203 : INVD1 port map( A => mult_21_C243_n221, Z => 
                           mult_21_C243_n219);
   mult_21_C243_U1202 : NAN2D1 port map( A1 => mult_21_C243_n223, A2 => 
                           mult_21_C243_n1528, Z => mult_21_C243_n216);
   mult_21_C243_U1201 : INVD1 port map( A => mult_21_C243_n264, Z => 
                           mult_21_C243_n263);
   mult_21_C243_U1200 : INVD1 port map( A => mult_21_C243_n231, Z => 
                           mult_21_C243_n229);
   mult_21_C243_U1199 : INVD1 port map( A => mult_21_C243_n230, Z => 
                           mult_21_C243_n313);
   mult_21_C243_U1198 : INVD1 port map( A => mult_21_C243_n255, Z => 
                           mult_21_C243_n254);
   mult_21_C243_U1197 : INVD1 port map( A => mult_21_C243_n242, Z => 
                           mult_21_C243_n241);
   mult_21_C243_U1196 : NAN2D1 port map( A1 => mult_21_C243_n313, A2 => 
                           mult_21_C243_n231, Z => mult_21_C243_n162);
   mult_21_C243_U1195 : INVD1 port map( A => mult_21_C243_n233, Z => 
                           mult_21_C243_n232);
   mult_21_C243_U1194 : INVD1 port map( A => mult_21_C243_n215, Z => 
                           mult_21_C243_n214);
   mult_21_C243_U1193 : OA21M20D1 port map( A1 => mult_21_C243_n1523, A2 => 
                           mult_21_C243_n197, B => mult_21_C243_n194, Z => 
                           mult_21_C243_n190);
   mult_21_C243_U1192 : OR2D1 port map( A1 => mult_21_C243_n1368, A2 => 
                           mult_21_C243_n1096, Z => mult_21_C243_n1522);
   mult_21_C243_U1191 : AO21D1 port map( A1 => mult_21_C243_n215, A2 => 
                           mult_21_C243_n187, B => mult_21_C243_n188, Z => 
                           mult_21_C243_n1521);
   mult_21_C243_U1190 : AND2D1 port map( A1 => mult_21_C243_n1522, A2 => 
                           mult_21_C243_n305, Z => N3265);
   mult_21_C243_U1189 : OAI21D1 port map( A1 => N2952, A2 => N2953, B => 
                           mult_21_C243_n1077, Z => mult_21_C243_n1519);
   mult_21_C243_U1188 : OAI21D1 port map( A1 => N2948, A2 => N2949, B => 
                           mult_21_C243_n1079, Z => mult_21_C243_n1518);
   mult_21_C243_U1187 : OAI21D1 port map( A1 => N2946, A2 => N2947, B => 
                           mult_21_C243_n1080, Z => mult_21_C243_n1517);
   mult_21_C243_U1186 : ADHALFDL port map( A => mult_21_C243_n1278, B => 
                           mult_21_C243_n1093, CO => mult_21_C243_n780, S => 
                           mult_21_C243_n781);
   mult_21_C243_U1135 : EXNOR2D1 port map( A1 => N2968, A2 => N2969, Z => 
                           mult_21_C243_n93);
   mult_21_C243_U1131 : EXNOR2D1 port map( A1 => N2970, A2 => N2971, Z => 
                           mult_21_C243_n98);
   mult_21_C243_U1129 : OAI21D1 port map( A1 => N2970, A2 => N2971, B => 
                           mult_21_C243_n1068, Z => mult_21_C243_n94);
   mult_21_C243_U1127 : EXNOR2D1 port map( A1 => N2972, A2 => N2973, Z => 
                           mult_21_C243_n103);
   mult_21_C243_U1125 : OAI21D1 port map( A1 => N2972, A2 => N2973, B => 
                           mult_21_C243_n1067, Z => mult_21_C243_n99);
   mult_21_C243_U1123 : EXNOR2D1 port map( A1 => N2974, A2 => N2975, Z => 
                           mult_21_C243_n106);
   mult_21_C243_U1121 : OAI21D1 port map( A1 => N2974, A2 => N2975, B => 
                           mult_21_C243_n1066, Z => mult_21_C243_n104);
   mult_21_C243_U1120 : NAN2M1D1 port map( A1 => mult_21_C243_n8, A2 => N3105, 
                           Z => mult_21_C243_n1065);
   mult_21_C243_U1119 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1065, Z => 
                           mult_21_C243_n1368);
   mult_21_C243_U1118 : MUXB2DL port map( A0 => N3106, A1 => N3105, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1064);
   mult_21_C243_U1117 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1064, Z => 
                           mult_21_C243_n1367);
   mult_21_C243_U1116 : MUXB2DL port map( A0 => N3107, A1 => mult_21_C243_n1545
                           , SL => mult_21_C243_n8, Z => mult_21_C243_n1063);
   mult_21_C243_U1115 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1063, Z => 
                           mult_21_C243_n1366);
   mult_21_C243_U1114 : MUXB2DL port map( A0 => N3108, A1 => N3107, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1062);
   mult_21_C243_U1113 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1062, Z => 
                           mult_21_C243_n1365);
   mult_21_C243_U1112 : MUXB2DL port map( A0 => N3109, A1 => mult_21_C243_n1543
                           , SL => mult_21_C243_n8, Z => mult_21_C243_n1061);
   mult_21_C243_U1111 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1061, Z => 
                           mult_21_C243_n1364);
   mult_21_C243_U1110 : MUXB2DL port map( A0 => N3110, A1 => N3109, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1060);
   mult_21_C243_U1109 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1060, Z => 
                           mult_21_C243_n1363);
   mult_21_C243_U1108 : MUXB2DL port map( A0 => N3111, A1 => N3110, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1059);
   mult_21_C243_U1107 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1059, Z => 
                           mult_21_C243_n1362);
   mult_21_C243_U1106 : MUXB2DL port map( A0 => N3112, A1 => N3111, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1058);
   mult_21_C243_U1105 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1058, Z => 
                           mult_21_C243_n1361);
   mult_21_C243_U1104 : MUXB2DL port map( A0 => N3113, A1 => N3112, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1057);
   mult_21_C243_U1103 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1057, Z => 
                           mult_21_C243_n1360);
   mult_21_C243_U1102 : MUXB2DL port map( A0 => N3114, A1 => N3113, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1056);
   mult_21_C243_U1101 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1056, Z => 
                           mult_21_C243_n1359);
   mult_21_C243_U1100 : MUXB2DL port map( A0 => N3115, A1 => N3114, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1055);
   mult_21_C243_U1099 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1055, Z => 
                           mult_21_C243_n1358);
   mult_21_C243_U1098 : MUXB2DL port map( A0 => N3116, A1 => N3115, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1054);
   mult_21_C243_U1097 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1054, Z => 
                           mult_21_C243_n1357);
   mult_21_C243_U1096 : MUXB2DL port map( A0 => N3117, A1 => N3116, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1053);
   mult_21_C243_U1095 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1053, Z => 
                           mult_21_C243_n1356);
   mult_21_C243_U1094 : MUXB2DL port map( A0 => N3118, A1 => N3117, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1052);
   mult_21_C243_U1093 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1052, Z => 
                           mult_21_C243_n1355);
   mult_21_C243_U1092 : MUXB2DL port map( A0 => N3119, A1 => N3118, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1051);
   mult_21_C243_U1091 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1051, Z => 
                           mult_21_C243_n1354);
   mult_21_C243_U1090 : MUXB2DL port map( A0 => N3120, A1 => N3119, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1050);
   mult_21_C243_U1089 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1050, Z => 
                           mult_21_C243_n1353);
   mult_21_C243_U1088 : MUXB2DL port map( A0 => N3121, A1 => N3120, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1049);
   mult_21_C243_U1087 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1049, Z => 
                           mult_21_C243_n1352);
   mult_21_C243_U1086 : MUXB2DL port map( A0 => N3122, A1 => N3121, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1048);
   mult_21_C243_U1085 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1048, Z => 
                           mult_21_C243_n1351);
   mult_21_C243_U1084 : MUXB2DL port map( A0 => N3123, A1 => N3122, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1047);
   mult_21_C243_U1083 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1047, Z => 
                           mult_21_C243_n1350);
   mult_21_C243_U1082 : MUXB2DL port map( A0 => N3124, A1 => N3123, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1046);
   mult_21_C243_U1081 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1046, Z => 
                           mult_21_C243_n1349);
   mult_21_C243_U1080 : MUXB2DL port map( A0 => N3125, A1 => N3124, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1045);
   mult_21_C243_U1079 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1045, Z => 
                           mult_21_C243_n1348);
   mult_21_C243_U1078 : MUXB2DL port map( A0 => N3126, A1 => N3125, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1044);
   mult_21_C243_U1077 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1044, Z => 
                           mult_21_C243_n1347);
   mult_21_C243_U1076 : MUXB2DL port map( A0 => N3127, A1 => N3126, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1043);
   mult_21_C243_U1075 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1043, Z => 
                           mult_21_C243_n1346);
   mult_21_C243_U1074 : MUXB2DL port map( A0 => N3128, A1 => N3127, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1042);
   mult_21_C243_U1073 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1042, Z => 
                           mult_21_C243_n1345);
   mult_21_C243_U1072 : MUXB2DL port map( A0 => N3129, A1 => N3128, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1041);
   mult_21_C243_U1071 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1041, Z => 
                           mult_21_C243_n1344);
   mult_21_C243_U1070 : MUXB2DL port map( A0 => N3130, A1 => N3129, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1040);
   mult_21_C243_U1069 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1040, Z => 
                           mult_21_C243_n1343);
   mult_21_C243_U1068 : MUXB2DL port map( A0 => N3131, A1 => N3130, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1039);
   mult_21_C243_U1067 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1039, Z => 
                           mult_21_C243_n1342);
   mult_21_C243_U1066 : MUXB2DL port map( A0 => N3132, A1 => N3131, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1038);
   mult_21_C243_U1065 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1038, Z => 
                           mult_21_C243_n1341);
   mult_21_C243_U1064 : MUXB2DL port map( A0 => N3133, A1 => N3132, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1037);
   mult_21_C243_U1063 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1037, Z => 
                           mult_21_C243_n1340);
   mult_21_C243_U1062 : MUXB2DL port map( A0 => N3134, A1 => N3133, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1036);
   mult_21_C243_U1061 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1036, Z => 
                           mult_21_C243_n1339);
   mult_21_C243_U1060 : MUXB2DL port map( A0 => N3135, A1 => N3134, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1035);
   mult_21_C243_U1059 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1035, Z => 
                           mult_21_C243_n1338);
   mult_21_C243_U1058 : MUXB2DL port map( A0 => N3136, A1 => N3135, SL => 
                           mult_21_C243_n8, Z => mult_21_C243_n1034);
   mult_21_C243_U1057 : MUXB2DL port map( A0 => mult_21_C243_n3, A1 => 
                           mult_21_C243_n6, SL => mult_21_C243_n1034, Z => 
                           mult_21_C243_n1337);
   mult_21_C243_U1056 : NOR2M1D1 port map( A1 => mult_21_C243_n3, A2 => 
                           mult_21_C243_n6, Z => mult_21_C243_n1096);
   mult_21_C243_U1055 : NAN2M1D1 port map( A1 => mult_21_C243_n1542, A2 => 
                           N3105, Z => mult_21_C243_n1033);
   mult_21_C243_U1054 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1033, Z => 
                           mult_21_C243_n1336);
   mult_21_C243_U1053 : MUXB2DL port map( A0 => N3106, A1 => N3105, SL => 
                           mult_21_C243_n1542, Z => mult_21_C243_n1032);
   mult_21_C243_U1052 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1032, Z => 
                           mult_21_C243_n1335);
   mult_21_C243_U1051 : MUXB2DL port map( A0 => N3107, A1 => mult_21_C243_n1545
                           , SL => mult_21_C243_n1542, Z => mult_21_C243_n1031)
                           ;
   mult_21_C243_U1050 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1031, Z => 
                           mult_21_C243_n1334);
   mult_21_C243_U1049 : MUXB2DL port map( A0 => N3108, A1 => N3107, SL => 
                           mult_21_C243_n1542, Z => mult_21_C243_n1030);
   mult_21_C243_U1048 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1030, Z => 
                           mult_21_C243_n1333);
   mult_21_C243_U1047 : MUXB2DL port map( A0 => N3109, A1 => mult_21_C243_n1543
                           , SL => mult_21_C243_n1542, Z => mult_21_C243_n1029)
                           ;
   mult_21_C243_U1046 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1029, Z => 
                           mult_21_C243_n1332);
   mult_21_C243_U1045 : MUXB2DL port map( A0 => N3110, A1 => N3109, SL => 
                           mult_21_C243_n1542, Z => mult_21_C243_n1028);
   mult_21_C243_U1044 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1028, Z => 
                           mult_21_C243_n1331);
   mult_21_C243_U1043 : MUXB2DL port map( A0 => N3111, A1 => N3110, SL => 
                           mult_21_C243_n1542, Z => mult_21_C243_n1027);
   mult_21_C243_U1042 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1027, Z => 
                           mult_21_C243_n1330);
   mult_21_C243_U1041 : MUXB2DL port map( A0 => N3112, A1 => N3111, SL => 
                           mult_21_C243_n1542, Z => mult_21_C243_n1026);
   mult_21_C243_U1040 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1026, Z => 
                           mult_21_C243_n1329);
   mult_21_C243_U1039 : MUXB2DL port map( A0 => N3113, A1 => N3112, SL => 
                           mult_21_C243_n1542, Z => mult_21_C243_n1025);
   mult_21_C243_U1038 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1025, Z => 
                           mult_21_C243_n1328);
   mult_21_C243_U1037 : MUXB2DL port map( A0 => N3114, A1 => N3113, SL => 
                           mult_21_C243_n1542, Z => mult_21_C243_n1024);
   mult_21_C243_U1036 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1024, Z => 
                           mult_21_C243_n1327);
   mult_21_C243_U1035 : MUXB2DL port map( A0 => N3115, A1 => N3114, SL => 
                           mult_21_C243_n1542, Z => mult_21_C243_n1023);
   mult_21_C243_U1034 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1023, Z => 
                           mult_21_C243_n1326);
   mult_21_C243_U1033 : MUXB2DL port map( A0 => N3116, A1 => N3115, SL => 
                           mult_21_C243_n1542, Z => mult_21_C243_n1022);
   mult_21_C243_U1032 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1022, Z => 
                           mult_21_C243_n1325);
   mult_21_C243_U1031 : MUXB2DL port map( A0 => N3117, A1 => N3116, SL => 
                           mult_21_C243_n1542, Z => mult_21_C243_n1021);
   mult_21_C243_U1030 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1021, Z => 
                           mult_21_C243_n1324);
   mult_21_C243_U1029 : MUXB2DL port map( A0 => N3118, A1 => N3117, SL => 
                           mult_21_C243_n1542, Z => mult_21_C243_n1020);
   mult_21_C243_U1028 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1020, Z => 
                           mult_21_C243_n1323);
   mult_21_C243_U1027 : MUXB2DL port map( A0 => N3119, A1 => N3118, SL => 
                           mult_21_C243_n1542, Z => mult_21_C243_n1019);
   mult_21_C243_U1026 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1019, Z => 
                           mult_21_C243_n1322);
   mult_21_C243_U1025 : MUXB2DL port map( A0 => N3120, A1 => N3119, SL => 
                           mult_21_C243_n1542, Z => mult_21_C243_n1018);
   mult_21_C243_U1024 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1018, Z => 
                           mult_21_C243_n1321);
   mult_21_C243_U1023 : MUXB2DL port map( A0 => N3121, A1 => N3120, SL => 
                           mult_21_C243_n1542, Z => mult_21_C243_n1017);
   mult_21_C243_U1022 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1017, Z => 
                           mult_21_C243_n1320);
   mult_21_C243_U1021 : MUXB2DL port map( A0 => N3122, A1 => N3121, SL => 
                           mult_21_C243_n1542, Z => mult_21_C243_n1016);
   mult_21_C243_U1020 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1016, Z => 
                           mult_21_C243_n1319);
   mult_21_C243_U1019 : MUXB2DL port map( A0 => N3123, A1 => N3122, SL => 
                           mult_21_C243_n1542, Z => mult_21_C243_n1015);
   mult_21_C243_U1018 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1015, Z => 
                           mult_21_C243_n1318);
   mult_21_C243_U1017 : MUXB2DL port map( A0 => N3124, A1 => N3123, SL => 
                           mult_21_C243_n1542, Z => mult_21_C243_n1014);
   mult_21_C243_U1016 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1014, Z => 
                           mult_21_C243_n1317);
   mult_21_C243_U1015 : MUXB2DL port map( A0 => N3125, A1 => N3124, SL => 
                           mult_21_C243_n1542, Z => mult_21_C243_n1013);
   mult_21_C243_U1014 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1013, Z => 
                           mult_21_C243_n1316);
   mult_21_C243_U1013 : MUXB2DL port map( A0 => N3126, A1 => N3125, SL => 
                           mult_21_C243_n1542, Z => mult_21_C243_n1012);
   mult_21_C243_U1012 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1012, Z => 
                           mult_21_C243_n1315);
   mult_21_C243_U1011 : MUXB2DL port map( A0 => N3127, A1 => N3126, SL => 
                           mult_21_C243_n1542, Z => mult_21_C243_n1011);
   mult_21_C243_U1010 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1011, Z => 
                           mult_21_C243_n1314);
   mult_21_C243_U1009 : MUXB2DL port map( A0 => N3128, A1 => N3127, SL => 
                           mult_21_C243_n1542, Z => mult_21_C243_n1010);
   mult_21_C243_U1008 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1010, Z => 
                           mult_21_C243_n1313);
   mult_21_C243_U1007 : MUXB2DL port map( A0 => N3129, A1 => N3128, SL => 
                           mult_21_C243_n1542, Z => mult_21_C243_n1009);
   mult_21_C243_U1006 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1009, Z => 
                           mult_21_C243_n1312);
   mult_21_C243_U1005 : MUXB2DL port map( A0 => N3130, A1 => N3129, SL => 
                           mult_21_C243_n1542, Z => mult_21_C243_n1008);
   mult_21_C243_U1004 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1008, Z => 
                           mult_21_C243_n1311);
   mult_21_C243_U1003 : MUXB2DL port map( A0 => N3131, A1 => N3130, SL => 
                           mult_21_C243_n1542, Z => mult_21_C243_n1007);
   mult_21_C243_U1002 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1007, Z => 
                           mult_21_C243_n1310);
   mult_21_C243_U1001 : MUXB2DL port map( A0 => N3132, A1 => N3131, SL => 
                           mult_21_C243_n1542, Z => mult_21_C243_n1006);
   mult_21_C243_U1000 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1006, Z => 
                           mult_21_C243_n1309);
   mult_21_C243_U999 : MUXB2DL port map( A0 => N3133, A1 => N3132, SL => 
                           mult_21_C243_n1542, Z => mult_21_C243_n1005);
   mult_21_C243_U998 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1005, Z => 
                           mult_21_C243_n1308);
   mult_21_C243_U997 : MUXB2DL port map( A0 => N3134, A1 => N3133, SL => 
                           mult_21_C243_n1542, Z => mult_21_C243_n1004);
   mult_21_C243_U996 : MUXB2DL port map( A0 => mult_21_C243_n1517, A1 => 
                           mult_21_C243_n14, SL => mult_21_C243_n1004, Z => 
                           mult_21_C243_n1307);
   mult_21_C243_U995 : NOR2M1D1 port map( A1 => mult_21_C243_n1517, A2 => 
                           mult_21_C243_n14, Z => mult_21_C243_n1095);
   mult_21_C243_U994 : NAN2M1D1 port map( A1 => mult_21_C243_n1541, A2 => N3105
                           , Z => mult_21_C243_n1003);
   mult_21_C243_U993 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n1003, Z => 
                           mult_21_C243_n1306);
   mult_21_C243_U992 : MUXB2DL port map( A0 => N3106, A1 => N3105, SL => 
                           mult_21_C243_n1541, Z => mult_21_C243_n1002);
   mult_21_C243_U991 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n1002, Z => 
                           mult_21_C243_n1305);
   mult_21_C243_U990 : MUXB2DL port map( A0 => N3107, A1 => mult_21_C243_n1545,
                           SL => mult_21_C243_n1541, Z => mult_21_C243_n1001);
   mult_21_C243_U989 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n1001, Z => 
                           mult_21_C243_n1304);
   mult_21_C243_U988 : MUXB2DL port map( A0 => N3108, A1 => N3107, SL => 
                           mult_21_C243_n1541, Z => mult_21_C243_n1000);
   mult_21_C243_U987 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n1000, Z => 
                           mult_21_C243_n1303);
   mult_21_C243_U986 : MUXB2DL port map( A0 => N3109, A1 => mult_21_C243_n1543,
                           SL => mult_21_C243_n1541, Z => mult_21_C243_n999);
   mult_21_C243_U985 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n999, Z => 
                           mult_21_C243_n1302);
   mult_21_C243_U984 : MUXB2DL port map( A0 => N3110, A1 => N3109, SL => 
                           mult_21_C243_n1541, Z => mult_21_C243_n998);
   mult_21_C243_U983 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n998, Z => 
                           mult_21_C243_n1301);
   mult_21_C243_U982 : MUXB2DL port map( A0 => N3111, A1 => N3110, SL => 
                           mult_21_C243_n1541, Z => mult_21_C243_n997);
   mult_21_C243_U981 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n997, Z => 
                           mult_21_C243_n1300);
   mult_21_C243_U980 : MUXB2DL port map( A0 => N3112, A1 => N3111, SL => 
                           mult_21_C243_n1541, Z => mult_21_C243_n996);
   mult_21_C243_U979 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n996, Z => 
                           mult_21_C243_n1299);
   mult_21_C243_U978 : MUXB2DL port map( A0 => N3113, A1 => N3112, SL => 
                           mult_21_C243_n1541, Z => mult_21_C243_n995);
   mult_21_C243_U977 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n995, Z => 
                           mult_21_C243_n1298);
   mult_21_C243_U976 : MUXB2DL port map( A0 => N3114, A1 => N3113, SL => 
                           mult_21_C243_n1541, Z => mult_21_C243_n994);
   mult_21_C243_U975 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n994, Z => 
                           mult_21_C243_n1297);
   mult_21_C243_U974 : MUXB2DL port map( A0 => N3115, A1 => N3114, SL => 
                           mult_21_C243_n1541, Z => mult_21_C243_n993);
   mult_21_C243_U973 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n993, Z => 
                           mult_21_C243_n1296);
   mult_21_C243_U972 : MUXB2DL port map( A0 => N3116, A1 => N3115, SL => 
                           mult_21_C243_n1541, Z => mult_21_C243_n992);
   mult_21_C243_U971 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n992, Z => 
                           mult_21_C243_n1295);
   mult_21_C243_U970 : MUXB2DL port map( A0 => N3117, A1 => N3116, SL => 
                           mult_21_C243_n1541, Z => mult_21_C243_n991);
   mult_21_C243_U969 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n991, Z => 
                           mult_21_C243_n1294);
   mult_21_C243_U968 : MUXB2DL port map( A0 => N3118, A1 => N3117, SL => 
                           mult_21_C243_n1541, Z => mult_21_C243_n990);
   mult_21_C243_U967 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n990, Z => 
                           mult_21_C243_n1293);
   mult_21_C243_U966 : MUXB2DL port map( A0 => N3119, A1 => N3118, SL => 
                           mult_21_C243_n1541, Z => mult_21_C243_n989);
   mult_21_C243_U965 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n989, Z => 
                           mult_21_C243_n1292);
   mult_21_C243_U964 : MUXB2DL port map( A0 => N3120, A1 => N3119, SL => 
                           mult_21_C243_n1541, Z => mult_21_C243_n988);
   mult_21_C243_U963 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n988, Z => 
                           mult_21_C243_n1291);
   mult_21_C243_U962 : MUXB2DL port map( A0 => N3121, A1 => N3120, SL => 
                           mult_21_C243_n1541, Z => mult_21_C243_n987);
   mult_21_C243_U961 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n987, Z => 
                           mult_21_C243_n1290);
   mult_21_C243_U960 : MUXB2DL port map( A0 => N3122, A1 => N3121, SL => 
                           mult_21_C243_n1541, Z => mult_21_C243_n986);
   mult_21_C243_U959 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n986, Z => 
                           mult_21_C243_n1289);
   mult_21_C243_U958 : MUXB2DL port map( A0 => N3123, A1 => N3122, SL => 
                           mult_21_C243_n1541, Z => mult_21_C243_n985);
   mult_21_C243_U957 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n985, Z => 
                           mult_21_C243_n1288);
   mult_21_C243_U956 : MUXB2DL port map( A0 => N3124, A1 => N3123, SL => 
                           mult_21_C243_n1541, Z => mult_21_C243_n984);
   mult_21_C243_U955 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n984, Z => 
                           mult_21_C243_n1287);
   mult_21_C243_U954 : MUXB2DL port map( A0 => N3125, A1 => N3124, SL => 
                           mult_21_C243_n1541, Z => mult_21_C243_n983);
   mult_21_C243_U953 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n983, Z => 
                           mult_21_C243_n1286);
   mult_21_C243_U952 : MUXB2DL port map( A0 => N3126, A1 => N3125, SL => 
                           mult_21_C243_n1541, Z => mult_21_C243_n982);
   mult_21_C243_U951 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n982, Z => 
                           mult_21_C243_n1285);
   mult_21_C243_U950 : MUXB2DL port map( A0 => N3127, A1 => N3126, SL => 
                           mult_21_C243_n1541, Z => mult_21_C243_n981);
   mult_21_C243_U949 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n981, Z => 
                           mult_21_C243_n1284);
   mult_21_C243_U948 : MUXB2DL port map( A0 => N3128, A1 => N3127, SL => 
                           mult_21_C243_n1541, Z => mult_21_C243_n980);
   mult_21_C243_U947 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n980, Z => 
                           mult_21_C243_n1283);
   mult_21_C243_U946 : MUXB2DL port map( A0 => N3129, A1 => N3128, SL => 
                           mult_21_C243_n1541, Z => mult_21_C243_n979);
   mult_21_C243_U945 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n979, Z => 
                           mult_21_C243_n1282);
   mult_21_C243_U944 : MUXB2DL port map( A0 => N3130, A1 => N3129, SL => 
                           mult_21_C243_n1541, Z => mult_21_C243_n978);
   mult_21_C243_U943 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n978, Z => 
                           mult_21_C243_n1281);
   mult_21_C243_U942 : MUXB2DL port map( A0 => N3131, A1 => N3130, SL => 
                           mult_21_C243_n1541, Z => mult_21_C243_n977);
   mult_21_C243_U941 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n977, Z => 
                           mult_21_C243_n1280);
   mult_21_C243_U940 : MUXB2DL port map( A0 => N3132, A1 => N3131, SL => 
                           mult_21_C243_n1541, Z => mult_21_C243_n976);
   mult_21_C243_U939 : MUXB2DL port map( A0 => mult_21_C243_n1518, A1 => 
                           mult_21_C243_n22, SL => mult_21_C243_n976, Z => 
                           mult_21_C243_n1279);
   mult_21_C243_U938 : NOR2M1D1 port map( A1 => mult_21_C243_n1518, A2 => 
                           mult_21_C243_n22, Z => mult_21_C243_n1094);
   mult_21_C243_U937 : NAN2M1D1 port map( A1 => mult_21_C243_n1539, A2 => N3105
                           , Z => mult_21_C243_n975);
   mult_21_C243_U936 : MUXB2DL port map( A0 => mult_21_C243_n1540, A1 => 
                           mult_21_C243_n30, SL => mult_21_C243_n975, Z => 
                           mult_21_C243_n1278);
   mult_21_C243_U935 : MUXB2DL port map( A0 => N3106, A1 => N3105, SL => 
                           mult_21_C243_n1539, Z => mult_21_C243_n974);
   mult_21_C243_U934 : MUXB2DL port map( A0 => mult_21_C243_n1540, A1 => 
                           mult_21_C243_n30, SL => mult_21_C243_n974, Z => 
                           mult_21_C243_n1277);
   mult_21_C243_U933 : MUXB2DL port map( A0 => N3107, A1 => mult_21_C243_n1545,
                           SL => mult_21_C243_n1539, Z => mult_21_C243_n973);
   mult_21_C243_U932 : MUXB2DL port map( A0 => mult_21_C243_n1540, A1 => 
                           mult_21_C243_n30, SL => mult_21_C243_n973, Z => 
                           mult_21_C243_n1276);
   mult_21_C243_U931 : MUXB2DL port map( A0 => N3108, A1 => N3107, SL => 
                           mult_21_C243_n1539, Z => mult_21_C243_n972);
   mult_21_C243_U930 : MUXB2DL port map( A0 => mult_21_C243_n1540, A1 => 
                           mult_21_C243_n30, SL => mult_21_C243_n972, Z => 
                           mult_21_C243_n1275);
   mult_21_C243_U929 : MUXB2DL port map( A0 => N3109, A1 => N3108, SL => 
                           mult_21_C243_n1539, Z => mult_21_C243_n971);
   mult_21_C243_U928 : MUXB2DL port map( A0 => mult_21_C243_n1540, A1 => 
                           mult_21_C243_n30, SL => mult_21_C243_n971, Z => 
                           mult_21_C243_n1274);
   mult_21_C243_U927 : MUXB2DL port map( A0 => N3110, A1 => N3109, SL => 
                           mult_21_C243_n1539, Z => mult_21_C243_n970);
   mult_21_C243_U926 : MUXB2DL port map( A0 => mult_21_C243_n1540, A1 => 
                           mult_21_C243_n30, SL => mult_21_C243_n970, Z => 
                           mult_21_C243_n1273);
   mult_21_C243_U925 : MUXB2DL port map( A0 => N3111, A1 => N3110, SL => 
                           mult_21_C243_n1539, Z => mult_21_C243_n969);
   mult_21_C243_U924 : MUXB2DL port map( A0 => mult_21_C243_n1540, A1 => 
                           mult_21_C243_n30, SL => mult_21_C243_n969, Z => 
                           mult_21_C243_n1272);
   mult_21_C243_U923 : MUXB2DL port map( A0 => N3112, A1 => N3111, SL => 
                           mult_21_C243_n1539, Z => mult_21_C243_n968);
   mult_21_C243_U922 : MUXB2DL port map( A0 => mult_21_C243_n1540, A1 => 
                           mult_21_C243_n30, SL => mult_21_C243_n968, Z => 
                           mult_21_C243_n1271);
   mult_21_C243_U921 : MUXB2DL port map( A0 => N3113, A1 => N3112, SL => 
                           mult_21_C243_n1539, Z => mult_21_C243_n967);
   mult_21_C243_U920 : MUXB2DL port map( A0 => mult_21_C243_n1540, A1 => 
                           mult_21_C243_n30, SL => mult_21_C243_n967, Z => 
                           mult_21_C243_n1270);
   mult_21_C243_U919 : MUXB2DL port map( A0 => N3114, A1 => N3113, SL => 
                           mult_21_C243_n1539, Z => mult_21_C243_n966);
   mult_21_C243_U918 : MUXB2DL port map( A0 => mult_21_C243_n1540, A1 => 
                           mult_21_C243_n30, SL => mult_21_C243_n966, Z => 
                           mult_21_C243_n1269);
   mult_21_C243_U917 : MUXB2DL port map( A0 => N3115, A1 => N3114, SL => 
                           mult_21_C243_n1539, Z => mult_21_C243_n965);
   mult_21_C243_U916 : MUXB2DL port map( A0 => mult_21_C243_n1540, A1 => 
                           mult_21_C243_n30, SL => mult_21_C243_n965, Z => 
                           mult_21_C243_n1268);
   mult_21_C243_U915 : MUXB2DL port map( A0 => N3116, A1 => N3115, SL => 
                           mult_21_C243_n1539, Z => mult_21_C243_n964);
   mult_21_C243_U914 : MUXB2DL port map( A0 => mult_21_C243_n1540, A1 => 
                           mult_21_C243_n30, SL => mult_21_C243_n964, Z => 
                           mult_21_C243_n1267);
   mult_21_C243_U913 : MUXB2DL port map( A0 => N3117, A1 => N3116, SL => 
                           mult_21_C243_n1539, Z => mult_21_C243_n963);
   mult_21_C243_U912 : MUXB2DL port map( A0 => mult_21_C243_n1540, A1 => 
                           mult_21_C243_n30, SL => mult_21_C243_n963, Z => 
                           mult_21_C243_n1266);
   mult_21_C243_U911 : MUXB2DL port map( A0 => N3118, A1 => N3117, SL => 
                           mult_21_C243_n1539, Z => mult_21_C243_n962);
   mult_21_C243_U910 : MUXB2DL port map( A0 => mult_21_C243_n1540, A1 => 
                           mult_21_C243_n30, SL => mult_21_C243_n962, Z => 
                           mult_21_C243_n1265);
   mult_21_C243_U909 : MUXB2DL port map( A0 => N3119, A1 => N3118, SL => 
                           mult_21_C243_n1539, Z => mult_21_C243_n961);
   mult_21_C243_U908 : MUXB2DL port map( A0 => mult_21_C243_n1540, A1 => 
                           mult_21_C243_n30, SL => mult_21_C243_n961, Z => 
                           mult_21_C243_n1264);
   mult_21_C243_U907 : MUXB2DL port map( A0 => N3120, A1 => N3119, SL => 
                           mult_21_C243_n1539, Z => mult_21_C243_n960);
   mult_21_C243_U906 : MUXB2DL port map( A0 => mult_21_C243_n1540, A1 => 
                           mult_21_C243_n30, SL => mult_21_C243_n960, Z => 
                           mult_21_C243_n1263);
   mult_21_C243_U905 : MUXB2DL port map( A0 => N3121, A1 => N3120, SL => 
                           mult_21_C243_n1539, Z => mult_21_C243_n959);
   mult_21_C243_U904 : MUXB2DL port map( A0 => mult_21_C243_n1540, A1 => 
                           mult_21_C243_n30, SL => mult_21_C243_n959, Z => 
                           mult_21_C243_n1262);
   mult_21_C243_U903 : MUXB2DL port map( A0 => N3122, A1 => N3121, SL => 
                           mult_21_C243_n1539, Z => mult_21_C243_n958);
   mult_21_C243_U902 : MUXB2DL port map( A0 => mult_21_C243_n1540, A1 => 
                           mult_21_C243_n30, SL => mult_21_C243_n958, Z => 
                           mult_21_C243_n1261);
   mult_21_C243_U901 : MUXB2DL port map( A0 => N3123, A1 => N3122, SL => 
                           mult_21_C243_n1539, Z => mult_21_C243_n957);
   mult_21_C243_U900 : MUXB2DL port map( A0 => mult_21_C243_n1540, A1 => 
                           mult_21_C243_n30, SL => mult_21_C243_n957, Z => 
                           mult_21_C243_n1260);
   mult_21_C243_U899 : MUXB2DL port map( A0 => N3124, A1 => N3123, SL => 
                           mult_21_C243_n1539, Z => mult_21_C243_n956);
   mult_21_C243_U898 : MUXB2DL port map( A0 => mult_21_C243_n1540, A1 => 
                           mult_21_C243_n30, SL => mult_21_C243_n956, Z => 
                           mult_21_C243_n1259);
   mult_21_C243_U897 : MUXB2DL port map( A0 => N3125, A1 => N3124, SL => 
                           mult_21_C243_n1539, Z => mult_21_C243_n955);
   mult_21_C243_U896 : MUXB2DL port map( A0 => mult_21_C243_n1540, A1 => 
                           mult_21_C243_n30, SL => mult_21_C243_n955, Z => 
                           mult_21_C243_n1258);
   mult_21_C243_U895 : MUXB2DL port map( A0 => N3126, A1 => N3125, SL => 
                           mult_21_C243_n1539, Z => mult_21_C243_n954);
   mult_21_C243_U894 : MUXB2DL port map( A0 => mult_21_C243_n1540, A1 => 
                           mult_21_C243_n30, SL => mult_21_C243_n954, Z => 
                           mult_21_C243_n1257);
   mult_21_C243_U893 : MUXB2DL port map( A0 => N3127, A1 => N3126, SL => 
                           mult_21_C243_n1539, Z => mult_21_C243_n953);
   mult_21_C243_U892 : MUXB2DL port map( A0 => mult_21_C243_n1540, A1 => 
                           mult_21_C243_n30, SL => mult_21_C243_n953, Z => 
                           mult_21_C243_n1256);
   mult_21_C243_U891 : MUXB2DL port map( A0 => N3128, A1 => N3127, SL => 
                           mult_21_C243_n1539, Z => mult_21_C243_n952);
   mult_21_C243_U890 : MUXB2DL port map( A0 => mult_21_C243_n1540, A1 => 
                           mult_21_C243_n30, SL => mult_21_C243_n952, Z => 
                           mult_21_C243_n1255);
   mult_21_C243_U889 : MUXB2DL port map( A0 => N3129, A1 => N3128, SL => 
                           mult_21_C243_n1539, Z => mult_21_C243_n951);
   mult_21_C243_U888 : MUXB2DL port map( A0 => mult_21_C243_n1540, A1 => 
                           mult_21_C243_n30, SL => mult_21_C243_n951, Z => 
                           mult_21_C243_n1254);
   mult_21_C243_U887 : MUXB2DL port map( A0 => N3130, A1 => N3129, SL => 
                           mult_21_C243_n1539, Z => mult_21_C243_n950);
   mult_21_C243_U886 : MUXB2DL port map( A0 => mult_21_C243_n1540, A1 => 
                           mult_21_C243_n30, SL => mult_21_C243_n950, Z => 
                           mult_21_C243_n1253);
   mult_21_C243_U884 : NAN2M1D1 port map( A1 => mult_21_C243_n1538, A2 => N3105
                           , Z => mult_21_C243_n949);
   mult_21_C243_U883 : MUXB2DL port map( A0 => mult_21_C243_n1519, A1 => 
                           mult_21_C243_n38, SL => mult_21_C243_n949, Z => 
                           mult_21_C243_n1252);
   mult_21_C243_U882 : MUXB2DL port map( A0 => N3106, A1 => N3105, SL => 
                           mult_21_C243_n1538, Z => mult_21_C243_n948);
   mult_21_C243_U881 : MUXB2DL port map( A0 => mult_21_C243_n1519, A1 => 
                           mult_21_C243_n38, SL => mult_21_C243_n948, Z => 
                           mult_21_C243_n1251);
   mult_21_C243_U880 : MUXB2DL port map( A0 => N3107, A1 => mult_21_C243_n1545,
                           SL => mult_21_C243_n1538, Z => mult_21_C243_n947);
   mult_21_C243_U879 : MUXB2DL port map( A0 => mult_21_C243_n1519, A1 => 
                           mult_21_C243_n38, SL => mult_21_C243_n947, Z => 
                           mult_21_C243_n1250);
   mult_21_C243_U878 : MUXB2DL port map( A0 => N3108, A1 => N3107, SL => 
                           mult_21_C243_n1538, Z => mult_21_C243_n946);
   mult_21_C243_U877 : MUXB2DL port map( A0 => mult_21_C243_n1519, A1 => 
                           mult_21_C243_n38, SL => mult_21_C243_n946, Z => 
                           mult_21_C243_n1249);
   mult_21_C243_U876 : MUXB2DL port map( A0 => N3109, A1 => N3108, SL => 
                           mult_21_C243_n1538, Z => mult_21_C243_n945);
   mult_21_C243_U875 : MUXB2DL port map( A0 => mult_21_C243_n1519, A1 => 
                           mult_21_C243_n38, SL => mult_21_C243_n945, Z => 
                           mult_21_C243_n1248);
   mult_21_C243_U874 : MUXB2DL port map( A0 => N3110, A1 => N3109, SL => 
                           mult_21_C243_n1538, Z => mult_21_C243_n944);
   mult_21_C243_U873 : MUXB2DL port map( A0 => mult_21_C243_n1519, A1 => 
                           mult_21_C243_n38, SL => mult_21_C243_n944, Z => 
                           mult_21_C243_n1247);
   mult_21_C243_U872 : MUXB2DL port map( A0 => N3111, A1 => N3110, SL => 
                           mult_21_C243_n1538, Z => mult_21_C243_n943);
   mult_21_C243_U871 : MUXB2DL port map( A0 => mult_21_C243_n1519, A1 => 
                           mult_21_C243_n38, SL => mult_21_C243_n943, Z => 
                           mult_21_C243_n1246);
   mult_21_C243_U870 : MUXB2DL port map( A0 => N3112, A1 => N3111, SL => 
                           mult_21_C243_n1538, Z => mult_21_C243_n942);
   mult_21_C243_U869 : MUXB2DL port map( A0 => mult_21_C243_n1519, A1 => 
                           mult_21_C243_n38, SL => mult_21_C243_n942, Z => 
                           mult_21_C243_n1245);
   mult_21_C243_U868 : MUXB2DL port map( A0 => N3113, A1 => N3112, SL => 
                           mult_21_C243_n1538, Z => mult_21_C243_n941);
   mult_21_C243_U867 : MUXB2DL port map( A0 => mult_21_C243_n1519, A1 => 
                           mult_21_C243_n38, SL => mult_21_C243_n941, Z => 
                           mult_21_C243_n1244);
   mult_21_C243_U866 : MUXB2DL port map( A0 => N3114, A1 => N3113, SL => 
                           mult_21_C243_n1538, Z => mult_21_C243_n940);
   mult_21_C243_U865 : MUXB2DL port map( A0 => mult_21_C243_n1519, A1 => 
                           mult_21_C243_n38, SL => mult_21_C243_n940, Z => 
                           mult_21_C243_n1243);
   mult_21_C243_U864 : MUXB2DL port map( A0 => N3115, A1 => N3114, SL => 
                           mult_21_C243_n1538, Z => mult_21_C243_n939);
   mult_21_C243_U863 : MUXB2DL port map( A0 => mult_21_C243_n1519, A1 => 
                           mult_21_C243_n38, SL => mult_21_C243_n939, Z => 
                           mult_21_C243_n1242);
   mult_21_C243_U862 : MUXB2DL port map( A0 => N3116, A1 => N3115, SL => 
                           mult_21_C243_n1538, Z => mult_21_C243_n938);
   mult_21_C243_U861 : MUXB2DL port map( A0 => mult_21_C243_n1519, A1 => 
                           mult_21_C243_n38, SL => mult_21_C243_n938, Z => 
                           mult_21_C243_n1241);
   mult_21_C243_U860 : MUXB2DL port map( A0 => N3117, A1 => N3116, SL => 
                           mult_21_C243_n1538, Z => mult_21_C243_n937);
   mult_21_C243_U859 : MUXB2DL port map( A0 => mult_21_C243_n1519, A1 => 
                           mult_21_C243_n38, SL => mult_21_C243_n937, Z => 
                           mult_21_C243_n1240);
   mult_21_C243_U858 : MUXB2DL port map( A0 => N3118, A1 => N3117, SL => 
                           mult_21_C243_n1538, Z => mult_21_C243_n936);
   mult_21_C243_U857 : MUXB2DL port map( A0 => mult_21_C243_n1519, A1 => 
                           mult_21_C243_n38, SL => mult_21_C243_n936, Z => 
                           mult_21_C243_n1239);
   mult_21_C243_U856 : MUXB2DL port map( A0 => N3119, A1 => N3118, SL => 
                           mult_21_C243_n1538, Z => mult_21_C243_n935);
   mult_21_C243_U855 : MUXB2DL port map( A0 => mult_21_C243_n1519, A1 => 
                           mult_21_C243_n38, SL => mult_21_C243_n935, Z => 
                           mult_21_C243_n1238);
   mult_21_C243_U854 : MUXB2DL port map( A0 => N3120, A1 => N3119, SL => 
                           mult_21_C243_n1538, Z => mult_21_C243_n934);
   mult_21_C243_U853 : MUXB2DL port map( A0 => mult_21_C243_n1519, A1 => 
                           mult_21_C243_n38, SL => mult_21_C243_n934, Z => 
                           mult_21_C243_n1237);
   mult_21_C243_U852 : MUXB2DL port map( A0 => N3121, A1 => N3120, SL => 
                           mult_21_C243_n1538, Z => mult_21_C243_n933);
   mult_21_C243_U851 : MUXB2DL port map( A0 => mult_21_C243_n1519, A1 => 
                           mult_21_C243_n38, SL => mult_21_C243_n933, Z => 
                           mult_21_C243_n1236);
   mult_21_C243_U850 : MUXB2DL port map( A0 => N3122, A1 => N3121, SL => 
                           mult_21_C243_n1538, Z => mult_21_C243_n932);
   mult_21_C243_U849 : MUXB2DL port map( A0 => mult_21_C243_n1519, A1 => 
                           mult_21_C243_n38, SL => mult_21_C243_n932, Z => 
                           mult_21_C243_n1235);
   mult_21_C243_U848 : MUXB2DL port map( A0 => N3123, A1 => N3122, SL => 
                           mult_21_C243_n1538, Z => mult_21_C243_n931);
   mult_21_C243_U847 : MUXB2DL port map( A0 => mult_21_C243_n1519, A1 => 
                           mult_21_C243_n38, SL => mult_21_C243_n931, Z => 
                           mult_21_C243_n1234);
   mult_21_C243_U846 : MUXB2DL port map( A0 => N3124, A1 => N3123, SL => 
                           mult_21_C243_n1538, Z => mult_21_C243_n930);
   mult_21_C243_U845 : MUXB2DL port map( A0 => mult_21_C243_n1519, A1 => 
                           mult_21_C243_n38, SL => mult_21_C243_n930, Z => 
                           mult_21_C243_n1233);
   mult_21_C243_U844 : MUXB2DL port map( A0 => N3125, A1 => N3124, SL => 
                           mult_21_C243_n1538, Z => mult_21_C243_n929);
   mult_21_C243_U843 : MUXB2DL port map( A0 => mult_21_C243_n1519, A1 => 
                           mult_21_C243_n38, SL => mult_21_C243_n929, Z => 
                           mult_21_C243_n1232);
   mult_21_C243_U842 : MUXB2DL port map( A0 => N3126, A1 => N3125, SL => 
                           mult_21_C243_n1538, Z => mult_21_C243_n928);
   mult_21_C243_U841 : MUXB2DL port map( A0 => mult_21_C243_n1519, A1 => 
                           mult_21_C243_n38, SL => mult_21_C243_n928, Z => 
                           mult_21_C243_n1231);
   mult_21_C243_U840 : MUXB2DL port map( A0 => N3127, A1 => N3126, SL => 
                           mult_21_C243_n1538, Z => mult_21_C243_n927);
   mult_21_C243_U839 : MUXB2DL port map( A0 => mult_21_C243_n1519, A1 => 
                           mult_21_C243_n38, SL => mult_21_C243_n927, Z => 
                           mult_21_C243_n1230);
   mult_21_C243_U838 : MUXB2DL port map( A0 => N3128, A1 => N3127, SL => 
                           mult_21_C243_n1538, Z => mult_21_C243_n926);
   mult_21_C243_U837 : MUXB2DL port map( A0 => mult_21_C243_n1519, A1 => 
                           mult_21_C243_n38, SL => mult_21_C243_n926, Z => 
                           mult_21_C243_n1229);
   mult_21_C243_U836 : NOR2M1D1 port map( A1 => mult_21_C243_n1519, A2 => 
                           mult_21_C243_n38, Z => mult_21_C243_n1092);
   mult_21_C243_U835 : NAN2M1D1 port map( A1 => mult_21_C243_n48, A2 => N3105, 
                           Z => mult_21_C243_n925);
   mult_21_C243_U834 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n45, SL => mult_21_C243_n925, Z => 
                           mult_21_C243_n1228);
   mult_21_C243_U833 : MUXB2DL port map( A0 => mult_21_C243_n1545, A1 => N3105,
                           SL => mult_21_C243_n48, Z => mult_21_C243_n924);
   mult_21_C243_U832 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n45, SL => mult_21_C243_n924, Z => 
                           mult_21_C243_n1227);
   mult_21_C243_U831 : MUXB2DL port map( A0 => N3107, A1 => mult_21_C243_n1545,
                           SL => mult_21_C243_n48, Z => mult_21_C243_n923);
   mult_21_C243_U830 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n45, SL => mult_21_C243_n923, Z => 
                           mult_21_C243_n1226);
   mult_21_C243_U829 : MUXB2DL port map( A0 => N3108, A1 => N3107, SL => 
                           mult_21_C243_n48, Z => mult_21_C243_n922);
   mult_21_C243_U828 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n45, SL => mult_21_C243_n922, Z => 
                           mult_21_C243_n1225);
   mult_21_C243_U827 : MUXB2DL port map( A0 => N3109, A1 => N3108, SL => 
                           mult_21_C243_n48, Z => mult_21_C243_n921);
   mult_21_C243_U826 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n45, SL => mult_21_C243_n921, Z => 
                           mult_21_C243_n1224);
   mult_21_C243_U825 : MUXB2DL port map( A0 => N3110, A1 => N3109, SL => 
                           mult_21_C243_n48, Z => mult_21_C243_n920);
   mult_21_C243_U824 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n45, SL => mult_21_C243_n920, Z => 
                           mult_21_C243_n1223);
   mult_21_C243_U823 : MUXB2DL port map( A0 => N3111, A1 => N3110, SL => 
                           mult_21_C243_n48, Z => mult_21_C243_n919);
   mult_21_C243_U822 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n45, SL => mult_21_C243_n919, Z => 
                           mult_21_C243_n1222);
   mult_21_C243_U821 : MUXB2DL port map( A0 => N3112, A1 => N3111, SL => 
                           mult_21_C243_n48, Z => mult_21_C243_n918);
   mult_21_C243_U820 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n45, SL => mult_21_C243_n918, Z => 
                           mult_21_C243_n1221);
   mult_21_C243_U819 : MUXB2DL port map( A0 => N3113, A1 => N3112, SL => 
                           mult_21_C243_n48, Z => mult_21_C243_n917);
   mult_21_C243_U818 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n45, SL => mult_21_C243_n917, Z => 
                           mult_21_C243_n1220);
   mult_21_C243_U817 : MUXB2DL port map( A0 => N3114, A1 => N3113, SL => 
                           mult_21_C243_n48, Z => mult_21_C243_n916);
   mult_21_C243_U816 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n45, SL => mult_21_C243_n916, Z => 
                           mult_21_C243_n1219);
   mult_21_C243_U815 : MUXB2DL port map( A0 => N3115, A1 => N3114, SL => 
                           mult_21_C243_n48, Z => mult_21_C243_n915);
   mult_21_C243_U814 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n45, SL => mult_21_C243_n915, Z => 
                           mult_21_C243_n1218);
   mult_21_C243_U813 : MUXB2DL port map( A0 => N3116, A1 => N3115, SL => 
                           mult_21_C243_n48, Z => mult_21_C243_n914);
   mult_21_C243_U812 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n45, SL => mult_21_C243_n914, Z => 
                           mult_21_C243_n1217);
   mult_21_C243_U811 : MUXB2DL port map( A0 => N3117, A1 => N3116, SL => 
                           mult_21_C243_n48, Z => mult_21_C243_n913);
   mult_21_C243_U810 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n45, SL => mult_21_C243_n913, Z => 
                           mult_21_C243_n1216);
   mult_21_C243_U809 : MUXB2DL port map( A0 => N3118, A1 => N3117, SL => 
                           mult_21_C243_n48, Z => mult_21_C243_n912);
   mult_21_C243_U808 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n45, SL => mult_21_C243_n912, Z => 
                           mult_21_C243_n1215);
   mult_21_C243_U807 : MUXB2DL port map( A0 => N3119, A1 => N3118, SL => 
                           mult_21_C243_n48, Z => mult_21_C243_n911);
   mult_21_C243_U806 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n45, SL => mult_21_C243_n911, Z => 
                           mult_21_C243_n1214);
   mult_21_C243_U805 : MUXB2DL port map( A0 => N3120, A1 => N3119, SL => 
                           mult_21_C243_n48, Z => mult_21_C243_n910);
   mult_21_C243_U804 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n45, SL => mult_21_C243_n910, Z => 
                           mult_21_C243_n1213);
   mult_21_C243_U803 : MUXB2DL port map( A0 => N3121, A1 => N3120, SL => 
                           mult_21_C243_n48, Z => mult_21_C243_n909);
   mult_21_C243_U802 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n45, SL => mult_21_C243_n909, Z => 
                           mult_21_C243_n1212);
   mult_21_C243_U801 : MUXB2DL port map( A0 => N3122, A1 => N3121, SL => 
                           mult_21_C243_n48, Z => mult_21_C243_n908);
   mult_21_C243_U800 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n45, SL => mult_21_C243_n908, Z => 
                           mult_21_C243_n1211);
   mult_21_C243_U799 : MUXB2DL port map( A0 => N3123, A1 => N3122, SL => 
                           mult_21_C243_n48, Z => mult_21_C243_n907);
   mult_21_C243_U798 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n45, SL => mult_21_C243_n907, Z => 
                           mult_21_C243_n1210);
   mult_21_C243_U797 : MUXB2DL port map( A0 => N3124, A1 => N3123, SL => 
                           mult_21_C243_n48, Z => mult_21_C243_n906);
   mult_21_C243_U796 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n45, SL => mult_21_C243_n906, Z => 
                           mult_21_C243_n1209);
   mult_21_C243_U795 : MUXB2DL port map( A0 => N3125, A1 => N3124, SL => 
                           mult_21_C243_n48, Z => mult_21_C243_n905);
   mult_21_C243_U794 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n45, SL => mult_21_C243_n905, Z => 
                           mult_21_C243_n1208);
   mult_21_C243_U793 : MUXB2DL port map( A0 => N3126, A1 => N3125, SL => 
                           mult_21_C243_n48, Z => mult_21_C243_n904);
   mult_21_C243_U792 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n45, SL => mult_21_C243_n904, Z => 
                           mult_21_C243_n1207);
   mult_21_C243_U791 : NOR2M1D1 port map( A1 => mult_21_C243_n42, A2 => 
                           mult_21_C243_n45, Z => mult_21_C243_n1091);
   mult_21_C243_U790 : NAN2M1D1 port map( A1 => mult_21_C243_n56, A2 => N3105, 
                           Z => mult_21_C243_n903);
   mult_21_C243_U789 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n53, SL => mult_21_C243_n903, Z => 
                           mult_21_C243_n1206);
   mult_21_C243_U788 : MUXB2DL port map( A0 => mult_21_C243_n1545, A1 => N3105,
                           SL => mult_21_C243_n56, Z => mult_21_C243_n902);
   mult_21_C243_U787 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n53, SL => mult_21_C243_n902, Z => 
                           mult_21_C243_n1205);
   mult_21_C243_U786 : MUXB2DL port map( A0 => N3107, A1 => mult_21_C243_n1545,
                           SL => mult_21_C243_n56, Z => mult_21_C243_n901);
   mult_21_C243_U785 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n53, SL => mult_21_C243_n901, Z => 
                           mult_21_C243_n1204);
   mult_21_C243_U784 : MUXB2DL port map( A0 => N3108, A1 => N3107, SL => 
                           mult_21_C243_n56, Z => mult_21_C243_n900);
   mult_21_C243_U783 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n53, SL => mult_21_C243_n900, Z => 
                           mult_21_C243_n1203);
   mult_21_C243_U782 : MUXB2DL port map( A0 => N3109, A1 => mult_21_C243_n1543,
                           SL => mult_21_C243_n56, Z => mult_21_C243_n899);
   mult_21_C243_U781 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n53, SL => mult_21_C243_n899, Z => 
                           mult_21_C243_n1202);
   mult_21_C243_U780 : MUXB2DL port map( A0 => N3110, A1 => N3109, SL => 
                           mult_21_C243_n56, Z => mult_21_C243_n898);
   mult_21_C243_U779 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n53, SL => mult_21_C243_n898, Z => 
                           mult_21_C243_n1201);
   mult_21_C243_U778 : MUXB2DL port map( A0 => N3111, A1 => N3110, SL => 
                           mult_21_C243_n56, Z => mult_21_C243_n897);
   mult_21_C243_U777 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n53, SL => mult_21_C243_n897, Z => 
                           mult_21_C243_n1200);
   mult_21_C243_U776 : MUXB2DL port map( A0 => N3112, A1 => N3111, SL => 
                           mult_21_C243_n56, Z => mult_21_C243_n896);
   mult_21_C243_U775 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n53, SL => mult_21_C243_n896, Z => 
                           mult_21_C243_n1199);
   mult_21_C243_U774 : MUXB2DL port map( A0 => N3113, A1 => N3112, SL => 
                           mult_21_C243_n56, Z => mult_21_C243_n895);
   mult_21_C243_U773 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n53, SL => mult_21_C243_n895, Z => 
                           mult_21_C243_n1198);
   mult_21_C243_U772 : MUXB2DL port map( A0 => N3114, A1 => N3113, SL => 
                           mult_21_C243_n56, Z => mult_21_C243_n894);
   mult_21_C243_U771 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n53, SL => mult_21_C243_n894, Z => 
                           mult_21_C243_n1197);
   mult_21_C243_U770 : MUXB2DL port map( A0 => N3115, A1 => N3114, SL => 
                           mult_21_C243_n56, Z => mult_21_C243_n893);
   mult_21_C243_U769 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n53, SL => mult_21_C243_n893, Z => 
                           mult_21_C243_n1196);
   mult_21_C243_U768 : MUXB2DL port map( A0 => N3116, A1 => N3115, SL => 
                           mult_21_C243_n56, Z => mult_21_C243_n892);
   mult_21_C243_U767 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n53, SL => mult_21_C243_n892, Z => 
                           mult_21_C243_n1195);
   mult_21_C243_U766 : MUXB2DL port map( A0 => N3117, A1 => N3116, SL => 
                           mult_21_C243_n56, Z => mult_21_C243_n891);
   mult_21_C243_U765 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n53, SL => mult_21_C243_n891, Z => 
                           mult_21_C243_n1194);
   mult_21_C243_U764 : MUXB2DL port map( A0 => N3118, A1 => N3117, SL => 
                           mult_21_C243_n56, Z => mult_21_C243_n890);
   mult_21_C243_U763 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n53, SL => mult_21_C243_n890, Z => 
                           mult_21_C243_n1193);
   mult_21_C243_U762 : MUXB2DL port map( A0 => N3119, A1 => N3118, SL => 
                           mult_21_C243_n56, Z => mult_21_C243_n889);
   mult_21_C243_U761 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n53, SL => mult_21_C243_n889, Z => 
                           mult_21_C243_n1192);
   mult_21_C243_U760 : MUXB2DL port map( A0 => N3120, A1 => N3119, SL => 
                           mult_21_C243_n56, Z => mult_21_C243_n888);
   mult_21_C243_U759 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n53, SL => mult_21_C243_n888, Z => 
                           mult_21_C243_n1191);
   mult_21_C243_U758 : MUXB2DL port map( A0 => N3121, A1 => N3120, SL => 
                           mult_21_C243_n56, Z => mult_21_C243_n887);
   mult_21_C243_U757 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n53, SL => mult_21_C243_n887, Z => 
                           mult_21_C243_n1190);
   mult_21_C243_U756 : MUXB2DL port map( A0 => N3122, A1 => N3121, SL => 
                           mult_21_C243_n56, Z => mult_21_C243_n886);
   mult_21_C243_U755 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n53, SL => mult_21_C243_n886, Z => 
                           mult_21_C243_n1189);
   mult_21_C243_U754 : MUXB2DL port map( A0 => N3123, A1 => N3122, SL => 
                           mult_21_C243_n56, Z => mult_21_C243_n885);
   mult_21_C243_U753 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n53, SL => mult_21_C243_n885, Z => 
                           mult_21_C243_n1188);
   mult_21_C243_U752 : MUXB2DL port map( A0 => N3124, A1 => N3123, SL => 
                           mult_21_C243_n56, Z => mult_21_C243_n884);
   mult_21_C243_U751 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n53, SL => mult_21_C243_n884, Z => 
                           mult_21_C243_n1187);
   mult_21_C243_U750 : NOR2M1D1 port map( A1 => mult_21_C243_n50, A2 => 
                           mult_21_C243_n53, Z => mult_21_C243_n1090);
   mult_21_C243_U749 : NAN2M1D1 port map( A1 => mult_21_C243_n63, A2 => N3105, 
                           Z => mult_21_C243_n883);
   mult_21_C243_U748 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n61, SL => mult_21_C243_n883, Z => 
                           mult_21_C243_n1186);
   mult_21_C243_U747 : MUXB2DL port map( A0 => mult_21_C243_n1545, A1 => N3105,
                           SL => mult_21_C243_n63, Z => mult_21_C243_n882);
   mult_21_C243_U746 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n61, SL => mult_21_C243_n882, Z => 
                           mult_21_C243_n1185);
   mult_21_C243_U745 : MUXB2DL port map( A0 => N3107, A1 => mult_21_C243_n1545,
                           SL => mult_21_C243_n63, Z => mult_21_C243_n881);
   mult_21_C243_U744 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n61, SL => mult_21_C243_n881, Z => 
                           mult_21_C243_n1184);
   mult_21_C243_U743 : MUXB2DL port map( A0 => N3108, A1 => N3107, SL => 
                           mult_21_C243_n63, Z => mult_21_C243_n880);
   mult_21_C243_U742 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n61, SL => mult_21_C243_n880, Z => 
                           mult_21_C243_n1183);
   mult_21_C243_U741 : MUXB2DL port map( A0 => N3109, A1 => mult_21_C243_n1543,
                           SL => mult_21_C243_n63, Z => mult_21_C243_n879);
   mult_21_C243_U740 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n61, SL => mult_21_C243_n879, Z => 
                           mult_21_C243_n1182);
   mult_21_C243_U739 : MUXB2DL port map( A0 => N3110, A1 => N3109, SL => 
                           mult_21_C243_n63, Z => mult_21_C243_n878);
   mult_21_C243_U738 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n61, SL => mult_21_C243_n878, Z => 
                           mult_21_C243_n1181);
   mult_21_C243_U737 : MUXB2DL port map( A0 => N3111, A1 => N3110, SL => 
                           mult_21_C243_n63, Z => mult_21_C243_n877);
   mult_21_C243_U736 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n61, SL => mult_21_C243_n877, Z => 
                           mult_21_C243_n1180);
   mult_21_C243_U735 : MUXB2DL port map( A0 => N3112, A1 => N3111, SL => 
                           mult_21_C243_n63, Z => mult_21_C243_n876);
   mult_21_C243_U734 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n61, SL => mult_21_C243_n876, Z => 
                           mult_21_C243_n1179);
   mult_21_C243_U733 : MUXB2DL port map( A0 => N3113, A1 => N3112, SL => 
                           mult_21_C243_n63, Z => mult_21_C243_n875);
   mult_21_C243_U732 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n61, SL => mult_21_C243_n875, Z => 
                           mult_21_C243_n1178);
   mult_21_C243_U731 : MUXB2DL port map( A0 => N3114, A1 => N3113, SL => 
                           mult_21_C243_n63, Z => mult_21_C243_n874);
   mult_21_C243_U730 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n61, SL => mult_21_C243_n874, Z => 
                           mult_21_C243_n1177);
   mult_21_C243_U729 : MUXB2DL port map( A0 => N3115, A1 => N3114, SL => 
                           mult_21_C243_n63, Z => mult_21_C243_n873);
   mult_21_C243_U728 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n61, SL => mult_21_C243_n873, Z => 
                           mult_21_C243_n1176);
   mult_21_C243_U727 : MUXB2DL port map( A0 => N3116, A1 => N3115, SL => 
                           mult_21_C243_n63, Z => mult_21_C243_n872);
   mult_21_C243_U726 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n61, SL => mult_21_C243_n872, Z => 
                           mult_21_C243_n1175);
   mult_21_C243_U725 : MUXB2DL port map( A0 => N3117, A1 => N3116, SL => 
                           mult_21_C243_n63, Z => mult_21_C243_n871);
   mult_21_C243_U724 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n61, SL => mult_21_C243_n871, Z => 
                           mult_21_C243_n1174);
   mult_21_C243_U723 : MUXB2DL port map( A0 => N3118, A1 => N3117, SL => 
                           mult_21_C243_n63, Z => mult_21_C243_n870);
   mult_21_C243_U722 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n61, SL => mult_21_C243_n870, Z => 
                           mult_21_C243_n1173);
   mult_21_C243_U721 : MUXB2DL port map( A0 => N3119, A1 => N3118, SL => 
                           mult_21_C243_n63, Z => mult_21_C243_n869);
   mult_21_C243_U720 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n61, SL => mult_21_C243_n869, Z => 
                           mult_21_C243_n1172);
   mult_21_C243_U719 : MUXB2DL port map( A0 => N3120, A1 => N3119, SL => 
                           mult_21_C243_n63, Z => mult_21_C243_n868);
   mult_21_C243_U718 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n61, SL => mult_21_C243_n868, Z => 
                           mult_21_C243_n1171);
   mult_21_C243_U717 : MUXB2DL port map( A0 => N3121, A1 => N3120, SL => 
                           mult_21_C243_n63, Z => mult_21_C243_n867);
   mult_21_C243_U716 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n61, SL => mult_21_C243_n867, Z => 
                           mult_21_C243_n1170);
   mult_21_C243_U715 : MUXB2DL port map( A0 => N3122, A1 => N3121, SL => 
                           mult_21_C243_n63, Z => mult_21_C243_n866);
   mult_21_C243_U714 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n61, SL => mult_21_C243_n866, Z => 
                           mult_21_C243_n1169);
   mult_21_C243_U713 : NOR2M1D1 port map( A1 => mult_21_C243_n58, A2 => 
                           mult_21_C243_n61, Z => mult_21_C243_n1089);
   mult_21_C243_U712 : NAN2M1D1 port map( A1 => mult_21_C243_n71, A2 => N3105, 
                           Z => mult_21_C243_n865);
   mult_21_C243_U711 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n69, SL => mult_21_C243_n865, Z => 
                           mult_21_C243_n1168);
   mult_21_C243_U710 : MUXB2DL port map( A0 => N3106, A1 => N3105, SL => 
                           mult_21_C243_n71, Z => mult_21_C243_n864);
   mult_21_C243_U709 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n69, SL => mult_21_C243_n864, Z => 
                           mult_21_C243_n1167);
   mult_21_C243_U708 : MUXB2DL port map( A0 => N3107, A1 => mult_21_C243_n1545,
                           SL => mult_21_C243_n71, Z => mult_21_C243_n863);
   mult_21_C243_U707 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n69, SL => mult_21_C243_n863, Z => 
                           mult_21_C243_n1166);
   mult_21_C243_U706 : MUXB2DL port map( A0 => mult_21_C243_n1543, A1 => N3107,
                           SL => mult_21_C243_n71, Z => mult_21_C243_n862);
   mult_21_C243_U705 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n69, SL => mult_21_C243_n862, Z => 
                           mult_21_C243_n1165);
   mult_21_C243_U704 : MUXB2DL port map( A0 => N3109, A1 => mult_21_C243_n1543,
                           SL => mult_21_C243_n71, Z => mult_21_C243_n861);
   mult_21_C243_U703 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n69, SL => mult_21_C243_n861, Z => 
                           mult_21_C243_n1164);
   mult_21_C243_U702 : MUXB2DL port map( A0 => N3110, A1 => N3109, SL => 
                           mult_21_C243_n71, Z => mult_21_C243_n860);
   mult_21_C243_U701 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n69, SL => mult_21_C243_n860, Z => 
                           mult_21_C243_n1163);
   mult_21_C243_U700 : MUXB2DL port map( A0 => N3111, A1 => N3110, SL => 
                           mult_21_C243_n71, Z => mult_21_C243_n859);
   mult_21_C243_U699 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n69, SL => mult_21_C243_n859, Z => 
                           mult_21_C243_n1162);
   mult_21_C243_U698 : MUXB2DL port map( A0 => N3112, A1 => N3111, SL => 
                           mult_21_C243_n71, Z => mult_21_C243_n858);
   mult_21_C243_U697 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n69, SL => mult_21_C243_n858, Z => 
                           mult_21_C243_n1161);
   mult_21_C243_U696 : MUXB2DL port map( A0 => N3113, A1 => N3112, SL => 
                           mult_21_C243_n71, Z => mult_21_C243_n857);
   mult_21_C243_U695 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n69, SL => mult_21_C243_n857, Z => 
                           mult_21_C243_n1160);
   mult_21_C243_U694 : MUXB2DL port map( A0 => N3114, A1 => N3113, SL => 
                           mult_21_C243_n71, Z => mult_21_C243_n856);
   mult_21_C243_U693 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n69, SL => mult_21_C243_n856, Z => 
                           mult_21_C243_n1159);
   mult_21_C243_U692 : MUXB2DL port map( A0 => N3115, A1 => N3114, SL => 
                           mult_21_C243_n71, Z => mult_21_C243_n855);
   mult_21_C243_U691 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n69, SL => mult_21_C243_n855, Z => 
                           mult_21_C243_n1158);
   mult_21_C243_U690 : MUXB2DL port map( A0 => N3116, A1 => N3115, SL => 
                           mult_21_C243_n71, Z => mult_21_C243_n854);
   mult_21_C243_U689 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n69, SL => mult_21_C243_n854, Z => 
                           mult_21_C243_n1157);
   mult_21_C243_U688 : MUXB2DL port map( A0 => N3117, A1 => N3116, SL => 
                           mult_21_C243_n71, Z => mult_21_C243_n853);
   mult_21_C243_U687 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n69, SL => mult_21_C243_n853, Z => 
                           mult_21_C243_n1156);
   mult_21_C243_U686 : MUXB2DL port map( A0 => N3118, A1 => N3117, SL => 
                           mult_21_C243_n71, Z => mult_21_C243_n852);
   mult_21_C243_U685 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n69, SL => mult_21_C243_n852, Z => 
                           mult_21_C243_n1155);
   mult_21_C243_U684 : MUXB2DL port map( A0 => N3119, A1 => N3118, SL => 
                           mult_21_C243_n71, Z => mult_21_C243_n851);
   mult_21_C243_U683 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n69, SL => mult_21_C243_n851, Z => 
                           mult_21_C243_n1154);
   mult_21_C243_U682 : MUXB2DL port map( A0 => N3120, A1 => N3119, SL => 
                           mult_21_C243_n71, Z => mult_21_C243_n850);
   mult_21_C243_U681 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n69, SL => mult_21_C243_n850, Z => 
                           mult_21_C243_n1153);
   mult_21_C243_U680 : NOR2M1D1 port map( A1 => mult_21_C243_n66, A2 => 
                           mult_21_C243_n69, Z => mult_21_C243_n1088);
   mult_21_C243_U679 : NAN2M1D1 port map( A1 => mult_21_C243_n78, A2 => N3105, 
                           Z => mult_21_C243_n849);
   mult_21_C243_U678 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n76, SL => mult_21_C243_n849, Z => 
                           mult_21_C243_n1152);
   mult_21_C243_U677 : MUXB2DL port map( A0 => N3106, A1 => N3105, SL => 
                           mult_21_C243_n78, Z => mult_21_C243_n848);
   mult_21_C243_U676 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n76, SL => mult_21_C243_n848, Z => 
                           mult_21_C243_n1151);
   mult_21_C243_U675 : MUXB2DL port map( A0 => N3107, A1 => mult_21_C243_n1545,
                           SL => mult_21_C243_n78, Z => mult_21_C243_n847);
   mult_21_C243_U674 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n76, SL => mult_21_C243_n847, Z => 
                           mult_21_C243_n1150);
   mult_21_C243_U673 : MUXB2DL port map( A0 => mult_21_C243_n1543, A1 => N3107,
                           SL => mult_21_C243_n78, Z => mult_21_C243_n846);
   mult_21_C243_U672 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n76, SL => mult_21_C243_n846, Z => 
                           mult_21_C243_n1149);
   mult_21_C243_U671 : MUXB2DL port map( A0 => N3109, A1 => mult_21_C243_n1543,
                           SL => mult_21_C243_n78, Z => mult_21_C243_n845);
   mult_21_C243_U670 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n76, SL => mult_21_C243_n845, Z => 
                           mult_21_C243_n1148);
   mult_21_C243_U669 : MUXB2DL port map( A0 => N3110, A1 => N3109, SL => 
                           mult_21_C243_n78, Z => mult_21_C243_n844);
   mult_21_C243_U668 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n76, SL => mult_21_C243_n844, Z => 
                           mult_21_C243_n1147);
   mult_21_C243_U667 : MUXB2DL port map( A0 => N3111, A1 => N3110, SL => 
                           mult_21_C243_n78, Z => mult_21_C243_n843);
   mult_21_C243_U666 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n76, SL => mult_21_C243_n843, Z => 
                           mult_21_C243_n1146);
   mult_21_C243_U665 : MUXB2DL port map( A0 => N3112, A1 => N3111, SL => 
                           mult_21_C243_n78, Z => mult_21_C243_n842);
   mult_21_C243_U664 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n76, SL => mult_21_C243_n842, Z => 
                           mult_21_C243_n1145);
   mult_21_C243_U663 : MUXB2DL port map( A0 => N3113, A1 => N3112, SL => 
                           mult_21_C243_n78, Z => mult_21_C243_n841);
   mult_21_C243_U662 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n76, SL => mult_21_C243_n841, Z => 
                           mult_21_C243_n1144);
   mult_21_C243_U661 : MUXB2DL port map( A0 => N3114, A1 => N3113, SL => 
                           mult_21_C243_n78, Z => mult_21_C243_n840);
   mult_21_C243_U660 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n76, SL => mult_21_C243_n840, Z => 
                           mult_21_C243_n1143);
   mult_21_C243_U659 : MUXB2DL port map( A0 => N3115, A1 => N3114, SL => 
                           mult_21_C243_n78, Z => mult_21_C243_n839);
   mult_21_C243_U658 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n76, SL => mult_21_C243_n839, Z => 
                           mult_21_C243_n1142);
   mult_21_C243_U657 : MUXB2DL port map( A0 => N3116, A1 => N3115, SL => 
                           mult_21_C243_n78, Z => mult_21_C243_n838);
   mult_21_C243_U656 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n76, SL => mult_21_C243_n838, Z => 
                           mult_21_C243_n1141);
   mult_21_C243_U655 : MUXB2DL port map( A0 => N3117, A1 => N3116, SL => 
                           mult_21_C243_n78, Z => mult_21_C243_n837);
   mult_21_C243_U654 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n76, SL => mult_21_C243_n837, Z => 
                           mult_21_C243_n1140);
   mult_21_C243_U653 : MUXB2DL port map( A0 => N3118, A1 => N3117, SL => 
                           mult_21_C243_n78, Z => mult_21_C243_n836);
   mult_21_C243_U652 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n76, SL => mult_21_C243_n836, Z => 
                           mult_21_C243_n1139);
   mult_21_C243_U651 : NOR2M1D1 port map( A1 => mult_21_C243_n73, A2 => 
                           mult_21_C243_n76, Z => mult_21_C243_n1087);
   mult_21_C243_U650 : NAN2M1D1 port map( A1 => mult_21_C243_n83, A2 => N3105, 
                           Z => mult_21_C243_n835);
   mult_21_C243_U649 : MUXB2DL port map( A0 => mult_21_C243_n79, A1 => 
                           mult_21_C243_n81, SL => mult_21_C243_n835, Z => 
                           mult_21_C243_n1138);
   mult_21_C243_U648 : MUXB2DL port map( A0 => N3106, A1 => N3105, SL => 
                           mult_21_C243_n83, Z => mult_21_C243_n834);
   mult_21_C243_U647 : MUXB2DL port map( A0 => mult_21_C243_n79, A1 => 
                           mult_21_C243_n81, SL => mult_21_C243_n834, Z => 
                           mult_21_C243_n1137);
   mult_21_C243_U646 : MUXB2DL port map( A0 => N3107, A1 => mult_21_C243_n1545,
                           SL => mult_21_C243_n83, Z => mult_21_C243_n833);
   mult_21_C243_U645 : MUXB2DL port map( A0 => mult_21_C243_n79, A1 => 
                           mult_21_C243_n81, SL => mult_21_C243_n833, Z => 
                           mult_21_C243_n1136);
   mult_21_C243_U644 : MUXB2DL port map( A0 => mult_21_C243_n1543, A1 => N3107,
                           SL => mult_21_C243_n83, Z => mult_21_C243_n832);
   mult_21_C243_U643 : MUXB2DL port map( A0 => mult_21_C243_n79, A1 => 
                           mult_21_C243_n81, SL => mult_21_C243_n832, Z => 
                           mult_21_C243_n1135);
   mult_21_C243_U642 : MUXB2DL port map( A0 => N3109, A1 => mult_21_C243_n1543,
                           SL => mult_21_C243_n83, Z => mult_21_C243_n831);
   mult_21_C243_U641 : MUXB2DL port map( A0 => mult_21_C243_n79, A1 => 
                           mult_21_C243_n81, SL => mult_21_C243_n831, Z => 
                           mult_21_C243_n1134);
   mult_21_C243_U640 : MUXB2DL port map( A0 => N3110, A1 => N3109, SL => 
                           mult_21_C243_n83, Z => mult_21_C243_n830);
   mult_21_C243_U639 : MUXB2DL port map( A0 => mult_21_C243_n79, A1 => 
                           mult_21_C243_n81, SL => mult_21_C243_n830, Z => 
                           mult_21_C243_n1133);
   mult_21_C243_U638 : MUXB2DL port map( A0 => N3111, A1 => N3110, SL => 
                           mult_21_C243_n83, Z => mult_21_C243_n829);
   mult_21_C243_U637 : MUXB2DL port map( A0 => mult_21_C243_n79, A1 => 
                           mult_21_C243_n81, SL => mult_21_C243_n829, Z => 
                           mult_21_C243_n1132);
   mult_21_C243_U636 : MUXB2DL port map( A0 => N3112, A1 => N3111, SL => 
                           mult_21_C243_n83, Z => mult_21_C243_n828);
   mult_21_C243_U635 : MUXB2DL port map( A0 => mult_21_C243_n79, A1 => 
                           mult_21_C243_n81, SL => mult_21_C243_n828, Z => 
                           mult_21_C243_n1131);
   mult_21_C243_U634 : MUXB2DL port map( A0 => N3113, A1 => N3112, SL => 
                           mult_21_C243_n83, Z => mult_21_C243_n827);
   mult_21_C243_U633 : MUXB2DL port map( A0 => mult_21_C243_n79, A1 => 
                           mult_21_C243_n81, SL => mult_21_C243_n827, Z => 
                           mult_21_C243_n1130);
   mult_21_C243_U632 : MUXB2DL port map( A0 => N3114, A1 => N3113, SL => 
                           mult_21_C243_n83, Z => mult_21_C243_n826);
   mult_21_C243_U631 : MUXB2DL port map( A0 => mult_21_C243_n79, A1 => 
                           mult_21_C243_n81, SL => mult_21_C243_n826, Z => 
                           mult_21_C243_n1129);
   mult_21_C243_U630 : MUXB2DL port map( A0 => N3115, A1 => N3114, SL => 
                           mult_21_C243_n83, Z => mult_21_C243_n825);
   mult_21_C243_U629 : MUXB2DL port map( A0 => mult_21_C243_n79, A1 => 
                           mult_21_C243_n81, SL => mult_21_C243_n825, Z => 
                           mult_21_C243_n1128);
   mult_21_C243_U628 : MUXB2DL port map( A0 => N3116, A1 => N3115, SL => 
                           mult_21_C243_n83, Z => mult_21_C243_n824);
   mult_21_C243_U627 : MUXB2DL port map( A0 => mult_21_C243_n79, A1 => 
                           mult_21_C243_n81, SL => mult_21_C243_n824, Z => 
                           mult_21_C243_n1127);
   mult_21_C243_U626 : NOR2M1D1 port map( A1 => mult_21_C243_n79, A2 => 
                           mult_21_C243_n81, Z => mult_21_C243_n1086);
   mult_21_C243_U625 : NAN2M1D1 port map( A1 => mult_21_C243_n88, A2 => N3105, 
                           Z => mult_21_C243_n823);
   mult_21_C243_U624 : MUXB2DL port map( A0 => mult_21_C243_n84, A1 => 
                           mult_21_C243_n86, SL => mult_21_C243_n823, Z => 
                           mult_21_C243_n1126);
   mult_21_C243_U623 : MUXB2DL port map( A0 => N3106, A1 => N3105, SL => 
                           mult_21_C243_n88, Z => mult_21_C243_n822);
   mult_21_C243_U622 : MUXB2DL port map( A0 => mult_21_C243_n84, A1 => 
                           mult_21_C243_n86, SL => mult_21_C243_n822, Z => 
                           mult_21_C243_n1125);
   mult_21_C243_U621 : MUXB2DL port map( A0 => N3107, A1 => mult_21_C243_n1545,
                           SL => mult_21_C243_n88, Z => mult_21_C243_n821);
   mult_21_C243_U620 : MUXB2DL port map( A0 => mult_21_C243_n84, A1 => 
                           mult_21_C243_n86, SL => mult_21_C243_n821, Z => 
                           mult_21_C243_n1124);
   mult_21_C243_U619 : MUXB2DL port map( A0 => N3108, A1 => N3107, SL => 
                           mult_21_C243_n88, Z => mult_21_C243_n820);
   mult_21_C243_U618 : MUXB2DL port map( A0 => mult_21_C243_n84, A1 => 
                           mult_21_C243_n86, SL => mult_21_C243_n820, Z => 
                           mult_21_C243_n1123);
   mult_21_C243_U617 : MUXB2DL port map( A0 => N3109, A1 => mult_21_C243_n1543,
                           SL => mult_21_C243_n88, Z => mult_21_C243_n819);
   mult_21_C243_U616 : MUXB2DL port map( A0 => mult_21_C243_n84, A1 => 
                           mult_21_C243_n86, SL => mult_21_C243_n819, Z => 
                           mult_21_C243_n1122);
   mult_21_C243_U615 : MUXB2DL port map( A0 => N3110, A1 => N3109, SL => 
                           mult_21_C243_n88, Z => mult_21_C243_n818);
   mult_21_C243_U614 : MUXB2DL port map( A0 => mult_21_C243_n84, A1 => 
                           mult_21_C243_n86, SL => mult_21_C243_n818, Z => 
                           mult_21_C243_n1121);
   mult_21_C243_U613 : MUXB2DL port map( A0 => N3111, A1 => N3110, SL => 
                           mult_21_C243_n88, Z => mult_21_C243_n817);
   mult_21_C243_U612 : MUXB2DL port map( A0 => mult_21_C243_n84, A1 => 
                           mult_21_C243_n86, SL => mult_21_C243_n817, Z => 
                           mult_21_C243_n1120);
   mult_21_C243_U611 : MUXB2DL port map( A0 => N3112, A1 => N3111, SL => 
                           mult_21_C243_n88, Z => mult_21_C243_n816);
   mult_21_C243_U610 : MUXB2DL port map( A0 => mult_21_C243_n84, A1 => 
                           mult_21_C243_n86, SL => mult_21_C243_n816, Z => 
                           mult_21_C243_n1119);
   mult_21_C243_U609 : MUXB2DL port map( A0 => N3113, A1 => N3112, SL => 
                           mult_21_C243_n88, Z => mult_21_C243_n815);
   mult_21_C243_U608 : MUXB2DL port map( A0 => mult_21_C243_n84, A1 => 
                           mult_21_C243_n86, SL => mult_21_C243_n815, Z => 
                           mult_21_C243_n1118);
   mult_21_C243_U607 : MUXB2DL port map( A0 => N3114, A1 => N3113, SL => 
                           mult_21_C243_n88, Z => mult_21_C243_n814);
   mult_21_C243_U606 : MUXB2DL port map( A0 => mult_21_C243_n84, A1 => 
                           mult_21_C243_n86, SL => mult_21_C243_n814, Z => 
                           mult_21_C243_n1117);
   mult_21_C243_U605 : NOR2M1D1 port map( A1 => mult_21_C243_n84, A2 => 
                           mult_21_C243_n86, Z => mult_21_C243_n1085);
   mult_21_C243_U604 : NAN2M1D1 port map( A1 => mult_21_C243_n93, A2 => N3105, 
                           Z => mult_21_C243_n813);
   mult_21_C243_U603 : MUXB2DL port map( A0 => mult_21_C243_n89, A1 => 
                           mult_21_C243_n91, SL => mult_21_C243_n813, Z => 
                           mult_21_C243_n1116);
   mult_21_C243_U602 : MUXB2DL port map( A0 => N3106, A1 => N3105, SL => 
                           mult_21_C243_n93, Z => mult_21_C243_n812);
   mult_21_C243_U601 : MUXB2DL port map( A0 => mult_21_C243_n89, A1 => 
                           mult_21_C243_n91, SL => mult_21_C243_n812, Z => 
                           mult_21_C243_n1115);
   mult_21_C243_U600 : MUXB2DL port map( A0 => N3107, A1 => mult_21_C243_n1545,
                           SL => mult_21_C243_n93, Z => mult_21_C243_n811);
   mult_21_C243_U599 : MUXB2DL port map( A0 => mult_21_C243_n89, A1 => 
                           mult_21_C243_n91, SL => mult_21_C243_n811, Z => 
                           mult_21_C243_n1114);
   mult_21_C243_U598 : MUXB2DL port map( A0 => N3108, A1 => N3107, SL => 
                           mult_21_C243_n93, Z => mult_21_C243_n810);
   mult_21_C243_U597 : MUXB2DL port map( A0 => mult_21_C243_n89, A1 => 
                           mult_21_C243_n91, SL => mult_21_C243_n810, Z => 
                           mult_21_C243_n1113);
   mult_21_C243_U596 : MUXB2DL port map( A0 => N3109, A1 => mult_21_C243_n1543,
                           SL => mult_21_C243_n93, Z => mult_21_C243_n809);
   mult_21_C243_U595 : MUXB2DL port map( A0 => mult_21_C243_n89, A1 => 
                           mult_21_C243_n91, SL => mult_21_C243_n809, Z => 
                           mult_21_C243_n1112);
   mult_21_C243_U594 : MUXB2DL port map( A0 => N3110, A1 => N3109, SL => 
                           mult_21_C243_n93, Z => mult_21_C243_n808);
   mult_21_C243_U593 : MUXB2DL port map( A0 => mult_21_C243_n89, A1 => 
                           mult_21_C243_n91, SL => mult_21_C243_n808, Z => 
                           mult_21_C243_n1111);
   mult_21_C243_U592 : MUXB2DL port map( A0 => N3111, A1 => N3110, SL => 
                           mult_21_C243_n93, Z => mult_21_C243_n807);
   mult_21_C243_U591 : MUXB2DL port map( A0 => mult_21_C243_n89, A1 => 
                           mult_21_C243_n91, SL => mult_21_C243_n807, Z => 
                           mult_21_C243_n1110);
   mult_21_C243_U590 : MUXB2DL port map( A0 => N3112, A1 => N3111, SL => 
                           mult_21_C243_n93, Z => mult_21_C243_n806);
   mult_21_C243_U589 : MUXB2DL port map( A0 => mult_21_C243_n89, A1 => 
                           mult_21_C243_n91, SL => mult_21_C243_n806, Z => 
                           mult_21_C243_n1109);
   mult_21_C243_U588 : NOR2M1D1 port map( A1 => mult_21_C243_n89, A2 => 
                           mult_21_C243_n91, Z => mult_21_C243_n1084);
   mult_21_C243_U587 : NAN2M1D1 port map( A1 => mult_21_C243_n98, A2 => N3105, 
                           Z => mult_21_C243_n805);
   mult_21_C243_U586 : MUXB2DL port map( A0 => mult_21_C243_n94, A1 => 
                           mult_21_C243_n96, SL => mult_21_C243_n805, Z => 
                           mult_21_C243_n1108);
   mult_21_C243_U585 : MUXB2DL port map( A0 => N3106, A1 => N3105, SL => 
                           mult_21_C243_n98, Z => mult_21_C243_n804);
   mult_21_C243_U584 : MUXB2DL port map( A0 => mult_21_C243_n94, A1 => 
                           mult_21_C243_n96, SL => mult_21_C243_n804, Z => 
                           mult_21_C243_n1107);
   mult_21_C243_U583 : MUXB2DL port map( A0 => N3107, A1 => mult_21_C243_n1545,
                           SL => mult_21_C243_n98, Z => mult_21_C243_n803);
   mult_21_C243_U582 : MUXB2DL port map( A0 => mult_21_C243_n94, A1 => 
                           mult_21_C243_n96, SL => mult_21_C243_n803, Z => 
                           mult_21_C243_n1106);
   mult_21_C243_U581 : MUXB2DL port map( A0 => N3108, A1 => N3107, SL => 
                           mult_21_C243_n98, Z => mult_21_C243_n802);
   mult_21_C243_U580 : MUXB2DL port map( A0 => mult_21_C243_n94, A1 => 
                           mult_21_C243_n96, SL => mult_21_C243_n802, Z => 
                           mult_21_C243_n1105);
   mult_21_C243_U579 : MUXB2DL port map( A0 => N3109, A1 => mult_21_C243_n1543,
                           SL => mult_21_C243_n98, Z => mult_21_C243_n801);
   mult_21_C243_U578 : MUXB2DL port map( A0 => mult_21_C243_n94, A1 => 
                           mult_21_C243_n96, SL => mult_21_C243_n801, Z => 
                           mult_21_C243_n1104);
   mult_21_C243_U577 : MUXB2DL port map( A0 => N3110, A1 => N3109, SL => 
                           mult_21_C243_n98, Z => mult_21_C243_n800);
   mult_21_C243_U576 : MUXB2DL port map( A0 => mult_21_C243_n94, A1 => 
                           mult_21_C243_n96, SL => mult_21_C243_n800, Z => 
                           mult_21_C243_n1103);
   mult_21_C243_U575 : NOR2M1D1 port map( A1 => mult_21_C243_n94, A2 => 
                           mult_21_C243_n96, Z => mult_21_C243_n1083);
   mult_21_C243_U574 : NAN2M1D1 port map( A1 => mult_21_C243_n103, A2 => N3105,
                           Z => mult_21_C243_n799);
   mult_21_C243_U573 : MUXB2DL port map( A0 => mult_21_C243_n99, A1 => 
                           mult_21_C243_n101, SL => mult_21_C243_n799, Z => 
                           mult_21_C243_n1102);
   mult_21_C243_U572 : MUXB2DL port map( A0 => N3106, A1 => N3105, SL => 
                           mult_21_C243_n103, Z => mult_21_C243_n798);
   mult_21_C243_U571 : MUXB2DL port map( A0 => mult_21_C243_n99, A1 => 
                           mult_21_C243_n101, SL => mult_21_C243_n798, Z => 
                           mult_21_C243_n1101);
   mult_21_C243_U570 : MUXB2DL port map( A0 => N3107, A1 => N3106, SL => 
                           mult_21_C243_n103, Z => mult_21_C243_n797);
   mult_21_C243_U569 : MUXB2DL port map( A0 => mult_21_C243_n99, A1 => 
                           mult_21_C243_n101, SL => mult_21_C243_n797, Z => 
                           mult_21_C243_n1100);
   mult_21_C243_U568 : MUXB2DL port map( A0 => N3108, A1 => N3107, SL => 
                           mult_21_C243_n103, Z => mult_21_C243_n796);
   mult_21_C243_U567 : MUXB2DL port map( A0 => mult_21_C243_n99, A1 => 
                           mult_21_C243_n101, SL => mult_21_C243_n796, Z => 
                           mult_21_C243_n1099);
   mult_21_C243_U566 : NOR2M1D1 port map( A1 => mult_21_C243_n99, A2 => 
                           mult_21_C243_n101, Z => mult_21_C243_n1082);
   mult_21_C243_U565 : NAN2M1D1 port map( A1 => mult_21_C243_n106, A2 => N3105,
                           Z => mult_21_C243_n795);
   mult_21_C243_U564 : MUXB2DL port map( A0 => mult_21_C243_n104, A1 => 
                           mult_21_C243_n105, SL => mult_21_C243_n795, Z => 
                           mult_21_C243_n1098);
   mult_21_C243_U563 : MUXB2DL port map( A0 => N3106, A1 => N3105, SL => 
                           mult_21_C243_n106, Z => mult_21_C243_n794);
   mult_21_C243_U562 : MUXB2DL port map( A0 => mult_21_C243_n104, A1 => 
                           mult_21_C243_n105, SL => mult_21_C243_n794, Z => 
                           mult_21_C243_n1097);
   mult_21_C243_U561 : NOR2M1D1 port map( A1 => mult_21_C243_n104, A2 => 
                           mult_21_C243_n105, Z => mult_21_C243_n1081);
   mult_21_C243_U557 : ADFULD1 port map( A => mult_21_C243_n1334, B => 
                           mult_21_C243_n1364, CI => mult_21_C243_n790, CO => 
                           mult_21_C243_n786, S => mult_21_C243_n787);
   mult_21_C243_U555 : ADFULD1 port map( A => mult_21_C243_n788, B => 
                           mult_21_C243_n1305, CI => mult_21_C243_n785, CO => 
                           mult_21_C243_n782, S => mult_21_C243_n783);
   mult_21_C243_U553 : ADFULD1 port map( A => mult_21_C243_n1304, B => 
                           mult_21_C243_n1362, CI => mult_21_C243_n1332, CO => 
                           mult_21_C243_n778, S => mult_21_C243_n779);
   mult_21_C243_U552 : ADFULD1 port map( A => mult_21_C243_n781, B => 
                           mult_21_C243_n784, CI => mult_21_C243_n779, CO => 
                           mult_21_C243_n776, S => mult_21_C243_n777);
   mult_21_C243_U550 : ADFULD1 port map( A => mult_21_C243_n1277, B => 
                           mult_21_C243_n1303, CI => mult_21_C243_n780, CO => 
                           mult_21_C243_n772, S => mult_21_C243_n773);
   mult_21_C243_U549 : ADFULD1 port map( A => mult_21_C243_n778, B => 
                           mult_21_C243_n775, CI => mult_21_C243_n773, CO => 
                           mult_21_C243_n770, S => mult_21_C243_n771);
   mult_21_C243_U547 : ADFULD1 port map( A => mult_21_C243_n1276, B => 
                           mult_21_C243_n1360, CI => mult_21_C243_n1330, CO => 
                           mult_21_C243_n766, S => mult_21_C243_n767);
   mult_21_C243_U546 : ADFULD1 port map( A => mult_21_C243_n774, B => 
                           mult_21_C243_n1302, CI => mult_21_C243_n769, CO => 
                           mult_21_C243_n764, S => mult_21_C243_n765);
   mult_21_C243_U545 : ADFULD1 port map( A => mult_21_C243_n767, B => 
                           mult_21_C243_n772, CI => mult_21_C243_n765, CO => 
                           mult_21_C243_n762, S => mult_21_C243_n763);
   mult_21_C243_U543 : ADFULD1 port map( A => mult_21_C243_n1275, B => 
                           mult_21_C243_n1251, CI => mult_21_C243_n1301, CO => 
                           mult_21_C243_n758, S => mult_21_C243_n759);
   mult_21_C243_U542 : ADFULD1 port map( A => mult_21_C243_n761, B => 
                           mult_21_C243_n768, CI => mult_21_C243_n766, CO => 
                           mult_21_C243_n756, S => mult_21_C243_n757);
   mult_21_C243_U541 : ADFULD1 port map( A => mult_21_C243_n764, B => 
                           mult_21_C243_n759, CI => mult_21_C243_n757, CO => 
                           mult_21_C243_n754, S => mult_21_C243_n755);
   mult_21_C243_U539 : ADFULD1 port map( A => mult_21_C243_n1250, B => 
                           mult_21_C243_n1358, CI => mult_21_C243_n1328, CO => 
                           mult_21_C243_n750, S => mult_21_C243_n751);
   mult_21_C243_U538 : ADFULD1 port map( A => mult_21_C243_n1274, B => 
                           mult_21_C243_n1300, CI => mult_21_C243_n760, CO => 
                           mult_21_C243_n748, S => mult_21_C243_n749);
   mult_21_C243_U537 : ADFULD1 port map( A => mult_21_C243_n758, B => 
                           mult_21_C243_n753, CI => mult_21_C243_n751, CO => 
                           mult_21_C243_n746, S => mult_21_C243_n747);
   mult_21_C243_U536 : ADFULD1 port map( A => mult_21_C243_n756, B => 
                           mult_21_C243_n749, CI => mult_21_C243_n747, CO => 
                           mult_21_C243_n744, S => mult_21_C243_n745);
   mult_21_C243_U534 : ADFULD1 port map( A => mult_21_C243_n1273, B => 
                           mult_21_C243_n1249, CI => mult_21_C243_n1227, CO => 
                           mult_21_C243_n740, S => mult_21_C243_n741);
   mult_21_C243_U533 : ADFULD1 port map( A => mult_21_C243_n752, B => 
                           mult_21_C243_n1299, CI => mult_21_C243_n743, CO => 
                           mult_21_C243_n738, S => mult_21_C243_n739);
   mult_21_C243_U532 : ADFULD1 port map( A => mult_21_C243_n748, B => 
                           mult_21_C243_n750, CI => mult_21_C243_n741, CO => 
                           mult_21_C243_n736, S => mult_21_C243_n737);
   mult_21_C243_U531 : ADFULD1 port map( A => mult_21_C243_n746, B => 
                           mult_21_C243_n739, CI => mult_21_C243_n737, CO => 
                           mult_21_C243_n734, S => mult_21_C243_n735);
   mult_21_C243_U529 : ADFULD1 port map( A => mult_21_C243_n1248, B => 
                           mult_21_C243_n1356, CI => mult_21_C243_n1326, CO => 
                           mult_21_C243_n730, S => mult_21_C243_n731);
   mult_21_C243_U528 : ADFULD1 port map( A => mult_21_C243_n1272, B => 
                           mult_21_C243_n1298, CI => mult_21_C243_n1226, CO => 
                           mult_21_C243_n728, S => mult_21_C243_n729);
   mult_21_C243_U527 : ADFULD1 port map( A => mult_21_C243_n733, B => 
                           mult_21_C243_n742, CI => mult_21_C243_n740, CO => 
                           mult_21_C243_n726, S => mult_21_C243_n727);
   mult_21_C243_U526 : ADFULD1 port map( A => mult_21_C243_n729, B => 
                           mult_21_C243_n731, CI => mult_21_C243_n738, CO => 
                           mult_21_C243_n724, S => mult_21_C243_n725);
   mult_21_C243_U525 : ADFULD1 port map( A => mult_21_C243_n736, B => 
                           mult_21_C243_n727, CI => mult_21_C243_n725, CO => 
                           mult_21_C243_n722, S => mult_21_C243_n723);
   mult_21_C243_U523 : ADFULD1 port map( A => mult_21_C243_n1271, B => 
                           mult_21_C243_n1297, CI => mult_21_C243_n1225, CO => 
                           mult_21_C243_n718, S => mult_21_C243_n719);
   mult_21_C243_U522 : ADFULD1 port map( A => mult_21_C243_n1205, B => 
                           mult_21_C243_n1247, CI => mult_21_C243_n732, CO => 
                           mult_21_C243_n716, S => mult_21_C243_n717);
   mult_21_C243_U521 : ADFULD1 port map( A => mult_21_C243_n730, B => 
                           mult_21_C243_n721, CI => mult_21_C243_n728, CO => 
                           mult_21_C243_n714, S => mult_21_C243_n715);
   mult_21_C243_U520 : ADFULD1 port map( A => mult_21_C243_n717, B => 
                           mult_21_C243_n719, CI => mult_21_C243_n726, CO => 
                           mult_21_C243_n712, S => mult_21_C243_n713);
   mult_21_C243_U519 : ADFULD1 port map( A => mult_21_C243_n724, B => 
                           mult_21_C243_n715, CI => mult_21_C243_n713, CO => 
                           mult_21_C243_n710, S => mult_21_C243_n711);
   mult_21_C243_U517 : ADFULD1 port map( A => mult_21_C243_n1204, B => 
                           mult_21_C243_n1354, CI => mult_21_C243_n1324, CO => 
                           mult_21_C243_n706, S => mult_21_C243_n707);
   mult_21_C243_U516 : ADFULD1 port map( A => mult_21_C243_n1246, B => 
                           mult_21_C243_n1296, CI => mult_21_C243_n1224, CO => 
                           mult_21_C243_n704, S => mult_21_C243_n705);
   mult_21_C243_U515 : ADFULD1 port map( A => mult_21_C243_n720, B => 
                           mult_21_C243_n1270, CI => mult_21_C243_n709, CO => 
                           mult_21_C243_n702, S => mult_21_C243_n703);
   mult_21_C243_U514 : ADFULD1 port map( A => mult_21_C243_n716, B => 
                           mult_21_C243_n718, CI => mult_21_C243_n707, CO => 
                           mult_21_C243_n700, S => mult_21_C243_n701);
   mult_21_C243_U513 : ADFULD1 port map( A => mult_21_C243_n703, B => 
                           mult_21_C243_n705, CI => mult_21_C243_n714, CO => 
                           mult_21_C243_n698, S => mult_21_C243_n699);
   mult_21_C243_U512 : ADFULD1 port map( A => mult_21_C243_n712, B => 
                           mult_21_C243_n701, CI => mult_21_C243_n699, CO => 
                           mult_21_C243_n696, S => mult_21_C243_n697);
   mult_21_C243_U510 : ADFULD1 port map( A => mult_21_C243_n1295, B => 
                           mult_21_C243_n1269, CI => mult_21_C243_n1223, CO => 
                           mult_21_C243_n692, S => mult_21_C243_n693);
   mult_21_C243_U509 : ADFULD1 port map( A => mult_21_C243_n1185, B => 
                           mult_21_C243_n1245, CI => mult_21_C243_n1203, CO => 
                           mult_21_C243_n690, S => mult_21_C243_n691);
   mult_21_C243_U508 : ADFULD1 port map( A => mult_21_C243_n695, B => 
                           mult_21_C243_n708, CI => mult_21_C243_n706, CO => 
                           mult_21_C243_n688, S => mult_21_C243_n689);
   mult_21_C243_U507 : ADFULD1 port map( A => mult_21_C243_n691, B => 
                           mult_21_C243_n704, CI => mult_21_C243_n693, CO => 
                           mult_21_C243_n686, S => mult_21_C243_n687);
   mult_21_C243_U506 : ADFULD1 port map( A => mult_21_C243_n700, B => 
                           mult_21_C243_n702, CI => mult_21_C243_n689, CO => 
                           mult_21_C243_n684, S => mult_21_C243_n685);
   mult_21_C243_U505 : ADFULD1 port map( A => mult_21_C243_n698, B => 
                           mult_21_C243_n687, CI => mult_21_C243_n685, CO => 
                           mult_21_C243_n682, S => mult_21_C243_n683);
   mult_21_C243_U503 : ADFULD1 port map( A => mult_21_C243_n1202, B => 
                           mult_21_C243_n1352, CI => mult_21_C243_n1322, CO => 
                           mult_21_C243_n678, S => mult_21_C243_n679);
   mult_21_C243_U502 : ADFULD1 port map( A => mult_21_C243_n1184, B => 
                           mult_21_C243_n1268, CI => mult_21_C243_n1222, CO => 
                           mult_21_C243_n676, S => mult_21_C243_n677);
   mult_21_C243_U501 : ADFULD1 port map( A => mult_21_C243_n1244, B => 
                           mult_21_C243_n1294, CI => mult_21_C243_n694, CO => 
                           mult_21_C243_n674, S => mult_21_C243_n675);
   mult_21_C243_U500 : ADFULD1 port map( A => mult_21_C243_n692, B => 
                           mult_21_C243_n681, CI => mult_21_C243_n690, CO => 
                           mult_21_C243_n672, S => mult_21_C243_n673);
   mult_21_C243_U499 : ADFULD1 port map( A => mult_21_C243_n677, B => 
                           mult_21_C243_n679, CI => mult_21_C243_n675, CO => 
                           mult_21_C243_n670, S => mult_21_C243_n671);
   mult_21_C243_U498 : ADFULD1 port map( A => mult_21_C243_n686, B => 
                           mult_21_C243_n688, CI => mult_21_C243_n673, CO => 
                           mult_21_C243_n668, S => mult_21_C243_n669);
   mult_21_C243_U497 : ADFULD1 port map( A => mult_21_C243_n684, B => 
                           mult_21_C243_n671, CI => mult_21_C243_n669, CO => 
                           mult_21_C243_n666, S => mult_21_C243_n667);
   mult_21_C243_U495 : ADFULD1 port map( A => mult_21_C243_n1293, B => 
                           mult_21_C243_n1201, CI => mult_21_C243_n1221, CO => 
                           mult_21_C243_n662, S => mult_21_C243_n663);
   mult_21_C243_U494 : ADFULD1 port map( A => mult_21_C243_n1183, B => 
                           mult_21_C243_n1167, CI => mult_21_C243_n1243, CO => 
                           mult_21_C243_n660, S => mult_21_C243_n661);
   mult_21_C243_U493 : ADFULD1 port map( A => mult_21_C243_n680, B => 
                           mult_21_C243_n1267, CI => mult_21_C243_n665, CO => 
                           mult_21_C243_n658, S => mult_21_C243_n659);
   mult_21_C243_U492 : ADFULD1 port map( A => mult_21_C243_n676, B => 
                           mult_21_C243_n678, CI => mult_21_C243_n674, CO => 
                           mult_21_C243_n656, S => mult_21_C243_n657);
   mult_21_C243_U491 : ADFULD1 port map( A => mult_21_C243_n663, B => 
                           mult_21_C243_n661, CI => mult_21_C243_n672, CO => 
                           mult_21_C243_n654, S => mult_21_C243_n655);
   mult_21_C243_U490 : ADFULD1 port map( A => mult_21_C243_n670, B => 
                           mult_21_C243_n659, CI => mult_21_C243_n657, CO => 
                           mult_21_C243_n652, S => mult_21_C243_n653);
   mult_21_C243_U489 : ADFULD1 port map( A => mult_21_C243_n668, B => 
                           mult_21_C243_n655, CI => mult_21_C243_n653, CO => 
                           mult_21_C243_n650, S => mult_21_C243_n651);
   mult_21_C243_U487 : ADFULD1 port map( A => mult_21_C243_n1200, B => 
                           mult_21_C243_n1350, CI => mult_21_C243_n1320, CO => 
                           mult_21_C243_n646, S => mult_21_C243_n647);
   mult_21_C243_U486 : ADFULD1 port map( A => mult_21_C243_n1166, B => 
                           mult_21_C243_n1266, CI => mult_21_C243_n1220, CO => 
                           mult_21_C243_n644, S => mult_21_C243_n645);
   mult_21_C243_U485 : ADFULD1 port map( A => mult_21_C243_n1182, B => 
                           mult_21_C243_n1292, CI => mult_21_C243_n1242, CO => 
                           mult_21_C243_n642, S => mult_21_C243_n643);
   mult_21_C243_U484 : ADFULD1 port map( A => mult_21_C243_n649, B => 
                           mult_21_C243_n664, CI => mult_21_C243_n662, CO => 
                           mult_21_C243_n640, S => mult_21_C243_n641);
   mult_21_C243_U483 : ADFULD1 port map( A => mult_21_C243_n647, B => 
                           mult_21_C243_n660, CI => mult_21_C243_n643, CO => 
                           mult_21_C243_n638, S => mult_21_C243_n639);
   mult_21_C243_U482 : ADFULD1 port map( A => mult_21_C243_n658, B => 
                           mult_21_C243_n645, CI => mult_21_C243_n656, CO => 
                           mult_21_C243_n636, S => mult_21_C243_n637);
   mult_21_C243_U481 : ADFULD1 port map( A => mult_21_C243_n639, B => 
                           mult_21_C243_n641, CI => mult_21_C243_n654, CO => 
                           mult_21_C243_n634, S => mult_21_C243_n635);
   mult_21_C243_U480 : ADFULD1 port map( A => mult_21_C243_n652, B => 
                           mult_21_C243_n637, CI => mult_21_C243_n635, CO => 
                           mult_21_C243_n632, S => mult_21_C243_n633);
   mult_21_C243_U478 : ADFULD1 port map( A => mult_21_C243_n1151, B => 
                           mult_21_C243_n1199, CI => mult_21_C243_n1219, CO => 
                           mult_21_C243_n628, S => mult_21_C243_n629);
   mult_21_C243_U477 : ADFULD1 port map( A => mult_21_C243_n1291, B => 
                           mult_21_C243_n1181, CI => mult_21_C243_n1165, CO => 
                           mult_21_C243_n626, S => mult_21_C243_n627);
   mult_21_C243_U476 : ADFULD1 port map( A => mult_21_C243_n1241, B => 
                           mult_21_C243_n1265, CI => mult_21_C243_n648, CO => 
                           mult_21_C243_n624, S => mult_21_C243_n625);
   mult_21_C243_U475 : ADFULD1 port map( A => mult_21_C243_n646, B => 
                           mult_21_C243_n631, CI => mult_21_C243_n642, CO => 
                           mult_21_C243_n622, S => mult_21_C243_n623);
   mult_21_C243_U474 : ADFULD1 port map( A => mult_21_C243_n627, B => 
                           mult_21_C243_n644, CI => mult_21_C243_n629, CO => 
                           mult_21_C243_n620, S => mult_21_C243_n621);
   mult_21_C243_U473 : ADFULD1 port map( A => mult_21_C243_n640, B => 
                           mult_21_C243_n625, CI => mult_21_C243_n638, CO => 
                           mult_21_C243_n618, S => mult_21_C243_n619);
   mult_21_C243_U472 : ADFULD1 port map( A => mult_21_C243_n621, B => 
                           mult_21_C243_n623, CI => mult_21_C243_n636, CO => 
                           mult_21_C243_n616, S => mult_21_C243_n617);
   mult_21_C243_U471 : ADFULD1 port map( A => mult_21_C243_n634, B => 
                           mult_21_C243_n619, CI => mult_21_C243_n617, CO => 
                           mult_21_C243_n614, S => mult_21_C243_n615);
   mult_21_C243_U469 : ADFULD1 port map( A => mult_21_C243_n1164, B => 
                           mult_21_C243_n1348, CI => mult_21_C243_n1318, CO => 
                           mult_21_C243_n610, S => mult_21_C243_n611);
   mult_21_C243_U468 : ADFULD1 port map( A => mult_21_C243_n1290, B => 
                           mult_21_C243_n1198, CI => mult_21_C243_n1218, CO => 
                           mult_21_C243_n608, S => mult_21_C243_n609);
   mult_21_C243_U467 : ADFULD1 port map( A => mult_21_C243_n1150, B => 
                           mult_21_C243_n1264, CI => mult_21_C243_n1180, CO => 
                           mult_21_C243_n606, S => mult_21_C243_n607);
   mult_21_C243_U466 : ADFULD1 port map( A => mult_21_C243_n630, B => 
                           mult_21_C243_n1240, CI => mult_21_C243_n613, CO => 
                           mult_21_C243_n604, S => mult_21_C243_n605);
   mult_21_C243_U465 : ADFULD1 port map( A => mult_21_C243_n626, B => 
                           mult_21_C243_n628, CI => mult_21_C243_n624, CO => 
                           mult_21_C243_n602, S => mult_21_C243_n603);
   mult_21_C243_U464 : ADFULD1 port map( A => mult_21_C243_n609, B => 
                           mult_21_C243_n611, CI => mult_21_C243_n607, CO => 
                           mult_21_C243_n600, S => mult_21_C243_n601);
   mult_21_C243_U463 : ADFULD1 port map( A => mult_21_C243_n622, B => 
                           mult_21_C243_n605, CI => mult_21_C243_n620, CO => 
                           mult_21_C243_n598, S => mult_21_C243_n599);
   mult_21_C243_U462 : ADFULD1 port map( A => mult_21_C243_n601, B => 
                           mult_21_C243_n603, CI => mult_21_C243_n618, CO => 
                           mult_21_C243_n596, S => mult_21_C243_n597);
   mult_21_C243_U461 : ADFULD1 port map( A => mult_21_C243_n616, B => 
                           mult_21_C243_n599, CI => mult_21_C243_n597, CO => 
                           mult_21_C243_n594, S => mult_21_C243_n595);
   mult_21_C243_U459 : ADFULD1 port map( A => mult_21_C243_n1289, B => 
                           mult_21_C243_n1179, CI => mult_21_C243_n1217, CO => 
                           mult_21_C243_n590, S => mult_21_C243_n591);
   mult_21_C243_U458 : ADFULD1 port map( A => mult_21_C243_n1263, B => 
                           mult_21_C243_n1149, CI => mult_21_C243_n1137, CO => 
                           mult_21_C243_n588, S => mult_21_C243_n589);
   mult_21_C243_U457 : ADFULD1 port map( A => mult_21_C243_n1163, B => 
                           mult_21_C243_n1239, CI => mult_21_C243_n1197, CO => 
                           mult_21_C243_n586, S => mult_21_C243_n587);
   mult_21_C243_U456 : ADFULD1 port map( A => mult_21_C243_n593, B => 
                           mult_21_C243_n612, CI => mult_21_C243_n610, CO => 
                           mult_21_C243_n584, S => mult_21_C243_n585);
   mult_21_C243_U455 : ADFULD1 port map( A => mult_21_C243_n606, B => 
                           mult_21_C243_n608, CI => mult_21_C243_n587, CO => 
                           mult_21_C243_n582, S => mult_21_C243_n583);
   mult_21_C243_U454 : ADFULD1 port map( A => mult_21_C243_n591, B => 
                           mult_21_C243_n589, CI => mult_21_C243_n604, CO => 
                           mult_21_C243_n580, S => mult_21_C243_n581);
   mult_21_C243_U453 : ADFULD1 port map( A => mult_21_C243_n585, B => 
                           mult_21_C243_n602, CI => mult_21_C243_n600, CO => 
                           mult_21_C243_n578, S => mult_21_C243_n579);
   mult_21_C243_U452 : ADFULD1 port map( A => mult_21_C243_n581, B => 
                           mult_21_C243_n583, CI => mult_21_C243_n598, CO => 
                           mult_21_C243_n576, S => mult_21_C243_n577);
   mult_21_C243_U451 : ADFULD1 port map( A => mult_21_C243_n596, B => 
                           mult_21_C243_n579, CI => mult_21_C243_n577, CO => 
                           mult_21_C243_n574, S => mult_21_C243_n575);
   mult_21_C243_U449 : ADFULD1 port map( A => mult_21_C243_n1136, B => 
                           mult_21_C243_n1346, CI => mult_21_C243_n1316, CO => 
                           mult_21_C243_n570, S => mult_21_C243_n571);
   mult_21_C243_U448 : ADFULD1 port map( A => mult_21_C243_n1288, B => 
                           mult_21_C243_n1178, CI => mult_21_C243_n1216, CO => 
                           mult_21_C243_n568, S => mult_21_C243_n569);
   mult_21_C243_U447 : ADFULD1 port map( A => mult_21_C243_n1148, B => 
                           mult_21_C243_n1262, CI => mult_21_C243_n1162, CO => 
                           mult_21_C243_n566, S => mult_21_C243_n567);
   mult_21_C243_U446 : ADFULD1 port map( A => mult_21_C243_n1196, B => 
                           mult_21_C243_n1238, CI => mult_21_C243_n592, CO => 
                           mult_21_C243_n564, S => mult_21_C243_n565);
   mult_21_C243_U445 : ADFULD1 port map( A => mult_21_C243_n590, B => 
                           mult_21_C243_n573, CI => mult_21_C243_n588, CO => 
                           mult_21_C243_n562, S => mult_21_C243_n563);
   mult_21_C243_U444 : ADFULD1 port map( A => mult_21_C243_n571, B => 
                           mult_21_C243_n586, CI => mult_21_C243_n567, CO => 
                           mult_21_C243_n560, S => mult_21_C243_n561);
   mult_21_C243_U443 : ADFULD1 port map( A => mult_21_C243_n565, B => 
                           mult_21_C243_n569, CI => mult_21_C243_n584, CO => 
                           mult_21_C243_n558, S => mult_21_C243_n559);
   mult_21_C243_U442 : ADFULD1 port map( A => mult_21_C243_n563, B => 
                           mult_21_C243_n582, CI => mult_21_C243_n580, CO => 
                           mult_21_C243_n556, S => mult_21_C243_n557);
   mult_21_C243_U441 : ADFULD1 port map( A => mult_21_C243_n559, B => 
                           mult_21_C243_n561, CI => mult_21_C243_n578, CO => 
                           mult_21_C243_n554, S => mult_21_C243_n555);
   mult_21_C243_U440 : ADFULD1 port map( A => mult_21_C243_n576, B => 
                           mult_21_C243_n557, CI => mult_21_C243_n555, CO => 
                           mult_21_C243_n552, S => mult_21_C243_n553);
   mult_21_C243_U438 : ADFULD1 port map( A => mult_21_C243_n1125, B => 
                           mult_21_C243_n1177, CI => mult_21_C243_n1215, CO => 
                           mult_21_C243_n548, S => mult_21_C243_n549);
   mult_21_C243_U437 : ADFULD1 port map( A => mult_21_C243_n1287, B => 
                           mult_21_C243_n1161, CI => mult_21_C243_n1261, CO => 
                           mult_21_C243_n546, S => mult_21_C243_n547);
   mult_21_C243_U436 : ADFULD1 port map( A => mult_21_C243_n1135, B => 
                           mult_21_C243_n1237, CI => mult_21_C243_n1147, CO => 
                           mult_21_C243_n544, S => mult_21_C243_n545);
   mult_21_C243_U435 : ADFULD1 port map( A => mult_21_C243_n572, B => 
                           mult_21_C243_n1195, CI => mult_21_C243_n551, CO => 
                           mult_21_C243_n542, S => mult_21_C243_n543);
   mult_21_C243_U434 : ADFULD1 port map( A => mult_21_C243_n566, B => 
                           mult_21_C243_n570, CI => mult_21_C243_n568, CO => 
                           mult_21_C243_n540, S => mult_21_C243_n541);
   mult_21_C243_U433 : ADFULD1 port map( A => mult_21_C243_n549, B => 
                           mult_21_C243_n564, CI => mult_21_C243_n547, CO => 
                           mult_21_C243_n538, S => mult_21_C243_n539);
   mult_21_C243_U432 : ADFULD1 port map( A => mult_21_C243_n562, B => 
                           mult_21_C243_n545, CI => mult_21_C243_n543, CO => 
                           mult_21_C243_n536, S => mult_21_C243_n537);
   mult_21_C243_U431 : ADFULD1 port map( A => mult_21_C243_n541, B => 
                           mult_21_C243_n560, CI => mult_21_C243_n558, CO => 
                           mult_21_C243_n534, S => mult_21_C243_n535);
   mult_21_C243_U430 : ADFULD1 port map( A => mult_21_C243_n556, B => 
                           mult_21_C243_n539, CI => mult_21_C243_n537, CO => 
                           mult_21_C243_n532, S => mult_21_C243_n533);
   mult_21_C243_U429 : ADFULD1 port map( A => mult_21_C243_n554, B => 
                           mult_21_C243_n535, CI => mult_21_C243_n533, CO => 
                           mult_21_C243_n530, S => mult_21_C243_n531);
   mult_21_C243_U427 : ADFULD1 port map( A => mult_21_C243_n1146, B => 
                           mult_21_C243_n1344, CI => mult_21_C243_n1314, CO => 
                           mult_21_C243_n526, S => mult_21_C243_n527);
   mult_21_C243_U426 : ADFULD1 port map( A => mult_21_C243_n1124, B => 
                           mult_21_C243_n1176, CI => mult_21_C243_n1214, CO => 
                           mult_21_C243_n524, S => mult_21_C243_n525);
   mult_21_C243_U425 : ADFULD1 port map( A => mult_21_C243_n1134, B => 
                           mult_21_C243_n1286, CI => mult_21_C243_n1160, CO => 
                           mult_21_C243_n522, S => mult_21_C243_n523);
   mult_21_C243_U424 : ADFULD1 port map( A => mult_21_C243_n1194, B => 
                           mult_21_C243_n1260, CI => mult_21_C243_n1236, CO => 
                           mult_21_C243_n520, S => mult_21_C243_n521);
   mult_21_C243_U423 : ADFULD1 port map( A => mult_21_C243_n529, B => 
                           mult_21_C243_n550, CI => mult_21_C243_n548, CO => 
                           mult_21_C243_n518, S => mult_21_C243_n519);
   mult_21_C243_U422 : ADFULD1 port map( A => mult_21_C243_n544, B => 
                           mult_21_C243_n546, CI => mult_21_C243_n527, CO => 
                           mult_21_C243_n516, S => mult_21_C243_n517);
   mult_21_C243_U421 : ADFULD1 port map( A => mult_21_C243_n525, B => 
                           mult_21_C243_n521, CI => mult_21_C243_n523, CO => 
                           mult_21_C243_n514, S => mult_21_C243_n515);
   mult_21_C243_U420 : ADFULD1 port map( A => mult_21_C243_n540, B => 
                           mult_21_C243_n542, CI => mult_21_C243_n519, CO => 
                           mult_21_C243_n512, S => mult_21_C243_n513);
   mult_21_C243_U419 : ADFULD1 port map( A => mult_21_C243_n517, B => 
                           mult_21_C243_n538, CI => mult_21_C243_n515, CO => 
                           mult_21_C243_n510, S => mult_21_C243_n511);
   mult_21_C243_U418 : ADFULD1 port map( A => mult_21_C243_n513, B => 
                           mult_21_C243_n536, CI => mult_21_C243_n534, CO => 
                           mult_21_C243_n508, S => mult_21_C243_n509);
   mult_21_C243_U417 : ADFULD1 port map( A => mult_21_C243_n532, B => 
                           mult_21_C243_n511, CI => mult_21_C243_n509, CO => 
                           mult_21_C243_n506, S => mult_21_C243_n507);
   mult_21_C243_U415 : ADFULD1 port map( A => mult_21_C243_n1115, B => 
                           mult_21_C243_n1175, CI => mult_21_C243_n1213, CO => 
                           mult_21_C243_n502, S => mult_21_C243_n503);
   mult_21_C243_U414 : ADFULD1 port map( A => mult_21_C243_n1123, B => 
                           mult_21_C243_n1145, CI => mult_21_C243_n1133, CO => 
                           mult_21_C243_n500, S => mult_21_C243_n501);
   mult_21_C243_U413 : ADFULD1 port map( A => mult_21_C243_n1159, B => 
                           mult_21_C243_n1285, CI => mult_21_C243_n1193, CO => 
                           mult_21_C243_n498, S => mult_21_C243_n499);
   mult_21_C243_U412 : ADFULD1 port map( A => mult_21_C243_n1235, B => 
                           mult_21_C243_n1259, CI => mult_21_C243_n528, CO => 
                           mult_21_C243_n496, S => mult_21_C243_n497);
   mult_21_C243_U411 : ADFULD1 port map( A => mult_21_C243_n526, B => 
                           mult_21_C243_n505, CI => mult_21_C243_n520, CO => 
                           mult_21_C243_n494, S => mult_21_C243_n495);
   mult_21_C243_U410 : ADFULD1 port map( A => mult_21_C243_n522, B => 
                           mult_21_C243_n524, CI => mult_21_C243_n499, CO => 
                           mult_21_C243_n492, S => mult_21_C243_n493);
   mult_21_C243_U409 : ADFULD1 port map( A => mult_21_C243_n501, B => 
                           mult_21_C243_n503, CI => mult_21_C243_n497, CO => 
                           mult_21_C243_n490, S => mult_21_C243_n491);
   mult_21_C243_U408 : ADFULD1 port map( A => mult_21_C243_n516, B => 
                           mult_21_C243_n518, CI => mult_21_C243_n495, CO => 
                           mult_21_C243_n488, S => mult_21_C243_n489);
   mult_21_C243_U407 : ADFULD1 port map( A => mult_21_C243_n493, B => 
                           mult_21_C243_n514, CI => mult_21_C243_n491, CO => 
                           mult_21_C243_n486, S => mult_21_C243_n487);
   mult_21_C243_U406 : ADFULD1 port map( A => mult_21_C243_n510, B => 
                           mult_21_C243_n512, CI => mult_21_C243_n489, CO => 
                           mult_21_C243_n484, S => mult_21_C243_n485);
   mult_21_C243_U405 : ADFULD1 port map( A => mult_21_C243_n508, B => 
                           mult_21_C243_n487, CI => mult_21_C243_n485, CO => 
                           mult_21_C243_n482, S => mult_21_C243_n483);
   mult_21_C243_U403 : ADFULD1 port map( A => mult_21_C243_n1114, B => 
                           mult_21_C243_n1342, CI => mult_21_C243_n1312, CO => 
                           mult_21_C243_n478, S => mult_21_C243_n479);
   mult_21_C243_U402 : ADFULD1 port map( A => mult_21_C243_n1284, B => 
                           mult_21_C243_n1174, CI => mult_21_C243_n1212, CO => 
                           mult_21_C243_n476, S => mult_21_C243_n477);
   mult_21_C243_U401 : ADFULD1 port map( A => mult_21_C243_n1258, B => 
                           mult_21_C243_n1132, CI => mult_21_C243_n1122, CO => 
                           mult_21_C243_n474, S => mult_21_C243_n475);
   mult_21_C243_U400 : ADFULD1 port map( A => mult_21_C243_n1144, B => 
                           mult_21_C243_n1234, CI => mult_21_C243_n1158, CO => 
                           mult_21_C243_n472, S => mult_21_C243_n473);
   mult_21_C243_U399 : ADFULD1 port map( A => mult_21_C243_n504, B => 
                           mult_21_C243_n1192, CI => mult_21_C243_n481, CO => 
                           mult_21_C243_n470, S => mult_21_C243_n471);
   mult_21_C243_U398 : ADFULD1 port map( A => mult_21_C243_n498, B => 
                           mult_21_C243_n502, CI => mult_21_C243_n496, CO => 
                           mult_21_C243_n468, S => mult_21_C243_n469);
   mult_21_C243_U397 : ADFULD1 port map( A => mult_21_C243_n479, B => 
                           mult_21_C243_n500, CI => mult_21_C243_n473, CO => 
                           mult_21_C243_n466, S => mult_21_C243_n467);
   mult_21_C243_U396 : ADFULD1 port map( A => mult_21_C243_n475, B => 
                           mult_21_C243_n477, CI => mult_21_C243_n471, CO => 
                           mult_21_C243_n464, S => mult_21_C243_n465);
   mult_21_C243_U395 : ADFULD1 port map( A => mult_21_C243_n492, B => 
                           mult_21_C243_n494, CI => mult_21_C243_n490, CO => 
                           mult_21_C243_n462, S => mult_21_C243_n463);
   mult_21_C243_U394 : ADFULD1 port map( A => mult_21_C243_n467, B => 
                           mult_21_C243_n469, CI => mult_21_C243_n465, CO => 
                           mult_21_C243_n460, S => mult_21_C243_n461);
   mult_21_C243_U393 : ADFULD1 port map( A => mult_21_C243_n486, B => 
                           mult_21_C243_n488, CI => mult_21_C243_n463, CO => 
                           mult_21_C243_n458, S => mult_21_C243_n459);
   mult_21_C243_U392 : ADFULD1 port map( A => mult_21_C243_n484, B => 
                           mult_21_C243_n461, CI => mult_21_C243_n459, CO => 
                           mult_21_C243_n456, S => mult_21_C243_n457);
   mult_21_C243_U390 : ADFULD1 port map( A => mult_21_C243_n1107, B => 
                           mult_21_C243_n1157, CI => mult_21_C243_n1211, CO => 
                           mult_21_C243_n452, S => mult_21_C243_n453);
   mult_21_C243_U389 : ADFULD1 port map( A => mult_21_C243_n1283, B => 
                           mult_21_C243_n1143, CI => mult_21_C243_n1257, CO => 
                           mult_21_C243_n450, S => mult_21_C243_n451);
   mult_21_C243_U388 : ADFULD1 port map( A => mult_21_C243_n1113, B => 
                           mult_21_C243_n1233, CI => mult_21_C243_n1121, CO => 
                           mult_21_C243_n448, S => mult_21_C243_n449);
   mult_21_C243_U387 : ADFULD1 port map( A => mult_21_C243_n1131, B => 
                           mult_21_C243_n1191, CI => mult_21_C243_n1173, CO => 
                           mult_21_C243_n446, S => mult_21_C243_n447);
   mult_21_C243_U386 : ADFULD1 port map( A => mult_21_C243_n455, B => 
                           mult_21_C243_n480, CI => mult_21_C243_n478, CO => 
                           mult_21_C243_n444, S => mult_21_C243_n445);
   mult_21_C243_U385 : ADFULD1 port map( A => mult_21_C243_n474, B => 
                           mult_21_C243_n472, CI => mult_21_C243_n476, CO => 
                           mult_21_C243_n442, S => mult_21_C243_n443);
   mult_21_C243_U384 : ADFULD1 port map( A => mult_21_C243_n453, B => 
                           mult_21_C243_n447, CI => mult_21_C243_n470, CO => 
                           mult_21_C243_n440, S => mult_21_C243_n441);
   mult_21_C243_U383 : ADFULD1 port map( A => mult_21_C243_n449, B => 
                           mult_21_C243_n451, CI => mult_21_C243_n468, CO => 
                           mult_21_C243_n438, S => mult_21_C243_n439);
   mult_21_C243_U382 : ADFULD1 port map( A => mult_21_C243_n466, B => 
                           mult_21_C243_n445, CI => mult_21_C243_n443, CO => 
                           mult_21_C243_n436, S => mult_21_C243_n437);
   mult_21_C243_U381 : ADFULD1 port map( A => mult_21_C243_n441, B => 
                           mult_21_C243_n464, CI => mult_21_C243_n462, CO => 
                           mult_21_C243_n434, S => mult_21_C243_n435);
   mult_21_C243_U380 : ADFULD1 port map( A => mult_21_C243_n437, B => 
                           mult_21_C243_n439, CI => mult_21_C243_n460, CO => 
                           mult_21_C243_n432, S => mult_21_C243_n433);
   mult_21_C243_U379 : ADFULD1 port map( A => mult_21_C243_n458, B => 
                           mult_21_C243_n435, CI => mult_21_C243_n433, CO => 
                           mult_21_C243_n430, S => mult_21_C243_n431);
   mult_21_C243_U377 : ADFULD1 port map( A => mult_21_C243_n1106, B => 
                           mult_21_C243_n1340, CI => mult_21_C243_n1310, CO => 
                           mult_21_C243_n426, S => mult_21_C243_n427);
   mult_21_C243_U376 : ADFULD1 port map( A => mult_21_C243_n1282, B => 
                           mult_21_C243_n1156, CI => mult_21_C243_n1210, CO => 
                           mult_21_C243_n424, S => mult_21_C243_n425);
   mult_21_C243_U375 : ADFULD1 port map( A => mult_21_C243_n1112, B => 
                           mult_21_C243_n1130, CI => mult_21_C243_n1120, CO => 
                           mult_21_C243_n422, S => mult_21_C243_n423);
   mult_21_C243_U374 : ADFULD1 port map( A => mult_21_C243_n1142, B => 
                           mult_21_C243_n1256, CI => mult_21_C243_n1172, CO => 
                           mult_21_C243_n420, S => mult_21_C243_n421);
   mult_21_C243_U373 : ADFULD1 port map( A => mult_21_C243_n1232, B => 
                           mult_21_C243_n1190, CI => mult_21_C243_n454, CO => 
                           mult_21_C243_n418, S => mult_21_C243_n419);
   mult_21_C243_U372 : ADFULD1 port map( A => mult_21_C243_n452, B => 
                           mult_21_C243_n429, CI => mult_21_C243_n450, CO => 
                           mult_21_C243_n416, S => mult_21_C243_n417);
   mult_21_C243_U371 : ADFULD1 port map( A => mult_21_C243_n448, B => 
                           mult_21_C243_n446, CI => mult_21_C243_n427, CO => 
                           mult_21_C243_n414, S => mult_21_C243_n415);
   mult_21_C243_U370 : ADFULD1 port map( A => mult_21_C243_n421, B => 
                           mult_21_C243_n423, CI => mult_21_C243_n425, CO => 
                           mult_21_C243_n412, S => mult_21_C243_n413);
   mult_21_C243_U369 : ADFULD1 port map( A => mult_21_C243_n444, B => 
                           mult_21_C243_n419, CI => mult_21_C243_n442, CO => 
                           mult_21_C243_n410, S => mult_21_C243_n411);
   mult_21_C243_U368 : ADFULD1 port map( A => mult_21_C243_n440, B => 
                           mult_21_C243_n417, CI => mult_21_C243_n415, CO => 
                           mult_21_C243_n408, S => mult_21_C243_n409);
   mult_21_C243_U367 : ADFULD1 port map( A => mult_21_C243_n438, B => 
                           mult_21_C243_n413, CI => mult_21_C243_n411, CO => 
                           mult_21_C243_n406, S => mult_21_C243_n407);
   mult_21_C243_U366 : ADFULD1 port map( A => mult_21_C243_n409, B => 
                           mult_21_C243_n436, CI => mult_21_C243_n434, CO => 
                           mult_21_C243_n404, S => mult_21_C243_n405);
   mult_21_C243_U365 : ADFULD1 port map( A => mult_21_C243_n432, B => 
                           mult_21_C243_n407, CI => mult_21_C243_n405, CO => 
                           mult_21_C243_n402, S => mult_21_C243_n403);
   mult_21_C243_U363 : ADFULD1 port map( A => mult_21_C243_n1281, B => 
                           mult_21_C243_n1155, CI => mult_21_C243_n1209, CO => 
                           mult_21_C243_n398, S => mult_21_C243_n399);
   mult_21_C243_U362 : ADFULD1 port map( A => mult_21_C243_n1255, B => 
                           mult_21_C243_n1119, CI => mult_21_C243_n1101, CO => 
                           mult_21_C243_n396, S => mult_21_C243_n397);
   mult_21_C243_U361 : ADFULD1 port map( A => mult_21_C243_n1231, B => 
                           mult_21_C243_n1111, CI => mult_21_C243_n1105, CO => 
                           mult_21_C243_n394, S => mult_21_C243_n395);
   mult_21_C243_U360 : ADFULD1 port map( A => mult_21_C243_n1129, B => 
                           mult_21_C243_n1189, CI => mult_21_C243_n1141, CO => 
                           mult_21_C243_n392, S => mult_21_C243_n393);
   mult_21_C243_U359 : ADFULD1 port map( A => mult_21_C243_n428, B => 
                           mult_21_C243_n1171, CI => mult_21_C243_n401, CO => 
                           mult_21_C243_n390, S => mult_21_C243_n391);
   mult_21_C243_U358 : ADFULD1 port map( A => mult_21_C243_n424, B => 
                           mult_21_C243_n426, CI => mult_21_C243_n420, CO => 
                           mult_21_C243_n388, S => mult_21_C243_n389);
   mult_21_C243_U357 : ADFULD1 port map( A => mult_21_C243_n418, B => 
                           mult_21_C243_n422, CI => mult_21_C243_n393, CO => 
                           mult_21_C243_n386, S => mult_21_C243_n387);
   mult_21_C243_U356 : ADFULD1 port map( A => mult_21_C243_n395, B => 
                           mult_21_C243_n397, CI => mult_21_C243_n399, CO => 
                           mult_21_C243_n384, S => mult_21_C243_n385);
   mult_21_C243_U355 : ADFULD1 port map( A => mult_21_C243_n391, B => 
                           mult_21_C243_n416, CI => mult_21_C243_n414, CO => 
                           mult_21_C243_n382, S => mult_21_C243_n383);
   mult_21_C243_U354 : ADFULD1 port map( A => mult_21_C243_n412, B => 
                           mult_21_C243_n389, CI => mult_21_C243_n387, CO => 
                           mult_21_C243_n380, S => mult_21_C243_n381);
   mult_21_C243_U353 : ADFULD1 port map( A => mult_21_C243_n410, B => 
                           mult_21_C243_n385, CI => mult_21_C243_n383, CO => 
                           mult_21_C243_n378, S => mult_21_C243_n379);
   mult_21_C243_U352 : ADFULD1 port map( A => mult_21_C243_n381, B => 
                           mult_21_C243_n408, CI => mult_21_C243_n406, CO => 
                           mult_21_C243_n376, S => mult_21_C243_n377);
   mult_21_C243_U351 : ADFULD1 port map( A => mult_21_C243_n404, B => 
                           mult_21_C243_n379, CI => mult_21_C243_n377, CO => 
                           mult_21_C243_n374, S => mult_21_C243_n375);
   mult_21_C243_U349 : ADFULD1 port map( A => mult_21_C243_n1100, B => 
                           mult_21_C243_n1338, CI => mult_21_C243_n1308, CO => 
                           mult_21_C243_n370, S => mult_21_C243_n371);
   mult_21_C243_U348 : ADFULD1 port map( A => mult_21_C243_n1280, B => 
                           mult_21_C243_n1154, CI => mult_21_C243_n1208, CO => 
                           mult_21_C243_n368, S => mult_21_C243_n369);
   mult_21_C243_U347 : ADFULD1 port map( A => mult_21_C243_n1254, B => 
                           mult_21_C243_n1128, CI => mult_21_C243_n1230, CO => 
                           mult_21_C243_n366, S => mult_21_C243_n367);
   mult_21_C243_U346 : ADFULD1 port map( A => mult_21_C243_n1104, B => 
                           mult_21_C243_n1188, CI => mult_21_C243_n1110, CO => 
                           mult_21_C243_n364, S => mult_21_C243_n365);
   mult_21_C243_U345 : ADFULD1 port map( A => mult_21_C243_n1170, B => 
                           mult_21_C243_n1118, CI => mult_21_C243_n1140, CO => 
                           mult_21_C243_n362, S => mult_21_C243_n363);
   mult_21_C243_U344 : ADFULD1 port map( A => mult_21_C243_n373, B => 
                           mult_21_C243_n400, CI => mult_21_C243_n392, CO => 
                           mult_21_C243_n360, S => mult_21_C243_n361);
   mult_21_C243_U343 : ADFULD1 port map( A => mult_21_C243_n398, B => 
                           mult_21_C243_n394, CI => mult_21_C243_n396, CO => 
                           mult_21_C243_n358, S => mult_21_C243_n359);
   mult_21_C243_U342 : ADFULD1 port map( A => mult_21_C243_n369, B => 
                           mult_21_C243_n371, CI => mult_21_C243_n367, CO => 
                           mult_21_C243_n356, S => mult_21_C243_n357);
   mult_21_C243_U341 : ADFULD1 port map( A => mult_21_C243_n365, B => 
                           mult_21_C243_n363, CI => mult_21_C243_n390, CO => 
                           mult_21_C243_n354, S => mult_21_C243_n355);
   mult_21_C243_U340 : ADFULD1 port map( A => mult_21_C243_n361, B => 
                           mult_21_C243_n388, CI => mult_21_C243_n386, CO => 
                           mult_21_C243_n352, S => mult_21_C243_n353);
   mult_21_C243_U339 : ADFULD1 port map( A => mult_21_C243_n359, B => 
                           mult_21_C243_n384, CI => mult_21_C243_n357, CO => 
                           mult_21_C243_n350, S => mult_21_C243_n351);
   mult_21_C243_U338 : ADFULD1 port map( A => mult_21_C243_n382, B => 
                           mult_21_C243_n355, CI => mult_21_C243_n380, CO => 
                           mult_21_C243_n348, S => mult_21_C243_n349);
   mult_21_C243_U337 : ADFULD1 port map( A => mult_21_C243_n351, B => 
                           mult_21_C243_n353, CI => mult_21_C243_n378, CO => 
                           mult_21_C243_n346, S => mult_21_C243_n347);
   mult_21_C243_U336 : ADFULD1 port map( A => mult_21_C243_n376, B => 
                           mult_21_C243_n349, CI => mult_21_C243_n347, CO => 
                           mult_21_C243_n344, S => mult_21_C243_n345);
   mult_21_C243_U334 : EXOR3D1 port map( A1 => mult_21_C243_n1097, A2 => 
                           mult_21_C243_n1279, A3 => mult_21_C243_n1207, Z => 
                           mult_21_C243_n342);
   mult_21_C243_U333 : EXOR3D1 port map( A1 => mult_21_C243_n1253, A2 => 
                           mult_21_C243_n1127, A3 => mult_21_C243_n1099, Z => 
                           mult_21_C243_n341);
   mult_21_C243_U332 : EXOR3D1 port map( A1 => mult_21_C243_n1103, A2 => 
                           mult_21_C243_n1117, A3 => mult_21_C243_n1109, Z => 
                           mult_21_C243_n340);
   mult_21_C243_U331 : EXOR3D1 port map( A1 => mult_21_C243_n1139, A2 => 
                           mult_21_C243_n1229, A3 => mult_21_C243_n1153, Z => 
                           mult_21_C243_n339);
   mult_21_C243_U330 : EXOR3D1 port map( A1 => mult_21_C243_n1187, A2 => 
                           mult_21_C243_n1169, A3 => mult_21_C243_n372, Z => 
                           mult_21_C243_n338);
   mult_21_C243_U329 : EXOR3D1 port map( A1 => mult_21_C243_n368, A2 => 
                           mult_21_C243_n370, A3 => mult_21_C243_n364, Z => 
                           mult_21_C243_n337);
   mult_21_C243_U328 : EXOR3D1 port map( A1 => mult_21_C243_n366, A2 => 
                           mult_21_C243_n343, A3 => mult_21_C243_n362, Z => 
                           mult_21_C243_n336);
   mult_21_C243_U327 : EXOR3D1 port map( A1 => mult_21_C243_n342, A2 => 
                           mult_21_C243_n338, A3 => mult_21_C243_n341, Z => 
                           mult_21_C243_n335);
   mult_21_C243_U326 : EXOR3D1 port map( A1 => mult_21_C243_n339, A2 => 
                           mult_21_C243_n340, A3 => mult_21_C243_n360, Z => 
                           mult_21_C243_n334);
   mult_21_C243_U325 : EXOR3D1 port map( A1 => mult_21_C243_n337, A2 => 
                           mult_21_C243_n358, A3 => mult_21_C243_n336, Z => 
                           mult_21_C243_n333);
   mult_21_C243_U324 : EXOR3D1 port map( A1 => mult_21_C243_n354, A2 => 
                           mult_21_C243_n356, A3 => mult_21_C243_n335, Z => 
                           mult_21_C243_n332);
   mult_21_C243_U323 : EXOR3D1 port map( A1 => mult_21_C243_n352, A2 => 
                           mult_21_C243_n334, A3 => mult_21_C243_n333, Z => 
                           mult_21_C243_n331);
   mult_21_C243_U322 : EXOR3D1 port map( A1 => mult_21_C243_n332, A2 => 
                           mult_21_C243_n350, A3 => mult_21_C243_n348, Z => 
                           mult_21_C243_n330);
   mult_21_C243_U321 : EXOR3D1 port map( A1 => mult_21_C243_n346, A2 => 
                           mult_21_C243_n331, A3 => mult_21_C243_n330, Z => 
                           mult_21_C243_n329);
   mult_21_C243_U313 : EXOR2D1 port map( A1 => mult_21_C243_n303, A2 => 
                           mult_21_C243_n305, Z => N3266);
   mult_21_C243_U305 : EXNOR2D1 port map( A1 => mult_21_C243_n176, A2 => 
                           mult_21_C243_n302, Z => N3267);
   mult_21_C243_U300 : OAI21D1 port map( A1 => mult_21_C243_n297, A2 => 
                           mult_21_C243_n295, B => mult_21_C243_n296, Z => 
                           mult_21_C243_n294);
   mult_21_C243_U299 : EXOR2D1 port map( A1 => mult_21_C243_n297, A2 => 
                           mult_21_C243_n175, Z => N3268);
   mult_21_C243_U291 : EXNOR2D1 port map( A1 => mult_21_C243_n174, A2 => 
                           mult_21_C243_n294, Z => N3269);
   mult_21_C243_U286 : OAI21D1 port map( A1 => mult_21_C243_n289, A2 => 
                           mult_21_C243_n287, B => mult_21_C243_n288, Z => 
                           mult_21_C243_n286);
   mult_21_C243_U284 : EXOR2D1 port map( A1 => mult_21_C243_n173, A2 => 
                           mult_21_C243_n289, Z => N3270);
   mult_21_C243_U279 : OAI21D1 port map( A1 => mult_21_C243_n285, A2 => 
                           mult_21_C243_n283, B => mult_21_C243_n284, Z => 
                           mult_21_C243_n282);
   mult_21_C243_U278 : EXOR2D1 port map( A1 => mult_21_C243_n172, A2 => 
                           mult_21_C243_n285, Z => N3271);
   mult_21_C243_U273 : OAI21D1 port map( A1 => mult_21_C243_n280, A2 => 
                           mult_21_C243_n284, B => mult_21_C243_n281, Z => 
                           mult_21_C243_n279);
   mult_21_C243_U271 : AOI21D1 port map( A1 => mult_21_C243_n278, A2 => 
                           mult_21_C243_n286, B => mult_21_C243_n279, Z => 
                           mult_21_C243_n277);
   mult_21_C243_U269 : EXNOR2D1 port map( A1 => mult_21_C243_n282, A2 => 
                           mult_21_C243_n171, Z => N3272);
   mult_21_C243_U262 : AOI21D1 port map( A1 => mult_21_C243_n276, A2 => 
                           mult_21_C243_n1527, B => mult_21_C243_n273, Z => 
                           mult_21_C243_n271);
   mult_21_C243_U261 : EXNOR2D1 port map( A1 => mult_21_C243_n276, A2 => 
                           mult_21_C243_n170, Z => N3273);
   mult_21_C243_U254 : AOI21D1 port map( A1 => mult_21_C243_n1524, A2 => 
                           mult_21_C243_n273, B => mult_21_C243_n268, Z => 
                           mult_21_C243_n266);
   mult_21_C243_U252 : OAI21D1 port map( A1 => mult_21_C243_n265, A2 => 
                           mult_21_C243_n277, B => mult_21_C243_n266, Z => 
                           mult_21_C243_n264);
   mult_21_C243_U250 : EXOR2D1 port map( A1 => mult_21_C243_n271, A2 => 
                           mult_21_C243_n169, Z => N3274);
   mult_21_C243_U245 : OAI21D1 port map( A1 => mult_21_C243_n263, A2 => 
                           mult_21_C243_n261, B => mult_21_C243_n262, Z => 
                           mult_21_C243_n260);
   mult_21_C243_U244 : EXOR2D1 port map( A1 => mult_21_C243_n263, A2 => 
                           mult_21_C243_n168, Z => N3275);
   mult_21_C243_U239 : OAI21D1 port map( A1 => mult_21_C243_n258, A2 => 
                           mult_21_C243_n262, B => mult_21_C243_n259, Z => 
                           mult_21_C243_n257);
   mult_21_C243_U237 : AOI21D1 port map( A1 => mult_21_C243_n256, A2 => 
                           mult_21_C243_n264, B => mult_21_C243_n257, Z => 
                           mult_21_C243_n255);
   mult_21_C243_U235 : EXNOR2D1 port map( A1 => mult_21_C243_n260, A2 => 
                           mult_21_C243_n167, Z => N3276);
   mult_21_C243_U228 : AOI21D1 port map( A1 => mult_21_C243_n254, A2 => 
                           mult_21_C243_n1529, B => mult_21_C243_n251, Z => 
                           mult_21_C243_n249);
   mult_21_C243_U227 : EXNOR2D1 port map( A1 => mult_21_C243_n254, A2 => 
                           mult_21_C243_n166, Z => N3277);
   mult_21_C243_U220 : AOI21D1 port map( A1 => mult_21_C243_n1530, A2 => 
                           mult_21_C243_n251, B => mult_21_C243_n246, Z => 
                           mult_21_C243_n244);
   mult_21_C243_U218 : OAI21D1 port map( A1 => mult_21_C243_n255, A2 => 
                           mult_21_C243_n243, B => mult_21_C243_n244, Z => 
                           mult_21_C243_n242);
   mult_21_C243_U216 : EXOR2D1 port map( A1 => mult_21_C243_n249, A2 => 
                           mult_21_C243_n165, Z => N3278);
   mult_21_C243_U211 : OAI21D1 port map( A1 => mult_21_C243_n241, A2 => 
                           mult_21_C243_n239, B => mult_21_C243_n240, Z => 
                           mult_21_C243_n238);
   mult_21_C243_U210 : EXOR2D1 port map( A1 => mult_21_C243_n241, A2 => 
                           mult_21_C243_n164, Z => N3279);
   mult_21_C243_U205 : OAI21D1 port map( A1 => mult_21_C243_n236, A2 => 
                           mult_21_C243_n240, B => mult_21_C243_n237, Z => 
                           mult_21_C243_n235);
   mult_21_C243_U203 : AOI21D1 port map( A1 => mult_21_C243_n242, A2 => 
                           mult_21_C243_n234, B => mult_21_C243_n235, Z => 
                           mult_21_C243_n233);
   mult_21_C243_U201 : EXNOR2D1 port map( A1 => mult_21_C243_n238, A2 => 
                           mult_21_C243_n163, Z => N3280);
   mult_21_C243_U194 : AOI21D1 port map( A1 => mult_21_C243_n232, A2 => 
                           mult_21_C243_n313, B => mult_21_C243_n229, Z => 
                           mult_21_C243_n227);
   mult_21_C243_U193 : EXNOR2D1 port map( A1 => mult_21_C243_n232, A2 => 
                           mult_21_C243_n162, Z => N3281);
   mult_21_C243_U188 : OAI21D1 port map( A1 => mult_21_C243_n225, A2 => 
                           mult_21_C243_n231, B => mult_21_C243_n226, Z => 
                           mult_21_C243_n224);
   mult_21_C243_U186 : AOI21D1 port map( A1 => mult_21_C243_n232, A2 => 
                           mult_21_C243_n223, B => mult_21_C243_n224, Z => 
                           mult_21_C243_n222);
   mult_21_C243_U185 : EXOR2D1 port map( A1 => mult_21_C243_n227, A2 => 
                           mult_21_C243_n161, Z => N3282);
   mult_21_C243_U178 : AOI21D1 port map( A1 => mult_21_C243_n224, A2 => 
                           mult_21_C243_n1528, B => mult_21_C243_n219, Z => 
                           mult_21_C243_n217);
   mult_21_C243_U176 : OAI21D1 port map( A1 => mult_21_C243_n233, A2 => 
                           mult_21_C243_n216, B => mult_21_C243_n217, Z => 
                           mult_21_C243_n215);
   mult_21_C243_U174 : EXOR2D1 port map( A1 => mult_21_C243_n222, A2 => 
                           mult_21_C243_n160, Z => N3283);
   mult_21_C243_U165 : OAI21D1 port map( A1 => mult_21_C243_n214, A2 => 
                           mult_21_C243_n208, B => mult_21_C243_n209, Z => 
                           mult_21_C243_n207);
   mult_21_C243_U164 : EXOR2D1 port map( A1 => mult_21_C243_n214, A2 => 
                           mult_21_C243_n159, Z => N3284);
   mult_21_C243_U157 : AOI21D1 port map( A1 => mult_21_C243_n1525, A2 => 
                           mult_21_C243_n211, B => mult_21_C243_n204, Z => 
                           mult_21_C243_n202);
   mult_21_C243_U155 : OAI21D1 port map( A1 => mult_21_C243_n214, A2 => 
                           mult_21_C243_n201, B => mult_21_C243_n202, Z => 
                           mult_21_C243_n200);
   mult_21_C243_U154 : EXNOR2D1 port map( A1 => mult_21_C243_n207, A2 => 
                           mult_21_C243_n158, Z => N3285);
   mult_21_C243_U147 : AOI21D1 port map( A1 => mult_21_C243_n200, A2 => 
                           mult_21_C243_n1526, B => mult_21_C243_n197, Z => 
                           mult_21_C243_n195);
   mult_21_C243_U146 : EXNOR2D1 port map( A1 => mult_21_C243_n200, A2 => 
                           mult_21_C243_n157, Z => N3286);
   mult_21_C243_U137 : OAI21D1 port map( A1 => mult_21_C243_n202, A2 => 
                           mult_21_C243_n189, B => mult_21_C243_n190, Z => 
                           mult_21_C243_n188);
   mult_21_C243_U134 : EXOR2D1 port map( A1 => mult_21_C243_n195, A2 => 
                           mult_21_C243_n156, Z => N3287);
   mult_21_C243_U132 : ADFULD1 port map( A => mult_21_C243_n531, B => 
                           mult_21_C243_n552, CI => mult_21_C243_n1521, CO => 
                           mult_21_C243_n185, S => N3288);
   mult_21_C243_U131 : ADFULD1 port map( A => mult_21_C243_n507, B => 
                           mult_21_C243_n530, CI => mult_21_C243_n185, CO => 
                           mult_21_C243_n184, S => N3289);
   mult_21_C243_U130 : ADFULD1 port map( A => mult_21_C243_n483, B => 
                           mult_21_C243_n506, CI => mult_21_C243_n184, CO => 
                           mult_21_C243_n183, S => N3290);
   mult_21_C243_U129 : ADFULD1 port map( A => mult_21_C243_n457, B => 
                           mult_21_C243_n482, CI => mult_21_C243_n183, CO => 
                           mult_21_C243_n182, S => N3291);
   mult_21_C243_U128 : ADFULD1 port map( A => mult_21_C243_n431, B => 
                           mult_21_C243_n456, CI => mult_21_C243_n182, CO => 
                           mult_21_C243_n181, S => N3292);
   mult_21_C243_U127 : ADFULD1 port map( A => mult_21_C243_n403, B => 
                           mult_21_C243_n430, CI => mult_21_C243_n181, CO => 
                           mult_21_C243_n180, S => N3293);
   mult_21_C243_U126 : ADFULD1 port map( A => mult_21_C243_n375, B => 
                           mult_21_C243_n402, CI => mult_21_C243_n180, CO => 
                           mult_21_C243_n179, S => N3294);
   mult_21_C243_U125 : ADFULD1 port map( A => mult_21_C243_n345, B => 
                           mult_21_C243_n374, CI => mult_21_C243_n179, CO => 
                           mult_21_C243_n178, S => N3295);
   mult_21_C245_U1390 : INVD1 port map( A => N3008, Z => mult_21_C245_n1066);
   mult_21_C245_U1389 : INVD1 port map( A => N3137, Z => mult_21_C245_n1544);
   mult_21_C245_U1388 : AO21D1 port map( A1 => N3006, A2 => N3007, B => 
                           mult_21_C245_n1066, Z => mult_21_C245_n105);
   mult_21_C245_U1387 : INVD1 port map( A => N3006, Z => mult_21_C245_n1067);
   mult_21_C245_U1386 : AO21D1 port map( A1 => N3004, A2 => N3005, B => 
                           mult_21_C245_n1067, Z => mult_21_C245_n101);
   mult_21_C245_U1385 : EXOR2D1 port map( A1 => mult_21_C245_n1307, A2 => 
                           mult_21_C245_n1337, Z => mult_21_C245_n343);
   mult_21_C245_U1384 : INVD1 port map( A => N3004, Z => mult_21_C245_n1068);
   mult_21_C245_U1383 : AO21D1 port map( A1 => N3002, A2 => N3003, B => 
                           mult_21_C245_n1068, Z => mult_21_C245_n96);
   mult_21_C245_U1382 : ADHALFDL port map( A => mult_21_C245_n1309, B => 
                           mult_21_C245_n1339, CO => mult_21_C245_n400, S => 
                           mult_21_C245_n401);
   mult_21_C245_U1381 : AO21D1 port map( A1 => N3000, A2 => N3001, B => 
                           mult_21_C245_n1069, Z => mult_21_C245_n91);
   mult_21_C245_U1380 : INVD1 port map( A => N3002, Z => mult_21_C245_n1069);
   mult_21_C245_U1379 : OAI21D1 port map( A1 => N3000, A2 => N3001, B => 
                           mult_21_C245_n1069, Z => mult_21_C245_n89);
   mult_21_C245_U1378 : ADHALFDL port map( A => mult_21_C245_n1311, B => 
                           mult_21_C245_n1341, CO => mult_21_C245_n454, S => 
                           mult_21_C245_n455);
   mult_21_C245_U1377 : ADHALFDL port map( A => mult_21_C245_n1313, B => 
                           mult_21_C245_n1343, CO => mult_21_C245_n504, S => 
                           mult_21_C245_n505);
   mult_21_C245_U1376 : AO21D1 port map( A1 => N2998, A2 => N2999, B => 
                           mult_21_C245_n1070, Z => mult_21_C245_n86);
   mult_21_C245_U1375 : INVD1 port map( A => N3000, Z => mult_21_C245_n1070);
   mult_21_C245_U1374 : OAI21D1 port map( A1 => N2998, A2 => N2999, B => 
                           mult_21_C245_n1070, Z => mult_21_C245_n84);
   mult_21_C245_U1373 : AO21D1 port map( A1 => N2996, A2 => N2997, B => 
                           mult_21_C245_n1071, Z => mult_21_C245_n81);
   mult_21_C245_U1372 : INVD1 port map( A => N2998, Z => mult_21_C245_n1071);
   mult_21_C245_U1371 : OAI21D1 port map( A1 => N2996, A2 => N2997, B => 
                           mult_21_C245_n1071, Z => mult_21_C245_n79);
   mult_21_C245_U1370 : EXNOR2D1 port map( A1 => N2998, A2 => N2999, Z => 
                           mult_21_C245_n88);
   mult_21_C245_U1369 : AO21D1 port map( A1 => N2994, A2 => N2995, B => 
                           mult_21_C245_n1072, Z => mult_21_C245_n76);
   mult_21_C245_U1368 : OAI21D1 port map( A1 => N2986, A2 => N2987, B => 
                           mult_21_C245_n1076, Z => mult_21_C245_n42);
   mult_21_C245_U1367 : INVD1 port map( A => N2996, Z => mult_21_C245_n1072);
   mult_21_C245_U1366 : OAI21D1 port map( A1 => N2994, A2 => N2995, B => 
                           mult_21_C245_n1072, Z => mult_21_C245_n73);
   mult_21_C245_U1365 : INVD1 port map( A => N2988, Z => mult_21_C245_n1076);
   mult_21_C245_U1364 : AO21D1 port map( A1 => N2986, A2 => N2987, B => 
                           mult_21_C245_n1076, Z => mult_21_C245_n45);
   mult_21_C245_U1363 : OAI21D1 port map( A1 => N2992, A2 => N2993, B => 
                           mult_21_C245_n1073, Z => mult_21_C245_n66);
   mult_21_C245_U1362 : INVD1 port map( A => N2994, Z => mult_21_C245_n1073);
   mult_21_C245_U1361 : OAI21D1 port map( A1 => N2990, A2 => N2991, B => 
                           mult_21_C245_n1074, Z => mult_21_C245_n58);
   mult_21_C245_U1360 : INVD1 port map( A => N2992, Z => mult_21_C245_n1074);
   mult_21_C245_U1359 : AO21D1 port map( A1 => N2992, A2 => N2993, B => 
                           mult_21_C245_n1073, Z => mult_21_C245_n69);
   mult_21_C245_U1358 : AO21D1 port map( A1 => N2990, A2 => N2991, B => 
                           mult_21_C245_n1074, Z => mult_21_C245_n61);
   mult_21_C245_U1357 : OAI21D1 port map( A1 => N2988, A2 => N2989, B => 
                           mult_21_C245_n1075, Z => mult_21_C245_n50);
   mult_21_C245_U1356 : AO21D1 port map( A1 => N2984, A2 => N2985, B => 
                           mult_21_C245_n1077, Z => mult_21_C245_n38);
   mult_21_C245_U1355 : AO21D1 port map( A1 => N2980, A2 => N2981, B => 
                           mult_21_C245_n1079, Z => mult_21_C245_n22);
   mult_21_C245_U1354 : ADHALFDL port map( A => mult_21_C245_n1315, B => 
                           mult_21_C245_n1345, CO => mult_21_C245_n550, S => 
                           mult_21_C245_n551);
   mult_21_C245_U1353 : INVD1 port map( A => N2990, Z => mult_21_C245_n1075);
   mult_21_C245_U1352 : AO21D1 port map( A1 => N2988, A2 => N2989, B => 
                           mult_21_C245_n1075, Z => mult_21_C245_n53);
   mult_21_C245_U1351 : EXNOR2D1 port map( A1 => N2996, A2 => N2997, Z => 
                           mult_21_C245_n83);
   mult_21_C245_U1350 : INVD1 port map( A => N2977, Z => mult_21_C245_n8);
   mult_21_C245_U1349 : AO21D1 port map( A1 => N2982, A2 => N2983, B => 
                           mult_21_C245_n1078, Z => mult_21_C245_n30);
   mult_21_C245_U1348 : INVD1 port map( A => mult_21_C245_n1544, Z => 
                           mult_21_C245_n1543);
   mult_21_C245_U1347 : EXNOR2D1 port map( A1 => N2994, A2 => N2995, Z => 
                           mult_21_C245_n78);
   mult_21_C245_U1346 : AO21D1 port map( A1 => N2978, A2 => N2979, B => 
                           mult_21_C245_n1080, Z => mult_21_C245_n14);
   mult_21_C245_U1345 : EXNOR2D1 port map( A1 => N2986, A2 => N2987, Z => 
                           mult_21_C245_n48);
   mult_21_C245_U1344 : INVD1 port map( A => N2982, Z => mult_21_C245_n1079);
   mult_21_C245_U1343 : EXNOR2D1 port map( A1 => N2992, A2 => N2993, Z => 
                           mult_21_C245_n71);
   mult_21_C245_U1342 : EXNOR2D1 port map( A1 => N2990, A2 => N2991, Z => 
                           mult_21_C245_n63);
   mult_21_C245_U1341 : INVD1 port map( A => N2986, Z => mult_21_C245_n1077);
   mult_21_C245_U1340 : INVD1 port map( A => N2978, Z => mult_21_C245_n6);
   mult_21_C245_U1339 : NAN2D1 port map( A1 => N2977, A2 => mult_21_C245_n6, Z 
                           => mult_21_C245_n3);
   mult_21_C245_U1338 : INVD1 port map( A => N2984, Z => mult_21_C245_n1078);
   mult_21_C245_U1337 : EXNOR2D1 port map( A1 => N2988, A2 => N2989, Z => 
                           mult_21_C245_n56);
   mult_21_C245_U1336 : INVD1 port map( A => N2980, Z => mult_21_C245_n1080);
   mult_21_C245_U1335 : OA21D1 port map( A1 => N2982, A2 => N2983, B => 
                           mult_21_C245_n1078, Z => mult_21_C245_n1537);
   mult_21_C245_U1334 : ADHALFDL port map( A => mult_21_C245_n1325, B => 
                           mult_21_C245_n1355, CO => mult_21_C245_n720, S => 
                           mult_21_C245_n721);
   mult_21_C245_U1333 : ADHALFDL port map( A => mult_21_C245_n1321, B => 
                           mult_21_C245_n1351, CO => mult_21_C245_n664, S => 
                           mult_21_C245_n665);
   mult_21_C245_U1332 : ADHALFDL port map( A => mult_21_C245_n1319, B => 
                           mult_21_C245_n1349, CO => mult_21_C245_n630, S => 
                           mult_21_C245_n631);
   mult_21_C245_U1331 : ADHALFDL port map( A => mult_21_C245_n1327, B => 
                           mult_21_C245_n1357, CO => mult_21_C245_n742, S => 
                           mult_21_C245_n743);
   mult_21_C245_U1330 : ADHALFDL port map( A => mult_21_C245_n1317, B => 
                           mult_21_C245_n1347, CO => mult_21_C245_n592, S => 
                           mult_21_C245_n593);
   mult_21_C245_U1329 : EXOR2D1 port map( A1 => N2984, A2 => N2985, Z => 
                           mult_21_C245_n1536);
   mult_21_C245_U1328 : EXOR2D1 port map( A1 => N2980, A2 => N2981, Z => 
                           mult_21_C245_n1535);
   mult_21_C245_U1327 : EXOR2D1 port map( A1 => N2982, A2 => N2983, Z => 
                           mult_21_C245_n1534);
   mult_21_C245_U1326 : ADHALFDL port map( A => mult_21_C245_n1323, B => 
                           mult_21_C245_n1353, CO => mult_21_C245_n694, S => 
                           mult_21_C245_n695);
   mult_21_C245_U1325 : EXOR2D1 port map( A1 => N2978, A2 => N2979, Z => 
                           mult_21_C245_n1533);
   mult_21_C245_U1324 : ADHALFDL port map( A => mult_21_C245_n1329, B => 
                           mult_21_C245_n1359, CO => mult_21_C245_n760, S => 
                           mult_21_C245_n761);
   mult_21_C245_U1323 : ADHALFDL port map( A => mult_21_C245_n1098, B => 
                           mult_21_C245_n1081, CO => mult_21_C245_n372, S => 
                           mult_21_C245_n373);
   mult_21_C245_U1322 : ADHALFDL port map( A => mult_21_C245_n1102, B => 
                           mult_21_C245_n1082, CO => mult_21_C245_n428, S => 
                           mult_21_C245_n429);
   mult_21_C245_U1321 : ADHALFDL port map( A => mult_21_C245_n1108, B => 
                           mult_21_C245_n1083, CO => mult_21_C245_n480, S => 
                           mult_21_C245_n481);
   mult_21_C245_U1320 : ADHALFDL port map( A => mult_21_C245_n1116, B => 
                           mult_21_C245_n1084, CO => mult_21_C245_n528, S => 
                           mult_21_C245_n529);
   mult_21_C245_U1319 : ADHALFDL port map( A => mult_21_C245_n1126, B => 
                           mult_21_C245_n1085, CO => mult_21_C245_n572, S => 
                           mult_21_C245_n573);
   mult_21_C245_U1318 : INVD1 port map( A => mult_21_C245_n1367, Z => 
                           mult_21_C245_n303);
   mult_21_C245_U1317 : ADHALFDL port map( A => mult_21_C245_n1138, B => 
                           mult_21_C245_n1086, CO => mult_21_C245_n612, S => 
                           mult_21_C245_n613);
   mult_21_C245_U1316 : ADHALFDL port map( A => mult_21_C245_n1186, B => 
                           mult_21_C245_n1089, CO => mult_21_C245_n708, S => 
                           mult_21_C245_n709);
   mult_21_C245_U1315 : ADHALFDL port map( A => mult_21_C245_n1228, B => 
                           mult_21_C245_n1091, CO => mult_21_C245_n752, S => 
                           mult_21_C245_n753);
   mult_21_C245_U1314 : ADHALFDL port map( A => mult_21_C245_n1152, B => 
                           mult_21_C245_n1087, CO => mult_21_C245_n648, S => 
                           mult_21_C245_n649);
   mult_21_C245_U1313 : ADHALFDL port map( A => mult_21_C245_n1168, B => 
                           mult_21_C245_n1088, CO => mult_21_C245_n680, S => 
                           mult_21_C245_n681);
   mult_21_C245_U1312 : ADHALFDL port map( A => mult_21_C245_n1206, B => 
                           mult_21_C245_n1090, CO => mult_21_C245_n732, S => 
                           mult_21_C245_n733);
   mult_21_C245_U1311 : INVD1 port map( A => mult_21_C245_n1537, Z => 
                           mult_21_C245_n1540);
   mult_21_C245_U1310 : ADHALFDL port map( A => mult_21_C245_n1306, B => 
                           mult_21_C245_n1094, CO => mult_21_C245_n788, S => 
                           mult_21_C245_n789);
   mult_21_C245_U1309 : ADHALFDL port map( A => mult_21_C245_n1333, B => 
                           mult_21_C245_n1363, CO => mult_21_C245_n784, S => 
                           mult_21_C245_n785);
   mult_21_C245_U1308 : INVD1 port map( A => mult_21_C245_n1536, Z => 
                           mult_21_C245_n1538);
   mult_21_C245_U1307 : ADHALFDL port map( A => mult_21_C245_n1252, B => 
                           mult_21_C245_n1092, CO => mult_21_C245_n768, S => 
                           mult_21_C245_n769);
   mult_21_C245_U1306 : INVD1 port map( A => mult_21_C245_n1534, Z => 
                           mult_21_C245_n1539);
   mult_21_C245_U1305 : ADHALFDL port map( A => mult_21_C245_n1331, B => 
                           mult_21_C245_n1361, CO => mult_21_C245_n774, S => 
                           mult_21_C245_n775);
   mult_21_C245_U1304 : INVD1 port map( A => mult_21_C245_n1535, Z => 
                           mult_21_C245_n1541);
   mult_21_C245_U1303 : NOR2D1 port map( A1 => mult_21_C245_n1537, A2 => 
                           mult_21_C245_n30, Z => mult_21_C245_n1093);
   mult_21_C245_U1302 : ADHALFDL port map( A => mult_21_C245_n1336, B => 
                           mult_21_C245_n1095, CO => mult_21_C245_n792, S => 
                           mult_21_C245_n793);
   mult_21_C245_U1301 : ADHALFDL port map( A => mult_21_C245_n1335, B => 
                           mult_21_C245_n1365, CO => mult_21_C245_n790, S => 
                           mult_21_C245_n791);
   mult_21_C245_U1300 : EXOR2D1 port map( A1 => mult_21_C245_n329, A2 => 
                           mult_21_C245_n344, Z => mult_21_C245_n155);
   mult_21_C245_U1299 : EXOR2D1 port map( A1 => mult_21_C245_n178, A2 => 
                           mult_21_C245_n155, Z => N3328);
   mult_21_C245_U1298 : INVD1 port map( A => mult_21_C245_n1533, Z => 
                           mult_21_C245_n1542);
   mult_21_C245_U1297 : NOR2D1 port map( A1 => mult_21_C245_n303, A2 => 
                           mult_21_C245_n305, Z => mult_21_C245_n302);
   mult_21_C245_U1296 : NAN2D1 port map( A1 => mult_21_C245_n1368, A2 => 
                           mult_21_C245_n1096, Z => mult_21_C245_n305);
   mult_21_C245_U1295 : NAN2D1 port map( A1 => mult_21_C245_n791, A2 => 
                           mult_21_C245_n792, Z => mult_21_C245_n296);
   mult_21_C245_U1294 : NAN2D1 port map( A1 => mult_21_C245_n783, A2 => 
                           mult_21_C245_n786, Z => mult_21_C245_n288);
   mult_21_C245_U1293 : NOR2D1 port map( A1 => mult_21_C245_n791, A2 => 
                           mult_21_C245_n792, Z => mult_21_C245_n295);
   mult_21_C245_U1292 : NOR2D1 port map( A1 => mult_21_C245_n783, A2 => 
                           mult_21_C245_n786, Z => mult_21_C245_n287);
   mult_21_C245_U1291 : NAN2D1 port map( A1 => mult_21_C245_n777, A2 => 
                           mult_21_C245_n782, Z => mult_21_C245_n284);
   mult_21_C245_U1290 : NAN2D1 port map( A1 => mult_21_C245_n793, A2 => 
                           mult_21_C245_n1366, Z => mult_21_C245_n301);
   mult_21_C245_U1289 : NAN2D1 port map( A1 => mult_21_C245_n787, A2 => 
                           mult_21_C245_n789, Z => mult_21_C245_n293);
   mult_21_C245_U1288 : NOR2D1 port map( A1 => mult_21_C245_n777, A2 => 
                           mult_21_C245_n782, Z => mult_21_C245_n283);
   mult_21_C245_U1287 : OR2D1 port map( A1 => mult_21_C245_n793, A2 => 
                           mult_21_C245_n1366, Z => mult_21_C245_n1532);
   mult_21_C245_U1286 : OR2D1 port map( A1 => mult_21_C245_n787, A2 => 
                           mult_21_C245_n789, Z => mult_21_C245_n1531);
   mult_21_C245_U1285 : NAN2D1 port map( A1 => mult_21_C245_n1532, A2 => 
                           mult_21_C245_n301, Z => mult_21_C245_n176);
   mult_21_C245_U1284 : INVD1 port map( A => mult_21_C245_n295, Z => 
                           mult_21_C245_n326);
   mult_21_C245_U1283 : NAN2D1 port map( A1 => mult_21_C245_n326, A2 => 
                           mult_21_C245_n296, Z => mult_21_C245_n175);
   mult_21_C245_U1282 : NAN2D1 port map( A1 => mult_21_C245_n1531, A2 => 
                           mult_21_C245_n293, Z => mult_21_C245_n174);
   mult_21_C245_U1281 : INVD1 port map( A => mult_21_C245_n287, Z => 
                           mult_21_C245_n324);
   mult_21_C245_U1280 : NAN2D1 port map( A1 => mult_21_C245_n324, A2 => 
                           mult_21_C245_n288, Z => mult_21_C245_n173);
   mult_21_C245_U1279 : INVD1 port map( A => mult_21_C245_n283, Z => 
                           mult_21_C245_n323);
   mult_21_C245_U1278 : NAN2D1 port map( A1 => mult_21_C245_n323, A2 => 
                           mult_21_C245_n284, Z => mult_21_C245_n172);
   mult_21_C245_U1277 : INVD1 port map( A => mult_21_C245_n280, Z => 
                           mult_21_C245_n322);
   mult_21_C245_U1276 : NAN2D1 port map( A1 => mult_21_C245_n322, A2 => 
                           mult_21_C245_n281, Z => mult_21_C245_n171);
   mult_21_C245_U1275 : NAN2D1 port map( A1 => mult_21_C245_n697, A2 => 
                           mult_21_C245_n710, Z => mult_21_C245_n240);
   mult_21_C245_U1274 : NAN2D1 port map( A1 => mult_21_C245_n633, A2 => 
                           mult_21_C245_n650, Z => mult_21_C245_n221);
   mult_21_C245_U1273 : NAN2D1 port map( A1 => mult_21_C245_n711, A2 => 
                           mult_21_C245_n722, Z => mult_21_C245_n248);
   mult_21_C245_U1272 : NOR2D1 port map( A1 => mult_21_C245_n697, A2 => 
                           mult_21_C245_n710, Z => mult_21_C245_n239);
   mult_21_C245_U1271 : NOR2D1 port map( A1 => mult_21_C245_n615, A2 => 
                           mult_21_C245_n632, Z => mult_21_C245_n208);
   mult_21_C245_U1270 : NAN2D1 port map( A1 => mult_21_C245_n735, A2 => 
                           mult_21_C245_n744, Z => mult_21_C245_n259);
   mult_21_C245_U1269 : NAN2D1 port map( A1 => mult_21_C245_n771, A2 => 
                           mult_21_C245_n776, Z => mult_21_C245_n281);
   mult_21_C245_U1268 : NAN2D1 port map( A1 => mult_21_C245_n615, A2 => 
                           mult_21_C245_n632, Z => mult_21_C245_n209);
   mult_21_C245_U1267 : OR2D1 port map( A1 => mult_21_C245_n711, A2 => 
                           mult_21_C245_n722, Z => mult_21_C245_n1530);
   mult_21_C245_U1266 : NAN2D1 port map( A1 => mult_21_C245_n745, A2 => 
                           mult_21_C245_n754, Z => mult_21_C245_n262);
   mult_21_C245_U1265 : OR2D1 port map( A1 => mult_21_C245_n723, A2 => 
                           mult_21_C245_n734, Z => mult_21_C245_n1529);
   mult_21_C245_U1264 : OR2D1 port map( A1 => mult_21_C245_n633, A2 => 
                           mult_21_C245_n650, Z => mult_21_C245_n1528);
   mult_21_C245_U1263 : NAN2D1 port map( A1 => mult_21_C245_n595, A2 => 
                           mult_21_C245_n614, Z => mult_21_C245_n206);
   mult_21_C245_U1262 : OR2D1 port map( A1 => mult_21_C245_n763, A2 => 
                           mult_21_C245_n770, Z => mult_21_C245_n1527);
   mult_21_C245_U1261 : NAN2D1 port map( A1 => mult_21_C245_n651, A2 => 
                           mult_21_C245_n666, Z => mult_21_C245_n226);
   mult_21_C245_U1260 : NAN2D1 port map( A1 => mult_21_C245_n723, A2 => 
                           mult_21_C245_n734, Z => mult_21_C245_n253);
   mult_21_C245_U1259 : NAN2D1 port map( A1 => mult_21_C245_n575, A2 => 
                           mult_21_C245_n594, Z => mult_21_C245_n199);
   mult_21_C245_U1258 : OR2D1 port map( A1 => mult_21_C245_n575, A2 => 
                           mult_21_C245_n594, Z => mult_21_C245_n1526);
   mult_21_C245_U1257 : NAN2D1 port map( A1 => mult_21_C245_n763, A2 => 
                           mult_21_C245_n770, Z => mult_21_C245_n275);
   mult_21_C245_U1256 : NOR2D1 port map( A1 => mult_21_C245_n735, A2 => 
                           mult_21_C245_n744, Z => mult_21_C245_n258);
   mult_21_C245_U1255 : NOR2D1 port map( A1 => mult_21_C245_n745, A2 => 
                           mult_21_C245_n754, Z => mult_21_C245_n261);
   mult_21_C245_U1254 : NOR2D1 port map( A1 => mult_21_C245_n771, A2 => 
                           mult_21_C245_n776, Z => mult_21_C245_n280);
   mult_21_C245_U1253 : OR2D1 port map( A1 => mult_21_C245_n595, A2 => 
                           mult_21_C245_n614, Z => mult_21_C245_n1525);
   mult_21_C245_U1252 : OA21M20D1 port map( A1 => mult_21_C245_n1532, A2 => 
                           mult_21_C245_n302, B => mult_21_C245_n301, Z => 
                           mult_21_C245_n297);
   mult_21_C245_U1251 : NOR2D1 port map( A1 => mult_21_C245_n651, A2 => 
                           mult_21_C245_n666, Z => mult_21_C245_n225);
   mult_21_C245_U1250 : OA21M20D1 port map( A1 => mult_21_C245_n1531, A2 => 
                           mult_21_C245_n294, B => mult_21_C245_n293, Z => 
                           mult_21_C245_n289);
   mult_21_C245_U1249 : NOR2D1 port map( A1 => mult_21_C245_n280, A2 => 
                           mult_21_C245_n283, Z => mult_21_C245_n278);
   mult_21_C245_U1248 : NAN2D1 port map( A1 => mult_21_C245_n755, A2 => 
                           mult_21_C245_n762, Z => mult_21_C245_n270);
   mult_21_C245_U1247 : OR2D1 port map( A1 => mult_21_C245_n755, A2 => 
                           mult_21_C245_n762, Z => mult_21_C245_n1524);
   mult_21_C245_U1246 : INVD1 port map( A => mult_21_C245_n286, Z => 
                           mult_21_C245_n285);
   mult_21_C245_U1245 : NAN2D1 port map( A1 => mult_21_C245_n1527, A2 => 
                           mult_21_C245_n275, Z => mult_21_C245_n170);
   mult_21_C245_U1244 : NAN2D1 port map( A1 => mult_21_C245_n1524, A2 => 
                           mult_21_C245_n270, Z => mult_21_C245_n169);
   mult_21_C245_U1243 : INVD1 port map( A => mult_21_C245_n277, Z => 
                           mult_21_C245_n276);
   mult_21_C245_U1242 : INVD1 port map( A => mult_21_C245_n261, Z => 
                           mult_21_C245_n319);
   mult_21_C245_U1241 : NAN2D1 port map( A1 => mult_21_C245_n319, A2 => 
                           mult_21_C245_n262, Z => mult_21_C245_n168);
   mult_21_C245_U1240 : INVD1 port map( A => mult_21_C245_n258, Z => 
                           mult_21_C245_n318);
   mult_21_C245_U1239 : NAN2D1 port map( A1 => mult_21_C245_n318, A2 => 
                           mult_21_C245_n259, Z => mult_21_C245_n167);
   mult_21_C245_U1238 : NAN2D1 port map( A1 => mult_21_C245_n1529, A2 => 
                           mult_21_C245_n253, Z => mult_21_C245_n166);
   mult_21_C245_U1237 : INVD1 port map( A => mult_21_C245_n239, Z => 
                           mult_21_C245_n315);
   mult_21_C245_U1236 : NAN2D1 port map( A1 => mult_21_C245_n315, A2 => 
                           mult_21_C245_n240, Z => mult_21_C245_n164);
   mult_21_C245_U1235 : NAN2D1 port map( A1 => mult_21_C245_n1530, A2 => 
                           mult_21_C245_n248, Z => mult_21_C245_n165);
   mult_21_C245_U1234 : INVD1 port map( A => mult_21_C245_n236, Z => 
                           mult_21_C245_n314);
   mult_21_C245_U1233 : NAN2D1 port map( A1 => mult_21_C245_n314, A2 => 
                           mult_21_C245_n237, Z => mult_21_C245_n163);
   mult_21_C245_U1232 : NAN2D1 port map( A1 => mult_21_C245_n1528, A2 => 
                           mult_21_C245_n221, Z => mult_21_C245_n160);
   mult_21_C245_U1231 : INVD1 port map( A => mult_21_C245_n225, Z => 
                           mult_21_C245_n312);
   mult_21_C245_U1230 : NAN2D1 port map( A1 => mult_21_C245_n312, A2 => 
                           mult_21_C245_n226, Z => mult_21_C245_n161);
   mult_21_C245_U1229 : NAN2D1 port map( A1 => mult_21_C245_n310, A2 => 
                           mult_21_C245_n209, Z => mult_21_C245_n159);
   mult_21_C245_U1228 : NAN2D1 port map( A1 => mult_21_C245_n1525, A2 => 
                           mult_21_C245_n206, Z => mult_21_C245_n158);
   mult_21_C245_U1227 : NAN2D1 port map( A1 => mult_21_C245_n1526, A2 => 
                           mult_21_C245_n199, Z => mult_21_C245_n157);
   mult_21_C245_U1226 : NAN2D1 port map( A1 => mult_21_C245_n1523, A2 => 
                           mult_21_C245_n194, Z => mult_21_C245_n156);
   mult_21_C245_U1225 : NAN2D1 port map( A1 => mult_21_C245_n683, A2 => 
                           mult_21_C245_n696, Z => mult_21_C245_n237);
   mult_21_C245_U1224 : NOR2D1 port map( A1 => mult_21_C245_n667, A2 => 
                           mult_21_C245_n682, Z => mult_21_C245_n230);
   mult_21_C245_U1223 : INVD1 port map( A => mult_21_C245_n208, Z => 
                           mult_21_C245_n310);
   mult_21_C245_U1222 : NAN2D1 port map( A1 => mult_21_C245_n553, A2 => 
                           mult_21_C245_n574, Z => mult_21_C245_n194);
   mult_21_C245_U1221 : NOR2D1 port map( A1 => mult_21_C245_n683, A2 => 
                           mult_21_C245_n696, Z => mult_21_C245_n236);
   mult_21_C245_U1220 : NAN2D1 port map( A1 => mult_21_C245_n1525, A2 => 
                           mult_21_C245_n310, Z => mult_21_C245_n201);
   mult_21_C245_U1219 : NOR2D1 port map( A1 => mult_21_C245_n225, A2 => 
                           mult_21_C245_n230, Z => mult_21_C245_n223);
   mult_21_C245_U1218 : NAN2D1 port map( A1 => mult_21_C245_n667, A2 => 
                           mult_21_C245_n682, Z => mult_21_C245_n231);
   mult_21_C245_U1217 : INVD1 port map( A => mult_21_C245_n253, Z => 
                           mult_21_C245_n251);
   mult_21_C245_U1216 : INVD1 port map( A => mult_21_C245_n199, Z => 
                           mult_21_C245_n197);
   mult_21_C245_U1215 : NAN2D1 port map( A1 => mult_21_C245_n1523, A2 => 
                           mult_21_C245_n1526, Z => mult_21_C245_n189);
   mult_21_C245_U1214 : OR2D1 port map( A1 => mult_21_C245_n553, A2 => 
                           mult_21_C245_n574, Z => mult_21_C245_n1523);
   mult_21_C245_U1213 : INVD1 port map( A => mult_21_C245_n275, Z => 
                           mult_21_C245_n273);
   mult_21_C245_U1212 : INVD1 port map( A => mult_21_C245_n206, Z => 
                           mult_21_C245_n204);
   mult_21_C245_U1211 : INVD1 port map( A => mult_21_C245_n209, Z => 
                           mult_21_C245_n211);
   mult_21_C245_U1210 : NOR2D1 port map( A1 => mult_21_C245_n189, A2 => 
                           mult_21_C245_n201, Z => mult_21_C245_n187);
   mult_21_C245_U1209 : NOR2D1 port map( A1 => mult_21_C245_n236, A2 => 
                           mult_21_C245_n239, Z => mult_21_C245_n234);
   mult_21_C245_U1208 : NOR2D1 port map( A1 => mult_21_C245_n258, A2 => 
                           mult_21_C245_n261, Z => mult_21_C245_n256);
   mult_21_C245_U1207 : INVD1 port map( A => mult_21_C245_n270, Z => 
                           mult_21_C245_n268);
   mult_21_C245_U1206 : NAN2D1 port map( A1 => mult_21_C245_n1524, A2 => 
                           mult_21_C245_n1527, Z => mult_21_C245_n265);
   mult_21_C245_U1205 : INVD1 port map( A => mult_21_C245_n248, Z => 
                           mult_21_C245_n246);
   mult_21_C245_U1204 : NAN2D1 port map( A1 => mult_21_C245_n1530, A2 => 
                           mult_21_C245_n1529, Z => mult_21_C245_n243);
   mult_21_C245_U1203 : INVD1 port map( A => mult_21_C245_n221, Z => 
                           mult_21_C245_n219);
   mult_21_C245_U1202 : NAN2D1 port map( A1 => mult_21_C245_n223, A2 => 
                           mult_21_C245_n1528, Z => mult_21_C245_n216);
   mult_21_C245_U1201 : INVD1 port map( A => mult_21_C245_n264, Z => 
                           mult_21_C245_n263);
   mult_21_C245_U1200 : INVD1 port map( A => mult_21_C245_n231, Z => 
                           mult_21_C245_n229);
   mult_21_C245_U1199 : INVD1 port map( A => mult_21_C245_n230, Z => 
                           mult_21_C245_n313);
   mult_21_C245_U1198 : INVD1 port map( A => mult_21_C245_n255, Z => 
                           mult_21_C245_n254);
   mult_21_C245_U1197 : INVD1 port map( A => mult_21_C245_n242, Z => 
                           mult_21_C245_n241);
   mult_21_C245_U1196 : NAN2D1 port map( A1 => mult_21_C245_n313, A2 => 
                           mult_21_C245_n231, Z => mult_21_C245_n162);
   mult_21_C245_U1195 : INVD1 port map( A => mult_21_C245_n233, Z => 
                           mult_21_C245_n232);
   mult_21_C245_U1194 : INVD1 port map( A => mult_21_C245_n215, Z => 
                           mult_21_C245_n214);
   mult_21_C245_U1193 : OA21M20D1 port map( A1 => mult_21_C245_n1523, A2 => 
                           mult_21_C245_n197, B => mult_21_C245_n194, Z => 
                           mult_21_C245_n190);
   mult_21_C245_U1192 : OR2D1 port map( A1 => mult_21_C245_n1368, A2 => 
                           mult_21_C245_n1096, Z => mult_21_C245_n1522);
   mult_21_C245_U1191 : AO21D1 port map( A1 => mult_21_C245_n215, A2 => 
                           mult_21_C245_n187, B => mult_21_C245_n188, Z => 
                           mult_21_C245_n1521);
   mult_21_C245_U1190 : AND2D1 port map( A1 => mult_21_C245_n1522, A2 => 
                           mult_21_C245_n305, Z => N3297);
   mult_21_C245_U1189 : OAI21D1 port map( A1 => N2984, A2 => N2985, B => 
                           mult_21_C245_n1077, Z => mult_21_C245_n1519);
   mult_21_C245_U1188 : OAI21D1 port map( A1 => N2980, A2 => N2981, B => 
                           mult_21_C245_n1079, Z => mult_21_C245_n1518);
   mult_21_C245_U1187 : OAI21D1 port map( A1 => N2978, A2 => N2979, B => 
                           mult_21_C245_n1080, Z => mult_21_C245_n1517);
   mult_21_C245_U1186 : ADHALFDL port map( A => mult_21_C245_n1278, B => 
                           mult_21_C245_n1093, CO => mult_21_C245_n780, S => 
                           mult_21_C245_n781);
   mult_21_C245_U1135 : EXNOR2D1 port map( A1 => N3000, A2 => N3001, Z => 
                           mult_21_C245_n93);
   mult_21_C245_U1131 : EXNOR2D1 port map( A1 => N3002, A2 => N3003, Z => 
                           mult_21_C245_n98);
   mult_21_C245_U1129 : OAI21D1 port map( A1 => N3002, A2 => N3003, B => 
                           mult_21_C245_n1068, Z => mult_21_C245_n94);
   mult_21_C245_U1127 : EXNOR2D1 port map( A1 => N3004, A2 => N3005, Z => 
                           mult_21_C245_n103);
   mult_21_C245_U1125 : OAI21D1 port map( A1 => N3004, A2 => N3005, B => 
                           mult_21_C245_n1067, Z => mult_21_C245_n99);
   mult_21_C245_U1123 : EXNOR2D1 port map( A1 => N3006, A2 => N3007, Z => 
                           mult_21_C245_n106);
   mult_21_C245_U1121 : OAI21D1 port map( A1 => N3006, A2 => N3007, B => 
                           mult_21_C245_n1066, Z => mult_21_C245_n104);
   mult_21_C245_U1120 : NAN2M1D1 port map( A1 => mult_21_C245_n8, A2 => 
                           mult_21_C245_n1543, Z => mult_21_C245_n1065);
   mult_21_C245_U1119 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1065, Z => 
                           mult_21_C245_n1368);
   mult_21_C245_U1118 : MUXB2DL port map( A0 => N3138, A1 => mult_21_C245_n1543
                           , SL => mult_21_C245_n8, Z => mult_21_C245_n1064);
   mult_21_C245_U1117 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1064, Z => 
                           mult_21_C245_n1367);
   mult_21_C245_U1116 : MUXB2DL port map( A0 => N3139, A1 => N3138, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1063);
   mult_21_C245_U1115 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1063, Z => 
                           mult_21_C245_n1366);
   mult_21_C245_U1114 : MUXB2DL port map( A0 => N3140, A1 => N3139, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1062);
   mult_21_C245_U1113 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1062, Z => 
                           mult_21_C245_n1365);
   mult_21_C245_U1112 : MUXB2DL port map( A0 => N3141, A1 => N3140, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1061);
   mult_21_C245_U1111 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1061, Z => 
                           mult_21_C245_n1364);
   mult_21_C245_U1110 : MUXB2DL port map( A0 => N3142, A1 => N3141, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1060);
   mult_21_C245_U1109 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1060, Z => 
                           mult_21_C245_n1363);
   mult_21_C245_U1108 : MUXB2DL port map( A0 => N3143, A1 => N3142, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1059);
   mult_21_C245_U1107 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1059, Z => 
                           mult_21_C245_n1362);
   mult_21_C245_U1106 : MUXB2DL port map( A0 => N3144, A1 => N3143, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1058);
   mult_21_C245_U1105 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1058, Z => 
                           mult_21_C245_n1361);
   mult_21_C245_U1104 : MUXB2DL port map( A0 => N3145, A1 => N3144, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1057);
   mult_21_C245_U1103 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1057, Z => 
                           mult_21_C245_n1360);
   mult_21_C245_U1102 : MUXB2DL port map( A0 => N3146, A1 => N3145, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1056);
   mult_21_C245_U1101 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1056, Z => 
                           mult_21_C245_n1359);
   mult_21_C245_U1100 : MUXB2DL port map( A0 => N3147, A1 => N3146, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1055);
   mult_21_C245_U1099 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1055, Z => 
                           mult_21_C245_n1358);
   mult_21_C245_U1098 : MUXB2DL port map( A0 => N3148, A1 => N3147, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1054);
   mult_21_C245_U1097 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1054, Z => 
                           mult_21_C245_n1357);
   mult_21_C245_U1096 : MUXB2DL port map( A0 => N3149, A1 => N3148, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1053);
   mult_21_C245_U1095 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1053, Z => 
                           mult_21_C245_n1356);
   mult_21_C245_U1094 : MUXB2DL port map( A0 => N3150, A1 => N3149, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1052);
   mult_21_C245_U1093 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1052, Z => 
                           mult_21_C245_n1355);
   mult_21_C245_U1092 : MUXB2DL port map( A0 => N3151, A1 => N3150, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1051);
   mult_21_C245_U1091 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1051, Z => 
                           mult_21_C245_n1354);
   mult_21_C245_U1090 : MUXB2DL port map( A0 => N3152, A1 => N3151, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1050);
   mult_21_C245_U1089 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1050, Z => 
                           mult_21_C245_n1353);
   mult_21_C245_U1088 : MUXB2DL port map( A0 => N3153, A1 => N3152, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1049);
   mult_21_C245_U1087 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1049, Z => 
                           mult_21_C245_n1352);
   mult_21_C245_U1086 : MUXB2DL port map( A0 => N3154, A1 => N3153, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1048);
   mult_21_C245_U1085 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1048, Z => 
                           mult_21_C245_n1351);
   mult_21_C245_U1084 : MUXB2DL port map( A0 => N3155, A1 => N3154, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1047);
   mult_21_C245_U1083 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1047, Z => 
                           mult_21_C245_n1350);
   mult_21_C245_U1082 : MUXB2DL port map( A0 => N3156, A1 => N3155, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1046);
   mult_21_C245_U1081 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1046, Z => 
                           mult_21_C245_n1349);
   mult_21_C245_U1080 : MUXB2DL port map( A0 => N3157, A1 => N3156, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1045);
   mult_21_C245_U1079 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1045, Z => 
                           mult_21_C245_n1348);
   mult_21_C245_U1078 : MUXB2DL port map( A0 => N3158, A1 => N3157, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1044);
   mult_21_C245_U1077 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1044, Z => 
                           mult_21_C245_n1347);
   mult_21_C245_U1076 : MUXB2DL port map( A0 => N3159, A1 => N3158, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1043);
   mult_21_C245_U1075 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1043, Z => 
                           mult_21_C245_n1346);
   mult_21_C245_U1074 : MUXB2DL port map( A0 => N3160, A1 => N3159, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1042);
   mult_21_C245_U1073 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1042, Z => 
                           mult_21_C245_n1345);
   mult_21_C245_U1072 : MUXB2DL port map( A0 => N3161, A1 => N3160, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1041);
   mult_21_C245_U1071 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1041, Z => 
                           mult_21_C245_n1344);
   mult_21_C245_U1070 : MUXB2DL port map( A0 => N3162, A1 => N3161, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1040);
   mult_21_C245_U1069 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1040, Z => 
                           mult_21_C245_n1343);
   mult_21_C245_U1068 : MUXB2DL port map( A0 => N3163, A1 => N3162, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1039);
   mult_21_C245_U1067 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1039, Z => 
                           mult_21_C245_n1342);
   mult_21_C245_U1066 : MUXB2DL port map( A0 => N3164, A1 => N3163, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1038);
   mult_21_C245_U1065 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1038, Z => 
                           mult_21_C245_n1341);
   mult_21_C245_U1064 : MUXB2DL port map( A0 => N3165, A1 => N3164, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1037);
   mult_21_C245_U1063 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1037, Z => 
                           mult_21_C245_n1340);
   mult_21_C245_U1062 : MUXB2DL port map( A0 => N3166, A1 => N3165, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1036);
   mult_21_C245_U1061 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1036, Z => 
                           mult_21_C245_n1339);
   mult_21_C245_U1060 : MUXB2DL port map( A0 => N3167, A1 => N3166, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1035);
   mult_21_C245_U1059 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1035, Z => 
                           mult_21_C245_n1338);
   mult_21_C245_U1058 : MUXB2DL port map( A0 => N3168, A1 => N3167, SL => 
                           mult_21_C245_n8, Z => mult_21_C245_n1034);
   mult_21_C245_U1057 : MUXB2DL port map( A0 => mult_21_C245_n3, A1 => 
                           mult_21_C245_n6, SL => mult_21_C245_n1034, Z => 
                           mult_21_C245_n1337);
   mult_21_C245_U1056 : NOR2M1D1 port map( A1 => mult_21_C245_n3, A2 => 
                           mult_21_C245_n6, Z => mult_21_C245_n1096);
   mult_21_C245_U1055 : NAN2M1D1 port map( A1 => mult_21_C245_n1542, A2 => 
                           N3137, Z => mult_21_C245_n1033);
   mult_21_C245_U1054 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1033, Z => 
                           mult_21_C245_n1336);
   mult_21_C245_U1053 : MUXB2DL port map( A0 => N3138, A1 => mult_21_C245_n1543
                           , SL => mult_21_C245_n1542, Z => mult_21_C245_n1032)
                           ;
   mult_21_C245_U1052 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1032, Z => 
                           mult_21_C245_n1335);
   mult_21_C245_U1051 : MUXB2DL port map( A0 => N3139, A1 => N3138, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1031);
   mult_21_C245_U1050 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1031, Z => 
                           mult_21_C245_n1334);
   mult_21_C245_U1049 : MUXB2DL port map( A0 => N3140, A1 => N3139, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1030);
   mult_21_C245_U1048 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1030, Z => 
                           mult_21_C245_n1333);
   mult_21_C245_U1047 : MUXB2DL port map( A0 => N3141, A1 => N3140, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1029);
   mult_21_C245_U1046 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1029, Z => 
                           mult_21_C245_n1332);
   mult_21_C245_U1045 : MUXB2DL port map( A0 => N3142, A1 => N3141, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1028);
   mult_21_C245_U1044 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1028, Z => 
                           mult_21_C245_n1331);
   mult_21_C245_U1043 : MUXB2DL port map( A0 => N3143, A1 => N3142, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1027);
   mult_21_C245_U1042 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1027, Z => 
                           mult_21_C245_n1330);
   mult_21_C245_U1041 : MUXB2DL port map( A0 => N3144, A1 => N3143, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1026);
   mult_21_C245_U1040 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1026, Z => 
                           mult_21_C245_n1329);
   mult_21_C245_U1039 : MUXB2DL port map( A0 => N3145, A1 => N3144, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1025);
   mult_21_C245_U1038 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1025, Z => 
                           mult_21_C245_n1328);
   mult_21_C245_U1037 : MUXB2DL port map( A0 => N3146, A1 => N3145, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1024);
   mult_21_C245_U1036 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1024, Z => 
                           mult_21_C245_n1327);
   mult_21_C245_U1035 : MUXB2DL port map( A0 => N3147, A1 => N3146, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1023);
   mult_21_C245_U1034 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1023, Z => 
                           mult_21_C245_n1326);
   mult_21_C245_U1033 : MUXB2DL port map( A0 => N3148, A1 => N3147, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1022);
   mult_21_C245_U1032 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1022, Z => 
                           mult_21_C245_n1325);
   mult_21_C245_U1031 : MUXB2DL port map( A0 => N3149, A1 => N3148, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1021);
   mult_21_C245_U1030 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1021, Z => 
                           mult_21_C245_n1324);
   mult_21_C245_U1029 : MUXB2DL port map( A0 => N3150, A1 => N3149, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1020);
   mult_21_C245_U1028 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1020, Z => 
                           mult_21_C245_n1323);
   mult_21_C245_U1027 : MUXB2DL port map( A0 => N3151, A1 => N3150, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1019);
   mult_21_C245_U1026 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1019, Z => 
                           mult_21_C245_n1322);
   mult_21_C245_U1025 : MUXB2DL port map( A0 => N3152, A1 => N3151, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1018);
   mult_21_C245_U1024 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1018, Z => 
                           mult_21_C245_n1321);
   mult_21_C245_U1023 : MUXB2DL port map( A0 => N3153, A1 => N3152, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1017);
   mult_21_C245_U1022 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1017, Z => 
                           mult_21_C245_n1320);
   mult_21_C245_U1021 : MUXB2DL port map( A0 => N3154, A1 => N3153, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1016);
   mult_21_C245_U1020 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1016, Z => 
                           mult_21_C245_n1319);
   mult_21_C245_U1019 : MUXB2DL port map( A0 => N3155, A1 => N3154, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1015);
   mult_21_C245_U1018 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1015, Z => 
                           mult_21_C245_n1318);
   mult_21_C245_U1017 : MUXB2DL port map( A0 => N3156, A1 => N3155, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1014);
   mult_21_C245_U1016 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1014, Z => 
                           mult_21_C245_n1317);
   mult_21_C245_U1015 : MUXB2DL port map( A0 => N3157, A1 => N3156, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1013);
   mult_21_C245_U1014 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1013, Z => 
                           mult_21_C245_n1316);
   mult_21_C245_U1013 : MUXB2DL port map( A0 => N3158, A1 => N3157, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1012);
   mult_21_C245_U1012 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1012, Z => 
                           mult_21_C245_n1315);
   mult_21_C245_U1011 : MUXB2DL port map( A0 => N3159, A1 => N3158, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1011);
   mult_21_C245_U1010 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1011, Z => 
                           mult_21_C245_n1314);
   mult_21_C245_U1009 : MUXB2DL port map( A0 => N3160, A1 => N3159, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1010);
   mult_21_C245_U1008 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1010, Z => 
                           mult_21_C245_n1313);
   mult_21_C245_U1007 : MUXB2DL port map( A0 => N3161, A1 => N3160, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1009);
   mult_21_C245_U1006 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1009, Z => 
                           mult_21_C245_n1312);
   mult_21_C245_U1005 : MUXB2DL port map( A0 => N3162, A1 => N3161, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1008);
   mult_21_C245_U1004 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1008, Z => 
                           mult_21_C245_n1311);
   mult_21_C245_U1003 : MUXB2DL port map( A0 => N3163, A1 => N3162, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1007);
   mult_21_C245_U1002 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1007, Z => 
                           mult_21_C245_n1310);
   mult_21_C245_U1001 : MUXB2DL port map( A0 => N3164, A1 => N3163, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1006);
   mult_21_C245_U1000 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1006, Z => 
                           mult_21_C245_n1309);
   mult_21_C245_U999 : MUXB2DL port map( A0 => N3165, A1 => N3164, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1005);
   mult_21_C245_U998 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1005, Z => 
                           mult_21_C245_n1308);
   mult_21_C245_U997 : MUXB2DL port map( A0 => N3166, A1 => N3165, SL => 
                           mult_21_C245_n1542, Z => mult_21_C245_n1004);
   mult_21_C245_U996 : MUXB2DL port map( A0 => mult_21_C245_n1517, A1 => 
                           mult_21_C245_n14, SL => mult_21_C245_n1004, Z => 
                           mult_21_C245_n1307);
   mult_21_C245_U995 : NOR2M1D1 port map( A1 => mult_21_C245_n1517, A2 => 
                           mult_21_C245_n14, Z => mult_21_C245_n1095);
   mult_21_C245_U994 : NAN2M1D1 port map( A1 => mult_21_C245_n1541, A2 => N3137
                           , Z => mult_21_C245_n1003);
   mult_21_C245_U993 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n1003, Z => 
                           mult_21_C245_n1306);
   mult_21_C245_U992 : MUXB2DL port map( A0 => N3138, A1 => mult_21_C245_n1543,
                           SL => mult_21_C245_n1541, Z => mult_21_C245_n1002);
   mult_21_C245_U991 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n1002, Z => 
                           mult_21_C245_n1305);
   mult_21_C245_U990 : MUXB2DL port map( A0 => N3139, A1 => N3138, SL => 
                           mult_21_C245_n1541, Z => mult_21_C245_n1001);
   mult_21_C245_U989 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n1001, Z => 
                           mult_21_C245_n1304);
   mult_21_C245_U988 : MUXB2DL port map( A0 => N3140, A1 => N3139, SL => 
                           mult_21_C245_n1541, Z => mult_21_C245_n1000);
   mult_21_C245_U987 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n1000, Z => 
                           mult_21_C245_n1303);
   mult_21_C245_U986 : MUXB2DL port map( A0 => N3141, A1 => N3140, SL => 
                           mult_21_C245_n1541, Z => mult_21_C245_n999);
   mult_21_C245_U985 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n999, Z => 
                           mult_21_C245_n1302);
   mult_21_C245_U984 : MUXB2DL port map( A0 => N3142, A1 => N3141, SL => 
                           mult_21_C245_n1541, Z => mult_21_C245_n998);
   mult_21_C245_U983 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n998, Z => 
                           mult_21_C245_n1301);
   mult_21_C245_U982 : MUXB2DL port map( A0 => N3143, A1 => N3142, SL => 
                           mult_21_C245_n1541, Z => mult_21_C245_n997);
   mult_21_C245_U981 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n997, Z => 
                           mult_21_C245_n1300);
   mult_21_C245_U980 : MUXB2DL port map( A0 => N3144, A1 => N3143, SL => 
                           mult_21_C245_n1541, Z => mult_21_C245_n996);
   mult_21_C245_U979 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n996, Z => 
                           mult_21_C245_n1299);
   mult_21_C245_U978 : MUXB2DL port map( A0 => N3145, A1 => N3144, SL => 
                           mult_21_C245_n1541, Z => mult_21_C245_n995);
   mult_21_C245_U977 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n995, Z => 
                           mult_21_C245_n1298);
   mult_21_C245_U976 : MUXB2DL port map( A0 => N3146, A1 => N3145, SL => 
                           mult_21_C245_n1541, Z => mult_21_C245_n994);
   mult_21_C245_U975 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n994, Z => 
                           mult_21_C245_n1297);
   mult_21_C245_U974 : MUXB2DL port map( A0 => N3147, A1 => N3146, SL => 
                           mult_21_C245_n1541, Z => mult_21_C245_n993);
   mult_21_C245_U973 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n993, Z => 
                           mult_21_C245_n1296);
   mult_21_C245_U972 : MUXB2DL port map( A0 => N3148, A1 => N3147, SL => 
                           mult_21_C245_n1541, Z => mult_21_C245_n992);
   mult_21_C245_U971 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n992, Z => 
                           mult_21_C245_n1295);
   mult_21_C245_U970 : MUXB2DL port map( A0 => N3149, A1 => N3148, SL => 
                           mult_21_C245_n1541, Z => mult_21_C245_n991);
   mult_21_C245_U969 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n991, Z => 
                           mult_21_C245_n1294);
   mult_21_C245_U968 : MUXB2DL port map( A0 => N3150, A1 => N3149, SL => 
                           mult_21_C245_n1541, Z => mult_21_C245_n990);
   mult_21_C245_U967 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n990, Z => 
                           mult_21_C245_n1293);
   mult_21_C245_U966 : MUXB2DL port map( A0 => N3151, A1 => N3150, SL => 
                           mult_21_C245_n1541, Z => mult_21_C245_n989);
   mult_21_C245_U965 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n989, Z => 
                           mult_21_C245_n1292);
   mult_21_C245_U964 : MUXB2DL port map( A0 => N3152, A1 => N3151, SL => 
                           mult_21_C245_n1541, Z => mult_21_C245_n988);
   mult_21_C245_U963 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n988, Z => 
                           mult_21_C245_n1291);
   mult_21_C245_U962 : MUXB2DL port map( A0 => N3153, A1 => N3152, SL => 
                           mult_21_C245_n1541, Z => mult_21_C245_n987);
   mult_21_C245_U961 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n987, Z => 
                           mult_21_C245_n1290);
   mult_21_C245_U960 : MUXB2DL port map( A0 => N3154, A1 => N3153, SL => 
                           mult_21_C245_n1541, Z => mult_21_C245_n986);
   mult_21_C245_U959 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n986, Z => 
                           mult_21_C245_n1289);
   mult_21_C245_U958 : MUXB2DL port map( A0 => N3155, A1 => N3154, SL => 
                           mult_21_C245_n1541, Z => mult_21_C245_n985);
   mult_21_C245_U957 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n985, Z => 
                           mult_21_C245_n1288);
   mult_21_C245_U956 : MUXB2DL port map( A0 => N3156, A1 => N3155, SL => 
                           mult_21_C245_n1541, Z => mult_21_C245_n984);
   mult_21_C245_U955 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n984, Z => 
                           mult_21_C245_n1287);
   mult_21_C245_U954 : MUXB2DL port map( A0 => N3157, A1 => N3156, SL => 
                           mult_21_C245_n1541, Z => mult_21_C245_n983);
   mult_21_C245_U953 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n983, Z => 
                           mult_21_C245_n1286);
   mult_21_C245_U952 : MUXB2DL port map( A0 => N3158, A1 => N3157, SL => 
                           mult_21_C245_n1541, Z => mult_21_C245_n982);
   mult_21_C245_U951 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n982, Z => 
                           mult_21_C245_n1285);
   mult_21_C245_U950 : MUXB2DL port map( A0 => N3159, A1 => N3158, SL => 
                           mult_21_C245_n1541, Z => mult_21_C245_n981);
   mult_21_C245_U949 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n981, Z => 
                           mult_21_C245_n1284);
   mult_21_C245_U948 : MUXB2DL port map( A0 => N3160, A1 => N3159, SL => 
                           mult_21_C245_n1541, Z => mult_21_C245_n980);
   mult_21_C245_U947 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n980, Z => 
                           mult_21_C245_n1283);
   mult_21_C245_U946 : MUXB2DL port map( A0 => N3161, A1 => N3160, SL => 
                           mult_21_C245_n1541, Z => mult_21_C245_n979);
   mult_21_C245_U945 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n979, Z => 
                           mult_21_C245_n1282);
   mult_21_C245_U944 : MUXB2DL port map( A0 => N3162, A1 => N3161, SL => 
                           mult_21_C245_n1541, Z => mult_21_C245_n978);
   mult_21_C245_U943 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n978, Z => 
                           mult_21_C245_n1281);
   mult_21_C245_U942 : MUXB2DL port map( A0 => N3163, A1 => N3162, SL => 
                           mult_21_C245_n1541, Z => mult_21_C245_n977);
   mult_21_C245_U941 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n977, Z => 
                           mult_21_C245_n1280);
   mult_21_C245_U940 : MUXB2DL port map( A0 => N3164, A1 => N3163, SL => 
                           mult_21_C245_n1541, Z => mult_21_C245_n976);
   mult_21_C245_U939 : MUXB2DL port map( A0 => mult_21_C245_n1518, A1 => 
                           mult_21_C245_n22, SL => mult_21_C245_n976, Z => 
                           mult_21_C245_n1279);
   mult_21_C245_U938 : NOR2M1D1 port map( A1 => mult_21_C245_n1518, A2 => 
                           mult_21_C245_n22, Z => mult_21_C245_n1094);
   mult_21_C245_U937 : NAN2M1D1 port map( A1 => mult_21_C245_n1539, A2 => N3137
                           , Z => mult_21_C245_n975);
   mult_21_C245_U936 : MUXB2DL port map( A0 => mult_21_C245_n1540, A1 => 
                           mult_21_C245_n30, SL => mult_21_C245_n975, Z => 
                           mult_21_C245_n1278);
   mult_21_C245_U935 : MUXB2DL port map( A0 => N3138, A1 => N3137, SL => 
                           mult_21_C245_n1539, Z => mult_21_C245_n974);
   mult_21_C245_U934 : MUXB2DL port map( A0 => mult_21_C245_n1540, A1 => 
                           mult_21_C245_n30, SL => mult_21_C245_n974, Z => 
                           mult_21_C245_n1277);
   mult_21_C245_U933 : MUXB2DL port map( A0 => N3139, A1 => N3138, SL => 
                           mult_21_C245_n1539, Z => mult_21_C245_n973);
   mult_21_C245_U932 : MUXB2DL port map( A0 => mult_21_C245_n1540, A1 => 
                           mult_21_C245_n30, SL => mult_21_C245_n973, Z => 
                           mult_21_C245_n1276);
   mult_21_C245_U931 : MUXB2DL port map( A0 => N3140, A1 => N3139, SL => 
                           mult_21_C245_n1539, Z => mult_21_C245_n972);
   mult_21_C245_U930 : MUXB2DL port map( A0 => mult_21_C245_n1540, A1 => 
                           mult_21_C245_n30, SL => mult_21_C245_n972, Z => 
                           mult_21_C245_n1275);
   mult_21_C245_U929 : MUXB2DL port map( A0 => N3141, A1 => N3140, SL => 
                           mult_21_C245_n1539, Z => mult_21_C245_n971);
   mult_21_C245_U928 : MUXB2DL port map( A0 => mult_21_C245_n1540, A1 => 
                           mult_21_C245_n30, SL => mult_21_C245_n971, Z => 
                           mult_21_C245_n1274);
   mult_21_C245_U927 : MUXB2DL port map( A0 => N3142, A1 => N3141, SL => 
                           mult_21_C245_n1539, Z => mult_21_C245_n970);
   mult_21_C245_U926 : MUXB2DL port map( A0 => mult_21_C245_n1540, A1 => 
                           mult_21_C245_n30, SL => mult_21_C245_n970, Z => 
                           mult_21_C245_n1273);
   mult_21_C245_U925 : MUXB2DL port map( A0 => N3143, A1 => N3142, SL => 
                           mult_21_C245_n1539, Z => mult_21_C245_n969);
   mult_21_C245_U924 : MUXB2DL port map( A0 => mult_21_C245_n1540, A1 => 
                           mult_21_C245_n30, SL => mult_21_C245_n969, Z => 
                           mult_21_C245_n1272);
   mult_21_C245_U923 : MUXB2DL port map( A0 => N3144, A1 => N3143, SL => 
                           mult_21_C245_n1539, Z => mult_21_C245_n968);
   mult_21_C245_U922 : MUXB2DL port map( A0 => mult_21_C245_n1540, A1 => 
                           mult_21_C245_n30, SL => mult_21_C245_n968, Z => 
                           mult_21_C245_n1271);
   mult_21_C245_U921 : MUXB2DL port map( A0 => N3145, A1 => N3144, SL => 
                           mult_21_C245_n1539, Z => mult_21_C245_n967);
   mult_21_C245_U920 : MUXB2DL port map( A0 => mult_21_C245_n1540, A1 => 
                           mult_21_C245_n30, SL => mult_21_C245_n967, Z => 
                           mult_21_C245_n1270);
   mult_21_C245_U919 : MUXB2DL port map( A0 => N3146, A1 => N3145, SL => 
                           mult_21_C245_n1539, Z => mult_21_C245_n966);
   mult_21_C245_U918 : MUXB2DL port map( A0 => mult_21_C245_n1540, A1 => 
                           mult_21_C245_n30, SL => mult_21_C245_n966, Z => 
                           mult_21_C245_n1269);
   mult_21_C245_U917 : MUXB2DL port map( A0 => N3147, A1 => N3146, SL => 
                           mult_21_C245_n1539, Z => mult_21_C245_n965);
   mult_21_C245_U916 : MUXB2DL port map( A0 => mult_21_C245_n1540, A1 => 
                           mult_21_C245_n30, SL => mult_21_C245_n965, Z => 
                           mult_21_C245_n1268);
   mult_21_C245_U915 : MUXB2DL port map( A0 => N3148, A1 => N3147, SL => 
                           mult_21_C245_n1539, Z => mult_21_C245_n964);
   mult_21_C245_U914 : MUXB2DL port map( A0 => mult_21_C245_n1540, A1 => 
                           mult_21_C245_n30, SL => mult_21_C245_n964, Z => 
                           mult_21_C245_n1267);
   mult_21_C245_U913 : MUXB2DL port map( A0 => N3149, A1 => N3148, SL => 
                           mult_21_C245_n1539, Z => mult_21_C245_n963);
   mult_21_C245_U912 : MUXB2DL port map( A0 => mult_21_C245_n1540, A1 => 
                           mult_21_C245_n30, SL => mult_21_C245_n963, Z => 
                           mult_21_C245_n1266);
   mult_21_C245_U911 : MUXB2DL port map( A0 => N3150, A1 => N3149, SL => 
                           mult_21_C245_n1539, Z => mult_21_C245_n962);
   mult_21_C245_U910 : MUXB2DL port map( A0 => mult_21_C245_n1540, A1 => 
                           mult_21_C245_n30, SL => mult_21_C245_n962, Z => 
                           mult_21_C245_n1265);
   mult_21_C245_U909 : MUXB2DL port map( A0 => N3151, A1 => N3150, SL => 
                           mult_21_C245_n1539, Z => mult_21_C245_n961);
   mult_21_C245_U908 : MUXB2DL port map( A0 => mult_21_C245_n1540, A1 => 
                           mult_21_C245_n30, SL => mult_21_C245_n961, Z => 
                           mult_21_C245_n1264);
   mult_21_C245_U907 : MUXB2DL port map( A0 => N3152, A1 => N3151, SL => 
                           mult_21_C245_n1539, Z => mult_21_C245_n960);
   mult_21_C245_U906 : MUXB2DL port map( A0 => mult_21_C245_n1540, A1 => 
                           mult_21_C245_n30, SL => mult_21_C245_n960, Z => 
                           mult_21_C245_n1263);
   mult_21_C245_U905 : MUXB2DL port map( A0 => N3153, A1 => N3152, SL => 
                           mult_21_C245_n1539, Z => mult_21_C245_n959);
   mult_21_C245_U904 : MUXB2DL port map( A0 => mult_21_C245_n1540, A1 => 
                           mult_21_C245_n30, SL => mult_21_C245_n959, Z => 
                           mult_21_C245_n1262);
   mult_21_C245_U903 : MUXB2DL port map( A0 => N3154, A1 => N3153, SL => 
                           mult_21_C245_n1539, Z => mult_21_C245_n958);
   mult_21_C245_U902 : MUXB2DL port map( A0 => mult_21_C245_n1540, A1 => 
                           mult_21_C245_n30, SL => mult_21_C245_n958, Z => 
                           mult_21_C245_n1261);
   mult_21_C245_U901 : MUXB2DL port map( A0 => N3155, A1 => N3154, SL => 
                           mult_21_C245_n1539, Z => mult_21_C245_n957);
   mult_21_C245_U900 : MUXB2DL port map( A0 => mult_21_C245_n1540, A1 => 
                           mult_21_C245_n30, SL => mult_21_C245_n957, Z => 
                           mult_21_C245_n1260);
   mult_21_C245_U899 : MUXB2DL port map( A0 => N3156, A1 => N3155, SL => 
                           mult_21_C245_n1539, Z => mult_21_C245_n956);
   mult_21_C245_U898 : MUXB2DL port map( A0 => mult_21_C245_n1540, A1 => 
                           mult_21_C245_n30, SL => mult_21_C245_n956, Z => 
                           mult_21_C245_n1259);
   mult_21_C245_U897 : MUXB2DL port map( A0 => N3157, A1 => N3156, SL => 
                           mult_21_C245_n1539, Z => mult_21_C245_n955);
   mult_21_C245_U896 : MUXB2DL port map( A0 => mult_21_C245_n1540, A1 => 
                           mult_21_C245_n30, SL => mult_21_C245_n955, Z => 
                           mult_21_C245_n1258);
   mult_21_C245_U895 : MUXB2DL port map( A0 => N3158, A1 => N3157, SL => 
                           mult_21_C245_n1539, Z => mult_21_C245_n954);
   mult_21_C245_U894 : MUXB2DL port map( A0 => mult_21_C245_n1540, A1 => 
                           mult_21_C245_n30, SL => mult_21_C245_n954, Z => 
                           mult_21_C245_n1257);
   mult_21_C245_U893 : MUXB2DL port map( A0 => N3159, A1 => N3158, SL => 
                           mult_21_C245_n1539, Z => mult_21_C245_n953);
   mult_21_C245_U892 : MUXB2DL port map( A0 => mult_21_C245_n1540, A1 => 
                           mult_21_C245_n30, SL => mult_21_C245_n953, Z => 
                           mult_21_C245_n1256);
   mult_21_C245_U891 : MUXB2DL port map( A0 => N3160, A1 => N3159, SL => 
                           mult_21_C245_n1539, Z => mult_21_C245_n952);
   mult_21_C245_U890 : MUXB2DL port map( A0 => mult_21_C245_n1540, A1 => 
                           mult_21_C245_n30, SL => mult_21_C245_n952, Z => 
                           mult_21_C245_n1255);
   mult_21_C245_U889 : MUXB2DL port map( A0 => N3161, A1 => N3160, SL => 
                           mult_21_C245_n1539, Z => mult_21_C245_n951);
   mult_21_C245_U888 : MUXB2DL port map( A0 => mult_21_C245_n1540, A1 => 
                           mult_21_C245_n30, SL => mult_21_C245_n951, Z => 
                           mult_21_C245_n1254);
   mult_21_C245_U887 : MUXB2DL port map( A0 => N3162, A1 => N3161, SL => 
                           mult_21_C245_n1539, Z => mult_21_C245_n950);
   mult_21_C245_U886 : MUXB2DL port map( A0 => mult_21_C245_n1540, A1 => 
                           mult_21_C245_n30, SL => mult_21_C245_n950, Z => 
                           mult_21_C245_n1253);
   mult_21_C245_U884 : NAN2M1D1 port map( A1 => mult_21_C245_n1538, A2 => N3137
                           , Z => mult_21_C245_n949);
   mult_21_C245_U883 : MUXB2DL port map( A0 => mult_21_C245_n1519, A1 => 
                           mult_21_C245_n38, SL => mult_21_C245_n949, Z => 
                           mult_21_C245_n1252);
   mult_21_C245_U882 : MUXB2DL port map( A0 => N3138, A1 => N3137, SL => 
                           mult_21_C245_n1538, Z => mult_21_C245_n948);
   mult_21_C245_U881 : MUXB2DL port map( A0 => mult_21_C245_n1519, A1 => 
                           mult_21_C245_n38, SL => mult_21_C245_n948, Z => 
                           mult_21_C245_n1251);
   mult_21_C245_U880 : MUXB2DL port map( A0 => N3139, A1 => N3138, SL => 
                           mult_21_C245_n1538, Z => mult_21_C245_n947);
   mult_21_C245_U879 : MUXB2DL port map( A0 => mult_21_C245_n1519, A1 => 
                           mult_21_C245_n38, SL => mult_21_C245_n947, Z => 
                           mult_21_C245_n1250);
   mult_21_C245_U878 : MUXB2DL port map( A0 => N3140, A1 => N3139, SL => 
                           mult_21_C245_n1538, Z => mult_21_C245_n946);
   mult_21_C245_U877 : MUXB2DL port map( A0 => mult_21_C245_n1519, A1 => 
                           mult_21_C245_n38, SL => mult_21_C245_n946, Z => 
                           mult_21_C245_n1249);
   mult_21_C245_U876 : MUXB2DL port map( A0 => N3141, A1 => N3140, SL => 
                           mult_21_C245_n1538, Z => mult_21_C245_n945);
   mult_21_C245_U875 : MUXB2DL port map( A0 => mult_21_C245_n1519, A1 => 
                           mult_21_C245_n38, SL => mult_21_C245_n945, Z => 
                           mult_21_C245_n1248);
   mult_21_C245_U874 : MUXB2DL port map( A0 => N3142, A1 => N3141, SL => 
                           mult_21_C245_n1538, Z => mult_21_C245_n944);
   mult_21_C245_U873 : MUXB2DL port map( A0 => mult_21_C245_n1519, A1 => 
                           mult_21_C245_n38, SL => mult_21_C245_n944, Z => 
                           mult_21_C245_n1247);
   mult_21_C245_U872 : MUXB2DL port map( A0 => N3143, A1 => N3142, SL => 
                           mult_21_C245_n1538, Z => mult_21_C245_n943);
   mult_21_C245_U871 : MUXB2DL port map( A0 => mult_21_C245_n1519, A1 => 
                           mult_21_C245_n38, SL => mult_21_C245_n943, Z => 
                           mult_21_C245_n1246);
   mult_21_C245_U870 : MUXB2DL port map( A0 => N3144, A1 => N3143, SL => 
                           mult_21_C245_n1538, Z => mult_21_C245_n942);
   mult_21_C245_U869 : MUXB2DL port map( A0 => mult_21_C245_n1519, A1 => 
                           mult_21_C245_n38, SL => mult_21_C245_n942, Z => 
                           mult_21_C245_n1245);
   mult_21_C245_U868 : MUXB2DL port map( A0 => N3145, A1 => N3144, SL => 
                           mult_21_C245_n1538, Z => mult_21_C245_n941);
   mult_21_C245_U867 : MUXB2DL port map( A0 => mult_21_C245_n1519, A1 => 
                           mult_21_C245_n38, SL => mult_21_C245_n941, Z => 
                           mult_21_C245_n1244);
   mult_21_C245_U866 : MUXB2DL port map( A0 => N3146, A1 => N3145, SL => 
                           mult_21_C245_n1538, Z => mult_21_C245_n940);
   mult_21_C245_U865 : MUXB2DL port map( A0 => mult_21_C245_n1519, A1 => 
                           mult_21_C245_n38, SL => mult_21_C245_n940, Z => 
                           mult_21_C245_n1243);
   mult_21_C245_U864 : MUXB2DL port map( A0 => N3147, A1 => N3146, SL => 
                           mult_21_C245_n1538, Z => mult_21_C245_n939);
   mult_21_C245_U863 : MUXB2DL port map( A0 => mult_21_C245_n1519, A1 => 
                           mult_21_C245_n38, SL => mult_21_C245_n939, Z => 
                           mult_21_C245_n1242);
   mult_21_C245_U862 : MUXB2DL port map( A0 => N3148, A1 => N3147, SL => 
                           mult_21_C245_n1538, Z => mult_21_C245_n938);
   mult_21_C245_U861 : MUXB2DL port map( A0 => mult_21_C245_n1519, A1 => 
                           mult_21_C245_n38, SL => mult_21_C245_n938, Z => 
                           mult_21_C245_n1241);
   mult_21_C245_U860 : MUXB2DL port map( A0 => N3149, A1 => N3148, SL => 
                           mult_21_C245_n1538, Z => mult_21_C245_n937);
   mult_21_C245_U859 : MUXB2DL port map( A0 => mult_21_C245_n1519, A1 => 
                           mult_21_C245_n38, SL => mult_21_C245_n937, Z => 
                           mult_21_C245_n1240);
   mult_21_C245_U858 : MUXB2DL port map( A0 => N3150, A1 => N3149, SL => 
                           mult_21_C245_n1538, Z => mult_21_C245_n936);
   mult_21_C245_U857 : MUXB2DL port map( A0 => mult_21_C245_n1519, A1 => 
                           mult_21_C245_n38, SL => mult_21_C245_n936, Z => 
                           mult_21_C245_n1239);
   mult_21_C245_U856 : MUXB2DL port map( A0 => N3151, A1 => N3150, SL => 
                           mult_21_C245_n1538, Z => mult_21_C245_n935);
   mult_21_C245_U855 : MUXB2DL port map( A0 => mult_21_C245_n1519, A1 => 
                           mult_21_C245_n38, SL => mult_21_C245_n935, Z => 
                           mult_21_C245_n1238);
   mult_21_C245_U854 : MUXB2DL port map( A0 => N3152, A1 => N3151, SL => 
                           mult_21_C245_n1538, Z => mult_21_C245_n934);
   mult_21_C245_U853 : MUXB2DL port map( A0 => mult_21_C245_n1519, A1 => 
                           mult_21_C245_n38, SL => mult_21_C245_n934, Z => 
                           mult_21_C245_n1237);
   mult_21_C245_U852 : MUXB2DL port map( A0 => N3153, A1 => N3152, SL => 
                           mult_21_C245_n1538, Z => mult_21_C245_n933);
   mult_21_C245_U851 : MUXB2DL port map( A0 => mult_21_C245_n1519, A1 => 
                           mult_21_C245_n38, SL => mult_21_C245_n933, Z => 
                           mult_21_C245_n1236);
   mult_21_C245_U850 : MUXB2DL port map( A0 => N3154, A1 => N3153, SL => 
                           mult_21_C245_n1538, Z => mult_21_C245_n932);
   mult_21_C245_U849 : MUXB2DL port map( A0 => mult_21_C245_n1519, A1 => 
                           mult_21_C245_n38, SL => mult_21_C245_n932, Z => 
                           mult_21_C245_n1235);
   mult_21_C245_U848 : MUXB2DL port map( A0 => N3155, A1 => N3154, SL => 
                           mult_21_C245_n1538, Z => mult_21_C245_n931);
   mult_21_C245_U847 : MUXB2DL port map( A0 => mult_21_C245_n1519, A1 => 
                           mult_21_C245_n38, SL => mult_21_C245_n931, Z => 
                           mult_21_C245_n1234);
   mult_21_C245_U846 : MUXB2DL port map( A0 => N3156, A1 => N3155, SL => 
                           mult_21_C245_n1538, Z => mult_21_C245_n930);
   mult_21_C245_U845 : MUXB2DL port map( A0 => mult_21_C245_n1519, A1 => 
                           mult_21_C245_n38, SL => mult_21_C245_n930, Z => 
                           mult_21_C245_n1233);
   mult_21_C245_U844 : MUXB2DL port map( A0 => N3157, A1 => N3156, SL => 
                           mult_21_C245_n1538, Z => mult_21_C245_n929);
   mult_21_C245_U843 : MUXB2DL port map( A0 => mult_21_C245_n1519, A1 => 
                           mult_21_C245_n38, SL => mult_21_C245_n929, Z => 
                           mult_21_C245_n1232);
   mult_21_C245_U842 : MUXB2DL port map( A0 => N3158, A1 => N3157, SL => 
                           mult_21_C245_n1538, Z => mult_21_C245_n928);
   mult_21_C245_U841 : MUXB2DL port map( A0 => mult_21_C245_n1519, A1 => 
                           mult_21_C245_n38, SL => mult_21_C245_n928, Z => 
                           mult_21_C245_n1231);
   mult_21_C245_U840 : MUXB2DL port map( A0 => N3159, A1 => N3158, SL => 
                           mult_21_C245_n1538, Z => mult_21_C245_n927);
   mult_21_C245_U839 : MUXB2DL port map( A0 => mult_21_C245_n1519, A1 => 
                           mult_21_C245_n38, SL => mult_21_C245_n927, Z => 
                           mult_21_C245_n1230);
   mult_21_C245_U838 : MUXB2DL port map( A0 => N3160, A1 => N3159, SL => 
                           mult_21_C245_n1538, Z => mult_21_C245_n926);
   mult_21_C245_U837 : MUXB2DL port map( A0 => mult_21_C245_n1519, A1 => 
                           mult_21_C245_n38, SL => mult_21_C245_n926, Z => 
                           mult_21_C245_n1229);
   mult_21_C245_U836 : NOR2M1D1 port map( A1 => mult_21_C245_n1519, A2 => 
                           mult_21_C245_n38, Z => mult_21_C245_n1092);
   mult_21_C245_U835 : NAN2M1D1 port map( A1 => mult_21_C245_n48, A2 => N3137, 
                           Z => mult_21_C245_n925);
   mult_21_C245_U834 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n45, SL => mult_21_C245_n925, Z => 
                           mult_21_C245_n1228);
   mult_21_C245_U833 : MUXB2DL port map( A0 => N3138, A1 => N3137, SL => 
                           mult_21_C245_n48, Z => mult_21_C245_n924);
   mult_21_C245_U832 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n45, SL => mult_21_C245_n924, Z => 
                           mult_21_C245_n1227);
   mult_21_C245_U831 : MUXB2DL port map( A0 => N3139, A1 => N3138, SL => 
                           mult_21_C245_n48, Z => mult_21_C245_n923);
   mult_21_C245_U830 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n45, SL => mult_21_C245_n923, Z => 
                           mult_21_C245_n1226);
   mult_21_C245_U829 : MUXB2DL port map( A0 => N3140, A1 => N3139, SL => 
                           mult_21_C245_n48, Z => mult_21_C245_n922);
   mult_21_C245_U828 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n45, SL => mult_21_C245_n922, Z => 
                           mult_21_C245_n1225);
   mult_21_C245_U827 : MUXB2DL port map( A0 => N3141, A1 => N3140, SL => 
                           mult_21_C245_n48, Z => mult_21_C245_n921);
   mult_21_C245_U826 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n45, SL => mult_21_C245_n921, Z => 
                           mult_21_C245_n1224);
   mult_21_C245_U825 : MUXB2DL port map( A0 => N3142, A1 => N3141, SL => 
                           mult_21_C245_n48, Z => mult_21_C245_n920);
   mult_21_C245_U824 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n45, SL => mult_21_C245_n920, Z => 
                           mult_21_C245_n1223);
   mult_21_C245_U823 : MUXB2DL port map( A0 => N3143, A1 => N3142, SL => 
                           mult_21_C245_n48, Z => mult_21_C245_n919);
   mult_21_C245_U822 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n45, SL => mult_21_C245_n919, Z => 
                           mult_21_C245_n1222);
   mult_21_C245_U821 : MUXB2DL port map( A0 => N3144, A1 => N3143, SL => 
                           mult_21_C245_n48, Z => mult_21_C245_n918);
   mult_21_C245_U820 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n45, SL => mult_21_C245_n918, Z => 
                           mult_21_C245_n1221);
   mult_21_C245_U819 : MUXB2DL port map( A0 => N3145, A1 => N3144, SL => 
                           mult_21_C245_n48, Z => mult_21_C245_n917);
   mult_21_C245_U818 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n45, SL => mult_21_C245_n917, Z => 
                           mult_21_C245_n1220);
   mult_21_C245_U817 : MUXB2DL port map( A0 => N3146, A1 => N3145, SL => 
                           mult_21_C245_n48, Z => mult_21_C245_n916);
   mult_21_C245_U816 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n45, SL => mult_21_C245_n916, Z => 
                           mult_21_C245_n1219);
   mult_21_C245_U815 : MUXB2DL port map( A0 => N3147, A1 => N3146, SL => 
                           mult_21_C245_n48, Z => mult_21_C245_n915);
   mult_21_C245_U814 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n45, SL => mult_21_C245_n915, Z => 
                           mult_21_C245_n1218);
   mult_21_C245_U813 : MUXB2DL port map( A0 => N3148, A1 => N3147, SL => 
                           mult_21_C245_n48, Z => mult_21_C245_n914);
   mult_21_C245_U812 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n45, SL => mult_21_C245_n914, Z => 
                           mult_21_C245_n1217);
   mult_21_C245_U811 : MUXB2DL port map( A0 => N3149, A1 => N3148, SL => 
                           mult_21_C245_n48, Z => mult_21_C245_n913);
   mult_21_C245_U810 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n45, SL => mult_21_C245_n913, Z => 
                           mult_21_C245_n1216);
   mult_21_C245_U809 : MUXB2DL port map( A0 => N3150, A1 => N3149, SL => 
                           mult_21_C245_n48, Z => mult_21_C245_n912);
   mult_21_C245_U808 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n45, SL => mult_21_C245_n912, Z => 
                           mult_21_C245_n1215);
   mult_21_C245_U807 : MUXB2DL port map( A0 => N3151, A1 => N3150, SL => 
                           mult_21_C245_n48, Z => mult_21_C245_n911);
   mult_21_C245_U806 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n45, SL => mult_21_C245_n911, Z => 
                           mult_21_C245_n1214);
   mult_21_C245_U805 : MUXB2DL port map( A0 => N3152, A1 => N3151, SL => 
                           mult_21_C245_n48, Z => mult_21_C245_n910);
   mult_21_C245_U804 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n45, SL => mult_21_C245_n910, Z => 
                           mult_21_C245_n1213);
   mult_21_C245_U803 : MUXB2DL port map( A0 => N3153, A1 => N3152, SL => 
                           mult_21_C245_n48, Z => mult_21_C245_n909);
   mult_21_C245_U802 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n45, SL => mult_21_C245_n909, Z => 
                           mult_21_C245_n1212);
   mult_21_C245_U801 : MUXB2DL port map( A0 => N3154, A1 => N3153, SL => 
                           mult_21_C245_n48, Z => mult_21_C245_n908);
   mult_21_C245_U800 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n45, SL => mult_21_C245_n908, Z => 
                           mult_21_C245_n1211);
   mult_21_C245_U799 : MUXB2DL port map( A0 => N3155, A1 => N3154, SL => 
                           mult_21_C245_n48, Z => mult_21_C245_n907);
   mult_21_C245_U798 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n45, SL => mult_21_C245_n907, Z => 
                           mult_21_C245_n1210);
   mult_21_C245_U797 : MUXB2DL port map( A0 => N3156, A1 => N3155, SL => 
                           mult_21_C245_n48, Z => mult_21_C245_n906);
   mult_21_C245_U796 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n45, SL => mult_21_C245_n906, Z => 
                           mult_21_C245_n1209);
   mult_21_C245_U795 : MUXB2DL port map( A0 => N3157, A1 => N3156, SL => 
                           mult_21_C245_n48, Z => mult_21_C245_n905);
   mult_21_C245_U794 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n45, SL => mult_21_C245_n905, Z => 
                           mult_21_C245_n1208);
   mult_21_C245_U793 : MUXB2DL port map( A0 => N3158, A1 => N3157, SL => 
                           mult_21_C245_n48, Z => mult_21_C245_n904);
   mult_21_C245_U792 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n45, SL => mult_21_C245_n904, Z => 
                           mult_21_C245_n1207);
   mult_21_C245_U791 : NOR2M1D1 port map( A1 => mult_21_C245_n42, A2 => 
                           mult_21_C245_n45, Z => mult_21_C245_n1091);
   mult_21_C245_U790 : NAN2M1D1 port map( A1 => mult_21_C245_n56, A2 => 
                           mult_21_C245_n1543, Z => mult_21_C245_n903);
   mult_21_C245_U789 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n53, SL => mult_21_C245_n903, Z => 
                           mult_21_C245_n1206);
   mult_21_C245_U788 : MUXB2DL port map( A0 => N3138, A1 => N3137, SL => 
                           mult_21_C245_n56, Z => mult_21_C245_n902);
   mult_21_C245_U787 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n53, SL => mult_21_C245_n902, Z => 
                           mult_21_C245_n1205);
   mult_21_C245_U786 : MUXB2DL port map( A0 => N3139, A1 => N3138, SL => 
                           mult_21_C245_n56, Z => mult_21_C245_n901);
   mult_21_C245_U785 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n53, SL => mult_21_C245_n901, Z => 
                           mult_21_C245_n1204);
   mult_21_C245_U784 : MUXB2DL port map( A0 => N3140, A1 => N3139, SL => 
                           mult_21_C245_n56, Z => mult_21_C245_n900);
   mult_21_C245_U783 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n53, SL => mult_21_C245_n900, Z => 
                           mult_21_C245_n1203);
   mult_21_C245_U782 : MUXB2DL port map( A0 => N3141, A1 => N3140, SL => 
                           mult_21_C245_n56, Z => mult_21_C245_n899);
   mult_21_C245_U781 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n53, SL => mult_21_C245_n899, Z => 
                           mult_21_C245_n1202);
   mult_21_C245_U780 : MUXB2DL port map( A0 => N3142, A1 => N3141, SL => 
                           mult_21_C245_n56, Z => mult_21_C245_n898);
   mult_21_C245_U779 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n53, SL => mult_21_C245_n898, Z => 
                           mult_21_C245_n1201);
   mult_21_C245_U778 : MUXB2DL port map( A0 => N3143, A1 => N3142, SL => 
                           mult_21_C245_n56, Z => mult_21_C245_n897);
   mult_21_C245_U777 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n53, SL => mult_21_C245_n897, Z => 
                           mult_21_C245_n1200);
   mult_21_C245_U776 : MUXB2DL port map( A0 => N3144, A1 => N3143, SL => 
                           mult_21_C245_n56, Z => mult_21_C245_n896);
   mult_21_C245_U775 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n53, SL => mult_21_C245_n896, Z => 
                           mult_21_C245_n1199);
   mult_21_C245_U774 : MUXB2DL port map( A0 => N3145, A1 => N3144, SL => 
                           mult_21_C245_n56, Z => mult_21_C245_n895);
   mult_21_C245_U773 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n53, SL => mult_21_C245_n895, Z => 
                           mult_21_C245_n1198);
   mult_21_C245_U772 : MUXB2DL port map( A0 => N3146, A1 => N3145, SL => 
                           mult_21_C245_n56, Z => mult_21_C245_n894);
   mult_21_C245_U771 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n53, SL => mult_21_C245_n894, Z => 
                           mult_21_C245_n1197);
   mult_21_C245_U770 : MUXB2DL port map( A0 => N3147, A1 => N3146, SL => 
                           mult_21_C245_n56, Z => mult_21_C245_n893);
   mult_21_C245_U769 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n53, SL => mult_21_C245_n893, Z => 
                           mult_21_C245_n1196);
   mult_21_C245_U768 : MUXB2DL port map( A0 => N3148, A1 => N3147, SL => 
                           mult_21_C245_n56, Z => mult_21_C245_n892);
   mult_21_C245_U767 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n53, SL => mult_21_C245_n892, Z => 
                           mult_21_C245_n1195);
   mult_21_C245_U766 : MUXB2DL port map( A0 => N3149, A1 => N3148, SL => 
                           mult_21_C245_n56, Z => mult_21_C245_n891);
   mult_21_C245_U765 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n53, SL => mult_21_C245_n891, Z => 
                           mult_21_C245_n1194);
   mult_21_C245_U764 : MUXB2DL port map( A0 => N3150, A1 => N3149, SL => 
                           mult_21_C245_n56, Z => mult_21_C245_n890);
   mult_21_C245_U763 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n53, SL => mult_21_C245_n890, Z => 
                           mult_21_C245_n1193);
   mult_21_C245_U762 : MUXB2DL port map( A0 => N3151, A1 => N3150, SL => 
                           mult_21_C245_n56, Z => mult_21_C245_n889);
   mult_21_C245_U761 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n53, SL => mult_21_C245_n889, Z => 
                           mult_21_C245_n1192);
   mult_21_C245_U760 : MUXB2DL port map( A0 => N3152, A1 => N3151, SL => 
                           mult_21_C245_n56, Z => mult_21_C245_n888);
   mult_21_C245_U759 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n53, SL => mult_21_C245_n888, Z => 
                           mult_21_C245_n1191);
   mult_21_C245_U758 : MUXB2DL port map( A0 => N3153, A1 => N3152, SL => 
                           mult_21_C245_n56, Z => mult_21_C245_n887);
   mult_21_C245_U757 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n53, SL => mult_21_C245_n887, Z => 
                           mult_21_C245_n1190);
   mult_21_C245_U756 : MUXB2DL port map( A0 => N3154, A1 => N3153, SL => 
                           mult_21_C245_n56, Z => mult_21_C245_n886);
   mult_21_C245_U755 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n53, SL => mult_21_C245_n886, Z => 
                           mult_21_C245_n1189);
   mult_21_C245_U754 : MUXB2DL port map( A0 => N3155, A1 => N3154, SL => 
                           mult_21_C245_n56, Z => mult_21_C245_n885);
   mult_21_C245_U753 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n53, SL => mult_21_C245_n885, Z => 
                           mult_21_C245_n1188);
   mult_21_C245_U752 : MUXB2DL port map( A0 => N3156, A1 => N3155, SL => 
                           mult_21_C245_n56, Z => mult_21_C245_n884);
   mult_21_C245_U751 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n53, SL => mult_21_C245_n884, Z => 
                           mult_21_C245_n1187);
   mult_21_C245_U750 : NOR2M1D1 port map( A1 => mult_21_C245_n50, A2 => 
                           mult_21_C245_n53, Z => mult_21_C245_n1090);
   mult_21_C245_U749 : NAN2M1D1 port map( A1 => mult_21_C245_n63, A2 => N3137, 
                           Z => mult_21_C245_n883);
   mult_21_C245_U748 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n61, SL => mult_21_C245_n883, Z => 
                           mult_21_C245_n1186);
   mult_21_C245_U747 : MUXB2DL port map( A0 => N3138, A1 => mult_21_C245_n1543,
                           SL => mult_21_C245_n63, Z => mult_21_C245_n882);
   mult_21_C245_U746 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n61, SL => mult_21_C245_n882, Z => 
                           mult_21_C245_n1185);
   mult_21_C245_U745 : MUXB2DL port map( A0 => N3139, A1 => N3138, SL => 
                           mult_21_C245_n63, Z => mult_21_C245_n881);
   mult_21_C245_U744 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n61, SL => mult_21_C245_n881, Z => 
                           mult_21_C245_n1184);
   mult_21_C245_U743 : MUXB2DL port map( A0 => N3140, A1 => N3139, SL => 
                           mult_21_C245_n63, Z => mult_21_C245_n880);
   mult_21_C245_U742 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n61, SL => mult_21_C245_n880, Z => 
                           mult_21_C245_n1183);
   mult_21_C245_U741 : MUXB2DL port map( A0 => N3141, A1 => N3140, SL => 
                           mult_21_C245_n63, Z => mult_21_C245_n879);
   mult_21_C245_U740 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n61, SL => mult_21_C245_n879, Z => 
                           mult_21_C245_n1182);
   mult_21_C245_U739 : MUXB2DL port map( A0 => N3142, A1 => N3141, SL => 
                           mult_21_C245_n63, Z => mult_21_C245_n878);
   mult_21_C245_U738 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n61, SL => mult_21_C245_n878, Z => 
                           mult_21_C245_n1181);
   mult_21_C245_U737 : MUXB2DL port map( A0 => N3143, A1 => N3142, SL => 
                           mult_21_C245_n63, Z => mult_21_C245_n877);
   mult_21_C245_U736 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n61, SL => mult_21_C245_n877, Z => 
                           mult_21_C245_n1180);
   mult_21_C245_U735 : MUXB2DL port map( A0 => N3144, A1 => N3143, SL => 
                           mult_21_C245_n63, Z => mult_21_C245_n876);
   mult_21_C245_U734 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n61, SL => mult_21_C245_n876, Z => 
                           mult_21_C245_n1179);
   mult_21_C245_U733 : MUXB2DL port map( A0 => N3145, A1 => N3144, SL => 
                           mult_21_C245_n63, Z => mult_21_C245_n875);
   mult_21_C245_U732 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n61, SL => mult_21_C245_n875, Z => 
                           mult_21_C245_n1178);
   mult_21_C245_U731 : MUXB2DL port map( A0 => N3146, A1 => N3145, SL => 
                           mult_21_C245_n63, Z => mult_21_C245_n874);
   mult_21_C245_U730 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n61, SL => mult_21_C245_n874, Z => 
                           mult_21_C245_n1177);
   mult_21_C245_U729 : MUXB2DL port map( A0 => N3147, A1 => N3146, SL => 
                           mult_21_C245_n63, Z => mult_21_C245_n873);
   mult_21_C245_U728 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n61, SL => mult_21_C245_n873, Z => 
                           mult_21_C245_n1176);
   mult_21_C245_U727 : MUXB2DL port map( A0 => N3148, A1 => N3147, SL => 
                           mult_21_C245_n63, Z => mult_21_C245_n872);
   mult_21_C245_U726 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n61, SL => mult_21_C245_n872, Z => 
                           mult_21_C245_n1175);
   mult_21_C245_U725 : MUXB2DL port map( A0 => N3149, A1 => N3148, SL => 
                           mult_21_C245_n63, Z => mult_21_C245_n871);
   mult_21_C245_U724 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n61, SL => mult_21_C245_n871, Z => 
                           mult_21_C245_n1174);
   mult_21_C245_U723 : MUXB2DL port map( A0 => N3150, A1 => N3149, SL => 
                           mult_21_C245_n63, Z => mult_21_C245_n870);
   mult_21_C245_U722 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n61, SL => mult_21_C245_n870, Z => 
                           mult_21_C245_n1173);
   mult_21_C245_U721 : MUXB2DL port map( A0 => N3151, A1 => N3150, SL => 
                           mult_21_C245_n63, Z => mult_21_C245_n869);
   mult_21_C245_U720 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n61, SL => mult_21_C245_n869, Z => 
                           mult_21_C245_n1172);
   mult_21_C245_U719 : MUXB2DL port map( A0 => N3152, A1 => N3151, SL => 
                           mult_21_C245_n63, Z => mult_21_C245_n868);
   mult_21_C245_U718 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n61, SL => mult_21_C245_n868, Z => 
                           mult_21_C245_n1171);
   mult_21_C245_U717 : MUXB2DL port map( A0 => N3153, A1 => N3152, SL => 
                           mult_21_C245_n63, Z => mult_21_C245_n867);
   mult_21_C245_U716 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n61, SL => mult_21_C245_n867, Z => 
                           mult_21_C245_n1170);
   mult_21_C245_U715 : MUXB2DL port map( A0 => N3154, A1 => N3153, SL => 
                           mult_21_C245_n63, Z => mult_21_C245_n866);
   mult_21_C245_U714 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n61, SL => mult_21_C245_n866, Z => 
                           mult_21_C245_n1169);
   mult_21_C245_U713 : NOR2M1D1 port map( A1 => mult_21_C245_n58, A2 => 
                           mult_21_C245_n61, Z => mult_21_C245_n1089);
   mult_21_C245_U712 : NAN2M1D1 port map( A1 => mult_21_C245_n71, A2 => N3137, 
                           Z => mult_21_C245_n865);
   mult_21_C245_U711 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n69, SL => mult_21_C245_n865, Z => 
                           mult_21_C245_n1168);
   mult_21_C245_U710 : MUXB2DL port map( A0 => N3138, A1 => mult_21_C245_n1543,
                           SL => mult_21_C245_n71, Z => mult_21_C245_n864);
   mult_21_C245_U709 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n69, SL => mult_21_C245_n864, Z => 
                           mult_21_C245_n1167);
   mult_21_C245_U708 : MUXB2DL port map( A0 => N3139, A1 => N3138, SL => 
                           mult_21_C245_n71, Z => mult_21_C245_n863);
   mult_21_C245_U707 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n69, SL => mult_21_C245_n863, Z => 
                           mult_21_C245_n1166);
   mult_21_C245_U706 : MUXB2DL port map( A0 => N3140, A1 => N3139, SL => 
                           mult_21_C245_n71, Z => mult_21_C245_n862);
   mult_21_C245_U705 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n69, SL => mult_21_C245_n862, Z => 
                           mult_21_C245_n1165);
   mult_21_C245_U704 : MUXB2DL port map( A0 => N3141, A1 => N3140, SL => 
                           mult_21_C245_n71, Z => mult_21_C245_n861);
   mult_21_C245_U703 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n69, SL => mult_21_C245_n861, Z => 
                           mult_21_C245_n1164);
   mult_21_C245_U702 : MUXB2DL port map( A0 => N3142, A1 => N3141, SL => 
                           mult_21_C245_n71, Z => mult_21_C245_n860);
   mult_21_C245_U701 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n69, SL => mult_21_C245_n860, Z => 
                           mult_21_C245_n1163);
   mult_21_C245_U700 : MUXB2DL port map( A0 => N3143, A1 => N3142, SL => 
                           mult_21_C245_n71, Z => mult_21_C245_n859);
   mult_21_C245_U699 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n69, SL => mult_21_C245_n859, Z => 
                           mult_21_C245_n1162);
   mult_21_C245_U698 : MUXB2DL port map( A0 => N3144, A1 => N3143, SL => 
                           mult_21_C245_n71, Z => mult_21_C245_n858);
   mult_21_C245_U697 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n69, SL => mult_21_C245_n858, Z => 
                           mult_21_C245_n1161);
   mult_21_C245_U696 : MUXB2DL port map( A0 => N3145, A1 => N3144, SL => 
                           mult_21_C245_n71, Z => mult_21_C245_n857);
   mult_21_C245_U695 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n69, SL => mult_21_C245_n857, Z => 
                           mult_21_C245_n1160);
   mult_21_C245_U694 : MUXB2DL port map( A0 => N3146, A1 => N3145, SL => 
                           mult_21_C245_n71, Z => mult_21_C245_n856);
   mult_21_C245_U693 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n69, SL => mult_21_C245_n856, Z => 
                           mult_21_C245_n1159);
   mult_21_C245_U692 : MUXB2DL port map( A0 => N3147, A1 => N3146, SL => 
                           mult_21_C245_n71, Z => mult_21_C245_n855);
   mult_21_C245_U691 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n69, SL => mult_21_C245_n855, Z => 
                           mult_21_C245_n1158);
   mult_21_C245_U690 : MUXB2DL port map( A0 => N3148, A1 => N3147, SL => 
                           mult_21_C245_n71, Z => mult_21_C245_n854);
   mult_21_C245_U689 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n69, SL => mult_21_C245_n854, Z => 
                           mult_21_C245_n1157);
   mult_21_C245_U688 : MUXB2DL port map( A0 => N3149, A1 => N3148, SL => 
                           mult_21_C245_n71, Z => mult_21_C245_n853);
   mult_21_C245_U687 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n69, SL => mult_21_C245_n853, Z => 
                           mult_21_C245_n1156);
   mult_21_C245_U686 : MUXB2DL port map( A0 => N3150, A1 => N3149, SL => 
                           mult_21_C245_n71, Z => mult_21_C245_n852);
   mult_21_C245_U685 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n69, SL => mult_21_C245_n852, Z => 
                           mult_21_C245_n1155);
   mult_21_C245_U684 : MUXB2DL port map( A0 => N3151, A1 => N3150, SL => 
                           mult_21_C245_n71, Z => mult_21_C245_n851);
   mult_21_C245_U683 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n69, SL => mult_21_C245_n851, Z => 
                           mult_21_C245_n1154);
   mult_21_C245_U682 : MUXB2DL port map( A0 => N3152, A1 => N3151, SL => 
                           mult_21_C245_n71, Z => mult_21_C245_n850);
   mult_21_C245_U681 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n69, SL => mult_21_C245_n850, Z => 
                           mult_21_C245_n1153);
   mult_21_C245_U680 : NOR2M1D1 port map( A1 => mult_21_C245_n66, A2 => 
                           mult_21_C245_n69, Z => mult_21_C245_n1088);
   mult_21_C245_U679 : NAN2M1D1 port map( A1 => mult_21_C245_n78, A2 => 
                           mult_21_C245_n1543, Z => mult_21_C245_n849);
   mult_21_C245_U678 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n76, SL => mult_21_C245_n849, Z => 
                           mult_21_C245_n1152);
   mult_21_C245_U677 : MUXB2DL port map( A0 => N3138, A1 => mult_21_C245_n1543,
                           SL => mult_21_C245_n78, Z => mult_21_C245_n848);
   mult_21_C245_U676 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n76, SL => mult_21_C245_n848, Z => 
                           mult_21_C245_n1151);
   mult_21_C245_U675 : MUXB2DL port map( A0 => N3139, A1 => N3138, SL => 
                           mult_21_C245_n78, Z => mult_21_C245_n847);
   mult_21_C245_U674 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n76, SL => mult_21_C245_n847, Z => 
                           mult_21_C245_n1150);
   mult_21_C245_U673 : MUXB2DL port map( A0 => N3140, A1 => N3139, SL => 
                           mult_21_C245_n78, Z => mult_21_C245_n846);
   mult_21_C245_U672 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n76, SL => mult_21_C245_n846, Z => 
                           mult_21_C245_n1149);
   mult_21_C245_U671 : MUXB2DL port map( A0 => N3141, A1 => N3140, SL => 
                           mult_21_C245_n78, Z => mult_21_C245_n845);
   mult_21_C245_U670 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n76, SL => mult_21_C245_n845, Z => 
                           mult_21_C245_n1148);
   mult_21_C245_U669 : MUXB2DL port map( A0 => N3142, A1 => N3141, SL => 
                           mult_21_C245_n78, Z => mult_21_C245_n844);
   mult_21_C245_U668 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n76, SL => mult_21_C245_n844, Z => 
                           mult_21_C245_n1147);
   mult_21_C245_U667 : MUXB2DL port map( A0 => N3143, A1 => N3142, SL => 
                           mult_21_C245_n78, Z => mult_21_C245_n843);
   mult_21_C245_U666 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n76, SL => mult_21_C245_n843, Z => 
                           mult_21_C245_n1146);
   mult_21_C245_U665 : MUXB2DL port map( A0 => N3144, A1 => N3143, SL => 
                           mult_21_C245_n78, Z => mult_21_C245_n842);
   mult_21_C245_U664 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n76, SL => mult_21_C245_n842, Z => 
                           mult_21_C245_n1145);
   mult_21_C245_U663 : MUXB2DL port map( A0 => N3145, A1 => N3144, SL => 
                           mult_21_C245_n78, Z => mult_21_C245_n841);
   mult_21_C245_U662 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n76, SL => mult_21_C245_n841, Z => 
                           mult_21_C245_n1144);
   mult_21_C245_U661 : MUXB2DL port map( A0 => N3146, A1 => N3145, SL => 
                           mult_21_C245_n78, Z => mult_21_C245_n840);
   mult_21_C245_U660 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n76, SL => mult_21_C245_n840, Z => 
                           mult_21_C245_n1143);
   mult_21_C245_U659 : MUXB2DL port map( A0 => N3147, A1 => N3146, SL => 
                           mult_21_C245_n78, Z => mult_21_C245_n839);
   mult_21_C245_U658 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n76, SL => mult_21_C245_n839, Z => 
                           mult_21_C245_n1142);
   mult_21_C245_U657 : MUXB2DL port map( A0 => N3148, A1 => N3147, SL => 
                           mult_21_C245_n78, Z => mult_21_C245_n838);
   mult_21_C245_U656 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n76, SL => mult_21_C245_n838, Z => 
                           mult_21_C245_n1141);
   mult_21_C245_U655 : MUXB2DL port map( A0 => N3149, A1 => N3148, SL => 
                           mult_21_C245_n78, Z => mult_21_C245_n837);
   mult_21_C245_U654 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n76, SL => mult_21_C245_n837, Z => 
                           mult_21_C245_n1140);
   mult_21_C245_U653 : MUXB2DL port map( A0 => N3150, A1 => N3149, SL => 
                           mult_21_C245_n78, Z => mult_21_C245_n836);
   mult_21_C245_U652 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n76, SL => mult_21_C245_n836, Z => 
                           mult_21_C245_n1139);
   mult_21_C245_U651 : NOR2M1D1 port map( A1 => mult_21_C245_n73, A2 => 
                           mult_21_C245_n76, Z => mult_21_C245_n1087);
   mult_21_C245_U650 : NAN2M1D1 port map( A1 => mult_21_C245_n83, A2 => N3137, 
                           Z => mult_21_C245_n835);
   mult_21_C245_U649 : MUXB2DL port map( A0 => mult_21_C245_n79, A1 => 
                           mult_21_C245_n81, SL => mult_21_C245_n835, Z => 
                           mult_21_C245_n1138);
   mult_21_C245_U648 : MUXB2DL port map( A0 => N3138, A1 => mult_21_C245_n1543,
                           SL => mult_21_C245_n83, Z => mult_21_C245_n834);
   mult_21_C245_U647 : MUXB2DL port map( A0 => mult_21_C245_n79, A1 => 
                           mult_21_C245_n81, SL => mult_21_C245_n834, Z => 
                           mult_21_C245_n1137);
   mult_21_C245_U646 : MUXB2DL port map( A0 => N3139, A1 => N3138, SL => 
                           mult_21_C245_n83, Z => mult_21_C245_n833);
   mult_21_C245_U645 : MUXB2DL port map( A0 => mult_21_C245_n79, A1 => 
                           mult_21_C245_n81, SL => mult_21_C245_n833, Z => 
                           mult_21_C245_n1136);
   mult_21_C245_U644 : MUXB2DL port map( A0 => N3140, A1 => N3139, SL => 
                           mult_21_C245_n83, Z => mult_21_C245_n832);
   mult_21_C245_U643 : MUXB2DL port map( A0 => mult_21_C245_n79, A1 => 
                           mult_21_C245_n81, SL => mult_21_C245_n832, Z => 
                           mult_21_C245_n1135);
   mult_21_C245_U642 : MUXB2DL port map( A0 => N3141, A1 => N3140, SL => 
                           mult_21_C245_n83, Z => mult_21_C245_n831);
   mult_21_C245_U641 : MUXB2DL port map( A0 => mult_21_C245_n79, A1 => 
                           mult_21_C245_n81, SL => mult_21_C245_n831, Z => 
                           mult_21_C245_n1134);
   mult_21_C245_U640 : MUXB2DL port map( A0 => N3142, A1 => N3141, SL => 
                           mult_21_C245_n83, Z => mult_21_C245_n830);
   mult_21_C245_U639 : MUXB2DL port map( A0 => mult_21_C245_n79, A1 => 
                           mult_21_C245_n81, SL => mult_21_C245_n830, Z => 
                           mult_21_C245_n1133);
   mult_21_C245_U638 : MUXB2DL port map( A0 => N3143, A1 => N3142, SL => 
                           mult_21_C245_n83, Z => mult_21_C245_n829);
   mult_21_C245_U637 : MUXB2DL port map( A0 => mult_21_C245_n79, A1 => 
                           mult_21_C245_n81, SL => mult_21_C245_n829, Z => 
                           mult_21_C245_n1132);
   mult_21_C245_U636 : MUXB2DL port map( A0 => N3144, A1 => N3143, SL => 
                           mult_21_C245_n83, Z => mult_21_C245_n828);
   mult_21_C245_U635 : MUXB2DL port map( A0 => mult_21_C245_n79, A1 => 
                           mult_21_C245_n81, SL => mult_21_C245_n828, Z => 
                           mult_21_C245_n1131);
   mult_21_C245_U634 : MUXB2DL port map( A0 => N3145, A1 => N3144, SL => 
                           mult_21_C245_n83, Z => mult_21_C245_n827);
   mult_21_C245_U633 : MUXB2DL port map( A0 => mult_21_C245_n79, A1 => 
                           mult_21_C245_n81, SL => mult_21_C245_n827, Z => 
                           mult_21_C245_n1130);
   mult_21_C245_U632 : MUXB2DL port map( A0 => N3146, A1 => N3145, SL => 
                           mult_21_C245_n83, Z => mult_21_C245_n826);
   mult_21_C245_U631 : MUXB2DL port map( A0 => mult_21_C245_n79, A1 => 
                           mult_21_C245_n81, SL => mult_21_C245_n826, Z => 
                           mult_21_C245_n1129);
   mult_21_C245_U630 : MUXB2DL port map( A0 => N3147, A1 => N3146, SL => 
                           mult_21_C245_n83, Z => mult_21_C245_n825);
   mult_21_C245_U629 : MUXB2DL port map( A0 => mult_21_C245_n79, A1 => 
                           mult_21_C245_n81, SL => mult_21_C245_n825, Z => 
                           mult_21_C245_n1128);
   mult_21_C245_U628 : MUXB2DL port map( A0 => N3148, A1 => N3147, SL => 
                           mult_21_C245_n83, Z => mult_21_C245_n824);
   mult_21_C245_U627 : MUXB2DL port map( A0 => mult_21_C245_n79, A1 => 
                           mult_21_C245_n81, SL => mult_21_C245_n824, Z => 
                           mult_21_C245_n1127);
   mult_21_C245_U626 : NOR2M1D1 port map( A1 => mult_21_C245_n79, A2 => 
                           mult_21_C245_n81, Z => mult_21_C245_n1086);
   mult_21_C245_U625 : NAN2M1D1 port map( A1 => mult_21_C245_n88, A2 => 
                           mult_21_C245_n1543, Z => mult_21_C245_n823);
   mult_21_C245_U624 : MUXB2DL port map( A0 => mult_21_C245_n84, A1 => 
                           mult_21_C245_n86, SL => mult_21_C245_n823, Z => 
                           mult_21_C245_n1126);
   mult_21_C245_U623 : MUXB2DL port map( A0 => N3138, A1 => mult_21_C245_n1543,
                           SL => mult_21_C245_n88, Z => mult_21_C245_n822);
   mult_21_C245_U622 : MUXB2DL port map( A0 => mult_21_C245_n84, A1 => 
                           mult_21_C245_n86, SL => mult_21_C245_n822, Z => 
                           mult_21_C245_n1125);
   mult_21_C245_U621 : MUXB2DL port map( A0 => N3139, A1 => N3138, SL => 
                           mult_21_C245_n88, Z => mult_21_C245_n821);
   mult_21_C245_U620 : MUXB2DL port map( A0 => mult_21_C245_n84, A1 => 
                           mult_21_C245_n86, SL => mult_21_C245_n821, Z => 
                           mult_21_C245_n1124);
   mult_21_C245_U619 : MUXB2DL port map( A0 => N3140, A1 => N3139, SL => 
                           mult_21_C245_n88, Z => mult_21_C245_n820);
   mult_21_C245_U618 : MUXB2DL port map( A0 => mult_21_C245_n84, A1 => 
                           mult_21_C245_n86, SL => mult_21_C245_n820, Z => 
                           mult_21_C245_n1123);
   mult_21_C245_U617 : MUXB2DL port map( A0 => N3141, A1 => N3140, SL => 
                           mult_21_C245_n88, Z => mult_21_C245_n819);
   mult_21_C245_U616 : MUXB2DL port map( A0 => mult_21_C245_n84, A1 => 
                           mult_21_C245_n86, SL => mult_21_C245_n819, Z => 
                           mult_21_C245_n1122);
   mult_21_C245_U615 : MUXB2DL port map( A0 => N3142, A1 => N3141, SL => 
                           mult_21_C245_n88, Z => mult_21_C245_n818);
   mult_21_C245_U614 : MUXB2DL port map( A0 => mult_21_C245_n84, A1 => 
                           mult_21_C245_n86, SL => mult_21_C245_n818, Z => 
                           mult_21_C245_n1121);
   mult_21_C245_U613 : MUXB2DL port map( A0 => N3143, A1 => N3142, SL => 
                           mult_21_C245_n88, Z => mult_21_C245_n817);
   mult_21_C245_U612 : MUXB2DL port map( A0 => mult_21_C245_n84, A1 => 
                           mult_21_C245_n86, SL => mult_21_C245_n817, Z => 
                           mult_21_C245_n1120);
   mult_21_C245_U611 : MUXB2DL port map( A0 => N3144, A1 => N3143, SL => 
                           mult_21_C245_n88, Z => mult_21_C245_n816);
   mult_21_C245_U610 : MUXB2DL port map( A0 => mult_21_C245_n84, A1 => 
                           mult_21_C245_n86, SL => mult_21_C245_n816, Z => 
                           mult_21_C245_n1119);
   mult_21_C245_U609 : MUXB2DL port map( A0 => N3145, A1 => N3144, SL => 
                           mult_21_C245_n88, Z => mult_21_C245_n815);
   mult_21_C245_U608 : MUXB2DL port map( A0 => mult_21_C245_n84, A1 => 
                           mult_21_C245_n86, SL => mult_21_C245_n815, Z => 
                           mult_21_C245_n1118);
   mult_21_C245_U607 : MUXB2DL port map( A0 => N3146, A1 => N3145, SL => 
                           mult_21_C245_n88, Z => mult_21_C245_n814);
   mult_21_C245_U606 : MUXB2DL port map( A0 => mult_21_C245_n84, A1 => 
                           mult_21_C245_n86, SL => mult_21_C245_n814, Z => 
                           mult_21_C245_n1117);
   mult_21_C245_U605 : NOR2M1D1 port map( A1 => mult_21_C245_n84, A2 => 
                           mult_21_C245_n86, Z => mult_21_C245_n1085);
   mult_21_C245_U604 : NAN2M1D1 port map( A1 => mult_21_C245_n93, A2 => 
                           mult_21_C245_n1543, Z => mult_21_C245_n813);
   mult_21_C245_U603 : MUXB2DL port map( A0 => mult_21_C245_n89, A1 => 
                           mult_21_C245_n91, SL => mult_21_C245_n813, Z => 
                           mult_21_C245_n1116);
   mult_21_C245_U602 : MUXB2DL port map( A0 => N3138, A1 => mult_21_C245_n1543,
                           SL => mult_21_C245_n93, Z => mult_21_C245_n812);
   mult_21_C245_U601 : MUXB2DL port map( A0 => mult_21_C245_n89, A1 => 
                           mult_21_C245_n91, SL => mult_21_C245_n812, Z => 
                           mult_21_C245_n1115);
   mult_21_C245_U600 : MUXB2DL port map( A0 => N3139, A1 => N3138, SL => 
                           mult_21_C245_n93, Z => mult_21_C245_n811);
   mult_21_C245_U599 : MUXB2DL port map( A0 => mult_21_C245_n89, A1 => 
                           mult_21_C245_n91, SL => mult_21_C245_n811, Z => 
                           mult_21_C245_n1114);
   mult_21_C245_U598 : MUXB2DL port map( A0 => N3140, A1 => N3139, SL => 
                           mult_21_C245_n93, Z => mult_21_C245_n810);
   mult_21_C245_U597 : MUXB2DL port map( A0 => mult_21_C245_n89, A1 => 
                           mult_21_C245_n91, SL => mult_21_C245_n810, Z => 
                           mult_21_C245_n1113);
   mult_21_C245_U596 : MUXB2DL port map( A0 => N3141, A1 => N3140, SL => 
                           mult_21_C245_n93, Z => mult_21_C245_n809);
   mult_21_C245_U595 : MUXB2DL port map( A0 => mult_21_C245_n89, A1 => 
                           mult_21_C245_n91, SL => mult_21_C245_n809, Z => 
                           mult_21_C245_n1112);
   mult_21_C245_U594 : MUXB2DL port map( A0 => N3142, A1 => N3141, SL => 
                           mult_21_C245_n93, Z => mult_21_C245_n808);
   mult_21_C245_U593 : MUXB2DL port map( A0 => mult_21_C245_n89, A1 => 
                           mult_21_C245_n91, SL => mult_21_C245_n808, Z => 
                           mult_21_C245_n1111);
   mult_21_C245_U592 : MUXB2DL port map( A0 => N3143, A1 => N3142, SL => 
                           mult_21_C245_n93, Z => mult_21_C245_n807);
   mult_21_C245_U591 : MUXB2DL port map( A0 => mult_21_C245_n89, A1 => 
                           mult_21_C245_n91, SL => mult_21_C245_n807, Z => 
                           mult_21_C245_n1110);
   mult_21_C245_U590 : MUXB2DL port map( A0 => N3144, A1 => N3143, SL => 
                           mult_21_C245_n93, Z => mult_21_C245_n806);
   mult_21_C245_U589 : MUXB2DL port map( A0 => mult_21_C245_n89, A1 => 
                           mult_21_C245_n91, SL => mult_21_C245_n806, Z => 
                           mult_21_C245_n1109);
   mult_21_C245_U588 : NOR2M1D1 port map( A1 => mult_21_C245_n89, A2 => 
                           mult_21_C245_n91, Z => mult_21_C245_n1084);
   mult_21_C245_U587 : NAN2M1D1 port map( A1 => mult_21_C245_n98, A2 => N3137, 
                           Z => mult_21_C245_n805);
   mult_21_C245_U586 : MUXB2DL port map( A0 => mult_21_C245_n94, A1 => 
                           mult_21_C245_n96, SL => mult_21_C245_n805, Z => 
                           mult_21_C245_n1108);
   mult_21_C245_U585 : MUXB2DL port map( A0 => N3138, A1 => mult_21_C245_n1543,
                           SL => mult_21_C245_n98, Z => mult_21_C245_n804);
   mult_21_C245_U584 : MUXB2DL port map( A0 => mult_21_C245_n94, A1 => 
                           mult_21_C245_n96, SL => mult_21_C245_n804, Z => 
                           mult_21_C245_n1107);
   mult_21_C245_U583 : MUXB2DL port map( A0 => N3139, A1 => N3138, SL => 
                           mult_21_C245_n98, Z => mult_21_C245_n803);
   mult_21_C245_U582 : MUXB2DL port map( A0 => mult_21_C245_n94, A1 => 
                           mult_21_C245_n96, SL => mult_21_C245_n803, Z => 
                           mult_21_C245_n1106);
   mult_21_C245_U581 : MUXB2DL port map( A0 => N3140, A1 => N3139, SL => 
                           mult_21_C245_n98, Z => mult_21_C245_n802);
   mult_21_C245_U580 : MUXB2DL port map( A0 => mult_21_C245_n94, A1 => 
                           mult_21_C245_n96, SL => mult_21_C245_n802, Z => 
                           mult_21_C245_n1105);
   mult_21_C245_U579 : MUXB2DL port map( A0 => N3141, A1 => N3140, SL => 
                           mult_21_C245_n98, Z => mult_21_C245_n801);
   mult_21_C245_U578 : MUXB2DL port map( A0 => mult_21_C245_n94, A1 => 
                           mult_21_C245_n96, SL => mult_21_C245_n801, Z => 
                           mult_21_C245_n1104);
   mult_21_C245_U577 : MUXB2DL port map( A0 => N3142, A1 => N3141, SL => 
                           mult_21_C245_n98, Z => mult_21_C245_n800);
   mult_21_C245_U576 : MUXB2DL port map( A0 => mult_21_C245_n94, A1 => 
                           mult_21_C245_n96, SL => mult_21_C245_n800, Z => 
                           mult_21_C245_n1103);
   mult_21_C245_U575 : NOR2M1D1 port map( A1 => mult_21_C245_n94, A2 => 
                           mult_21_C245_n96, Z => mult_21_C245_n1083);
   mult_21_C245_U574 : NAN2M1D1 port map( A1 => mult_21_C245_n103, A2 => N3137,
                           Z => mult_21_C245_n799);
   mult_21_C245_U573 : MUXB2DL port map( A0 => mult_21_C245_n99, A1 => 
                           mult_21_C245_n101, SL => mult_21_C245_n799, Z => 
                           mult_21_C245_n1102);
   mult_21_C245_U572 : MUXB2DL port map( A0 => N3138, A1 => mult_21_C245_n1543,
                           SL => mult_21_C245_n103, Z => mult_21_C245_n798);
   mult_21_C245_U571 : MUXB2DL port map( A0 => mult_21_C245_n99, A1 => 
                           mult_21_C245_n101, SL => mult_21_C245_n798, Z => 
                           mult_21_C245_n1101);
   mult_21_C245_U570 : MUXB2DL port map( A0 => N3139, A1 => N3138, SL => 
                           mult_21_C245_n103, Z => mult_21_C245_n797);
   mult_21_C245_U569 : MUXB2DL port map( A0 => mult_21_C245_n99, A1 => 
                           mult_21_C245_n101, SL => mult_21_C245_n797, Z => 
                           mult_21_C245_n1100);
   mult_21_C245_U568 : MUXB2DL port map( A0 => N3140, A1 => N3139, SL => 
                           mult_21_C245_n103, Z => mult_21_C245_n796);
   mult_21_C245_U567 : MUXB2DL port map( A0 => mult_21_C245_n99, A1 => 
                           mult_21_C245_n101, SL => mult_21_C245_n796, Z => 
                           mult_21_C245_n1099);
   mult_21_C245_U566 : NOR2M1D1 port map( A1 => mult_21_C245_n99, A2 => 
                           mult_21_C245_n101, Z => mult_21_C245_n1082);
   mult_21_C245_U565 : NAN2M1D1 port map( A1 => mult_21_C245_n106, A2 => N3137,
                           Z => mult_21_C245_n795);
   mult_21_C245_U564 : MUXB2DL port map( A0 => mult_21_C245_n104, A1 => 
                           mult_21_C245_n105, SL => mult_21_C245_n795, Z => 
                           mult_21_C245_n1098);
   mult_21_C245_U563 : MUXB2DL port map( A0 => N3138, A1 => mult_21_C245_n1543,
                           SL => mult_21_C245_n106, Z => mult_21_C245_n794);
   mult_21_C245_U562 : MUXB2DL port map( A0 => mult_21_C245_n104, A1 => 
                           mult_21_C245_n105, SL => mult_21_C245_n794, Z => 
                           mult_21_C245_n1097);
   mult_21_C245_U561 : NOR2M1D1 port map( A1 => mult_21_C245_n104, A2 => 
                           mult_21_C245_n105, Z => mult_21_C245_n1081);
   mult_21_C245_U557 : ADFULD1 port map( A => mult_21_C245_n1334, B => 
                           mult_21_C245_n1364, CI => mult_21_C245_n790, CO => 
                           mult_21_C245_n786, S => mult_21_C245_n787);
   mult_21_C245_U555 : ADFULD1 port map( A => mult_21_C245_n788, B => 
                           mult_21_C245_n1305, CI => mult_21_C245_n785, CO => 
                           mult_21_C245_n782, S => mult_21_C245_n783);
   mult_21_C245_U553 : ADFULD1 port map( A => mult_21_C245_n1304, B => 
                           mult_21_C245_n1362, CI => mult_21_C245_n1332, CO => 
                           mult_21_C245_n778, S => mult_21_C245_n779);
   mult_21_C245_U552 : ADFULD1 port map( A => mult_21_C245_n781, B => 
                           mult_21_C245_n784, CI => mult_21_C245_n779, CO => 
                           mult_21_C245_n776, S => mult_21_C245_n777);
   mult_21_C245_U550 : ADFULD1 port map( A => mult_21_C245_n1277, B => 
                           mult_21_C245_n1303, CI => mult_21_C245_n780, CO => 
                           mult_21_C245_n772, S => mult_21_C245_n773);
   mult_21_C245_U549 : ADFULD1 port map( A => mult_21_C245_n778, B => 
                           mult_21_C245_n775, CI => mult_21_C245_n773, CO => 
                           mult_21_C245_n770, S => mult_21_C245_n771);
   mult_21_C245_U547 : ADFULD1 port map( A => mult_21_C245_n1276, B => 
                           mult_21_C245_n1360, CI => mult_21_C245_n1330, CO => 
                           mult_21_C245_n766, S => mult_21_C245_n767);
   mult_21_C245_U546 : ADFULD1 port map( A => mult_21_C245_n774, B => 
                           mult_21_C245_n1302, CI => mult_21_C245_n769, CO => 
                           mult_21_C245_n764, S => mult_21_C245_n765);
   mult_21_C245_U545 : ADFULD1 port map( A => mult_21_C245_n767, B => 
                           mult_21_C245_n772, CI => mult_21_C245_n765, CO => 
                           mult_21_C245_n762, S => mult_21_C245_n763);
   mult_21_C245_U543 : ADFULD1 port map( A => mult_21_C245_n1275, B => 
                           mult_21_C245_n1251, CI => mult_21_C245_n1301, CO => 
                           mult_21_C245_n758, S => mult_21_C245_n759);
   mult_21_C245_U542 : ADFULD1 port map( A => mult_21_C245_n761, B => 
                           mult_21_C245_n768, CI => mult_21_C245_n766, CO => 
                           mult_21_C245_n756, S => mult_21_C245_n757);
   mult_21_C245_U541 : ADFULD1 port map( A => mult_21_C245_n764, B => 
                           mult_21_C245_n759, CI => mult_21_C245_n757, CO => 
                           mult_21_C245_n754, S => mult_21_C245_n755);
   mult_21_C245_U539 : ADFULD1 port map( A => mult_21_C245_n1250, B => 
                           mult_21_C245_n1358, CI => mult_21_C245_n1328, CO => 
                           mult_21_C245_n750, S => mult_21_C245_n751);
   mult_21_C245_U538 : ADFULD1 port map( A => mult_21_C245_n1274, B => 
                           mult_21_C245_n1300, CI => mult_21_C245_n760, CO => 
                           mult_21_C245_n748, S => mult_21_C245_n749);
   mult_21_C245_U537 : ADFULD1 port map( A => mult_21_C245_n758, B => 
                           mult_21_C245_n753, CI => mult_21_C245_n751, CO => 
                           mult_21_C245_n746, S => mult_21_C245_n747);
   mult_21_C245_U536 : ADFULD1 port map( A => mult_21_C245_n756, B => 
                           mult_21_C245_n749, CI => mult_21_C245_n747, CO => 
                           mult_21_C245_n744, S => mult_21_C245_n745);
   mult_21_C245_U534 : ADFULD1 port map( A => mult_21_C245_n1273, B => 
                           mult_21_C245_n1249, CI => mult_21_C245_n1227, CO => 
                           mult_21_C245_n740, S => mult_21_C245_n741);
   mult_21_C245_U533 : ADFULD1 port map( A => mult_21_C245_n752, B => 
                           mult_21_C245_n1299, CI => mult_21_C245_n743, CO => 
                           mult_21_C245_n738, S => mult_21_C245_n739);
   mult_21_C245_U532 : ADFULD1 port map( A => mult_21_C245_n748, B => 
                           mult_21_C245_n750, CI => mult_21_C245_n741, CO => 
                           mult_21_C245_n736, S => mult_21_C245_n737);
   mult_21_C245_U531 : ADFULD1 port map( A => mult_21_C245_n746, B => 
                           mult_21_C245_n739, CI => mult_21_C245_n737, CO => 
                           mult_21_C245_n734, S => mult_21_C245_n735);
   mult_21_C245_U529 : ADFULD1 port map( A => mult_21_C245_n1248, B => 
                           mult_21_C245_n1356, CI => mult_21_C245_n1326, CO => 
                           mult_21_C245_n730, S => mult_21_C245_n731);
   mult_21_C245_U528 : ADFULD1 port map( A => mult_21_C245_n1272, B => 
                           mult_21_C245_n1298, CI => mult_21_C245_n1226, CO => 
                           mult_21_C245_n728, S => mult_21_C245_n729);
   mult_21_C245_U527 : ADFULD1 port map( A => mult_21_C245_n733, B => 
                           mult_21_C245_n742, CI => mult_21_C245_n740, CO => 
                           mult_21_C245_n726, S => mult_21_C245_n727);
   mult_21_C245_U526 : ADFULD1 port map( A => mult_21_C245_n729, B => 
                           mult_21_C245_n731, CI => mult_21_C245_n738, CO => 
                           mult_21_C245_n724, S => mult_21_C245_n725);
   mult_21_C245_U525 : ADFULD1 port map( A => mult_21_C245_n736, B => 
                           mult_21_C245_n727, CI => mult_21_C245_n725, CO => 
                           mult_21_C245_n722, S => mult_21_C245_n723);
   mult_21_C245_U523 : ADFULD1 port map( A => mult_21_C245_n1271, B => 
                           mult_21_C245_n1297, CI => mult_21_C245_n1225, CO => 
                           mult_21_C245_n718, S => mult_21_C245_n719);
   mult_21_C245_U522 : ADFULD1 port map( A => mult_21_C245_n1205, B => 
                           mult_21_C245_n1247, CI => mult_21_C245_n732, CO => 
                           mult_21_C245_n716, S => mult_21_C245_n717);
   mult_21_C245_U521 : ADFULD1 port map( A => mult_21_C245_n730, B => 
                           mult_21_C245_n721, CI => mult_21_C245_n728, CO => 
                           mult_21_C245_n714, S => mult_21_C245_n715);
   mult_21_C245_U520 : ADFULD1 port map( A => mult_21_C245_n717, B => 
                           mult_21_C245_n719, CI => mult_21_C245_n726, CO => 
                           mult_21_C245_n712, S => mult_21_C245_n713);
   mult_21_C245_U519 : ADFULD1 port map( A => mult_21_C245_n724, B => 
                           mult_21_C245_n715, CI => mult_21_C245_n713, CO => 
                           mult_21_C245_n710, S => mult_21_C245_n711);
   mult_21_C245_U517 : ADFULD1 port map( A => mult_21_C245_n1204, B => 
                           mult_21_C245_n1354, CI => mult_21_C245_n1324, CO => 
                           mult_21_C245_n706, S => mult_21_C245_n707);
   mult_21_C245_U516 : ADFULD1 port map( A => mult_21_C245_n1246, B => 
                           mult_21_C245_n1296, CI => mult_21_C245_n1224, CO => 
                           mult_21_C245_n704, S => mult_21_C245_n705);
   mult_21_C245_U515 : ADFULD1 port map( A => mult_21_C245_n720, B => 
                           mult_21_C245_n1270, CI => mult_21_C245_n709, CO => 
                           mult_21_C245_n702, S => mult_21_C245_n703);
   mult_21_C245_U514 : ADFULD1 port map( A => mult_21_C245_n716, B => 
                           mult_21_C245_n718, CI => mult_21_C245_n707, CO => 
                           mult_21_C245_n700, S => mult_21_C245_n701);
   mult_21_C245_U513 : ADFULD1 port map( A => mult_21_C245_n703, B => 
                           mult_21_C245_n705, CI => mult_21_C245_n714, CO => 
                           mult_21_C245_n698, S => mult_21_C245_n699);
   mult_21_C245_U512 : ADFULD1 port map( A => mult_21_C245_n712, B => 
                           mult_21_C245_n701, CI => mult_21_C245_n699, CO => 
                           mult_21_C245_n696, S => mult_21_C245_n697);
   mult_21_C245_U510 : ADFULD1 port map( A => mult_21_C245_n1295, B => 
                           mult_21_C245_n1269, CI => mult_21_C245_n1223, CO => 
                           mult_21_C245_n692, S => mult_21_C245_n693);
   mult_21_C245_U509 : ADFULD1 port map( A => mult_21_C245_n1185, B => 
                           mult_21_C245_n1245, CI => mult_21_C245_n1203, CO => 
                           mult_21_C245_n690, S => mult_21_C245_n691);
   mult_21_C245_U508 : ADFULD1 port map( A => mult_21_C245_n695, B => 
                           mult_21_C245_n708, CI => mult_21_C245_n706, CO => 
                           mult_21_C245_n688, S => mult_21_C245_n689);
   mult_21_C245_U507 : ADFULD1 port map( A => mult_21_C245_n691, B => 
                           mult_21_C245_n704, CI => mult_21_C245_n693, CO => 
                           mult_21_C245_n686, S => mult_21_C245_n687);
   mult_21_C245_U506 : ADFULD1 port map( A => mult_21_C245_n700, B => 
                           mult_21_C245_n702, CI => mult_21_C245_n689, CO => 
                           mult_21_C245_n684, S => mult_21_C245_n685);
   mult_21_C245_U505 : ADFULD1 port map( A => mult_21_C245_n698, B => 
                           mult_21_C245_n687, CI => mult_21_C245_n685, CO => 
                           mult_21_C245_n682, S => mult_21_C245_n683);
   mult_21_C245_U503 : ADFULD1 port map( A => mult_21_C245_n1202, B => 
                           mult_21_C245_n1352, CI => mult_21_C245_n1322, CO => 
                           mult_21_C245_n678, S => mult_21_C245_n679);
   mult_21_C245_U502 : ADFULD1 port map( A => mult_21_C245_n1184, B => 
                           mult_21_C245_n1268, CI => mult_21_C245_n1222, CO => 
                           mult_21_C245_n676, S => mult_21_C245_n677);
   mult_21_C245_U501 : ADFULD1 port map( A => mult_21_C245_n1244, B => 
                           mult_21_C245_n1294, CI => mult_21_C245_n694, CO => 
                           mult_21_C245_n674, S => mult_21_C245_n675);
   mult_21_C245_U500 : ADFULD1 port map( A => mult_21_C245_n692, B => 
                           mult_21_C245_n681, CI => mult_21_C245_n690, CO => 
                           mult_21_C245_n672, S => mult_21_C245_n673);
   mult_21_C245_U499 : ADFULD1 port map( A => mult_21_C245_n677, B => 
                           mult_21_C245_n679, CI => mult_21_C245_n675, CO => 
                           mult_21_C245_n670, S => mult_21_C245_n671);
   mult_21_C245_U498 : ADFULD1 port map( A => mult_21_C245_n686, B => 
                           mult_21_C245_n688, CI => mult_21_C245_n673, CO => 
                           mult_21_C245_n668, S => mult_21_C245_n669);
   mult_21_C245_U497 : ADFULD1 port map( A => mult_21_C245_n684, B => 
                           mult_21_C245_n671, CI => mult_21_C245_n669, CO => 
                           mult_21_C245_n666, S => mult_21_C245_n667);
   mult_21_C245_U495 : ADFULD1 port map( A => mult_21_C245_n1293, B => 
                           mult_21_C245_n1201, CI => mult_21_C245_n1221, CO => 
                           mult_21_C245_n662, S => mult_21_C245_n663);
   mult_21_C245_U494 : ADFULD1 port map( A => mult_21_C245_n1183, B => 
                           mult_21_C245_n1167, CI => mult_21_C245_n1243, CO => 
                           mult_21_C245_n660, S => mult_21_C245_n661);
   mult_21_C245_U493 : ADFULD1 port map( A => mult_21_C245_n680, B => 
                           mult_21_C245_n1267, CI => mult_21_C245_n665, CO => 
                           mult_21_C245_n658, S => mult_21_C245_n659);
   mult_21_C245_U492 : ADFULD1 port map( A => mult_21_C245_n676, B => 
                           mult_21_C245_n678, CI => mult_21_C245_n674, CO => 
                           mult_21_C245_n656, S => mult_21_C245_n657);
   mult_21_C245_U491 : ADFULD1 port map( A => mult_21_C245_n663, B => 
                           mult_21_C245_n661, CI => mult_21_C245_n672, CO => 
                           mult_21_C245_n654, S => mult_21_C245_n655);
   mult_21_C245_U490 : ADFULD1 port map( A => mult_21_C245_n670, B => 
                           mult_21_C245_n659, CI => mult_21_C245_n657, CO => 
                           mult_21_C245_n652, S => mult_21_C245_n653);
   mult_21_C245_U489 : ADFULD1 port map( A => mult_21_C245_n668, B => 
                           mult_21_C245_n655, CI => mult_21_C245_n653, CO => 
                           mult_21_C245_n650, S => mult_21_C245_n651);
   mult_21_C245_U487 : ADFULD1 port map( A => mult_21_C245_n1200, B => 
                           mult_21_C245_n1350, CI => mult_21_C245_n1320, CO => 
                           mult_21_C245_n646, S => mult_21_C245_n647);
   mult_21_C245_U486 : ADFULD1 port map( A => mult_21_C245_n1166, B => 
                           mult_21_C245_n1266, CI => mult_21_C245_n1220, CO => 
                           mult_21_C245_n644, S => mult_21_C245_n645);
   mult_21_C245_U485 : ADFULD1 port map( A => mult_21_C245_n1182, B => 
                           mult_21_C245_n1292, CI => mult_21_C245_n1242, CO => 
                           mult_21_C245_n642, S => mult_21_C245_n643);
   mult_21_C245_U484 : ADFULD1 port map( A => mult_21_C245_n649, B => 
                           mult_21_C245_n664, CI => mult_21_C245_n662, CO => 
                           mult_21_C245_n640, S => mult_21_C245_n641);
   mult_21_C245_U483 : ADFULD1 port map( A => mult_21_C245_n647, B => 
                           mult_21_C245_n660, CI => mult_21_C245_n643, CO => 
                           mult_21_C245_n638, S => mult_21_C245_n639);
   mult_21_C245_U482 : ADFULD1 port map( A => mult_21_C245_n658, B => 
                           mult_21_C245_n645, CI => mult_21_C245_n656, CO => 
                           mult_21_C245_n636, S => mult_21_C245_n637);
   mult_21_C245_U481 : ADFULD1 port map( A => mult_21_C245_n639, B => 
                           mult_21_C245_n641, CI => mult_21_C245_n654, CO => 
                           mult_21_C245_n634, S => mult_21_C245_n635);
   mult_21_C245_U480 : ADFULD1 port map( A => mult_21_C245_n652, B => 
                           mult_21_C245_n637, CI => mult_21_C245_n635, CO => 
                           mult_21_C245_n632, S => mult_21_C245_n633);
   mult_21_C245_U478 : ADFULD1 port map( A => mult_21_C245_n1151, B => 
                           mult_21_C245_n1199, CI => mult_21_C245_n1219, CO => 
                           mult_21_C245_n628, S => mult_21_C245_n629);
   mult_21_C245_U477 : ADFULD1 port map( A => mult_21_C245_n1291, B => 
                           mult_21_C245_n1181, CI => mult_21_C245_n1165, CO => 
                           mult_21_C245_n626, S => mult_21_C245_n627);
   mult_21_C245_U476 : ADFULD1 port map( A => mult_21_C245_n1241, B => 
                           mult_21_C245_n1265, CI => mult_21_C245_n648, CO => 
                           mult_21_C245_n624, S => mult_21_C245_n625);
   mult_21_C245_U475 : ADFULD1 port map( A => mult_21_C245_n646, B => 
                           mult_21_C245_n631, CI => mult_21_C245_n642, CO => 
                           mult_21_C245_n622, S => mult_21_C245_n623);
   mult_21_C245_U474 : ADFULD1 port map( A => mult_21_C245_n627, B => 
                           mult_21_C245_n644, CI => mult_21_C245_n629, CO => 
                           mult_21_C245_n620, S => mult_21_C245_n621);
   mult_21_C245_U473 : ADFULD1 port map( A => mult_21_C245_n640, B => 
                           mult_21_C245_n625, CI => mult_21_C245_n638, CO => 
                           mult_21_C245_n618, S => mult_21_C245_n619);
   mult_21_C245_U472 : ADFULD1 port map( A => mult_21_C245_n621, B => 
                           mult_21_C245_n623, CI => mult_21_C245_n636, CO => 
                           mult_21_C245_n616, S => mult_21_C245_n617);
   mult_21_C245_U471 : ADFULD1 port map( A => mult_21_C245_n634, B => 
                           mult_21_C245_n619, CI => mult_21_C245_n617, CO => 
                           mult_21_C245_n614, S => mult_21_C245_n615);
   mult_21_C245_U469 : ADFULD1 port map( A => mult_21_C245_n1164, B => 
                           mult_21_C245_n1348, CI => mult_21_C245_n1318, CO => 
                           mult_21_C245_n610, S => mult_21_C245_n611);
   mult_21_C245_U468 : ADFULD1 port map( A => mult_21_C245_n1290, B => 
                           mult_21_C245_n1198, CI => mult_21_C245_n1218, CO => 
                           mult_21_C245_n608, S => mult_21_C245_n609);
   mult_21_C245_U467 : ADFULD1 port map( A => mult_21_C245_n1150, B => 
                           mult_21_C245_n1264, CI => mult_21_C245_n1180, CO => 
                           mult_21_C245_n606, S => mult_21_C245_n607);
   mult_21_C245_U466 : ADFULD1 port map( A => mult_21_C245_n630, B => 
                           mult_21_C245_n1240, CI => mult_21_C245_n613, CO => 
                           mult_21_C245_n604, S => mult_21_C245_n605);
   mult_21_C245_U465 : ADFULD1 port map( A => mult_21_C245_n626, B => 
                           mult_21_C245_n628, CI => mult_21_C245_n624, CO => 
                           mult_21_C245_n602, S => mult_21_C245_n603);
   mult_21_C245_U464 : ADFULD1 port map( A => mult_21_C245_n609, B => 
                           mult_21_C245_n611, CI => mult_21_C245_n607, CO => 
                           mult_21_C245_n600, S => mult_21_C245_n601);
   mult_21_C245_U463 : ADFULD1 port map( A => mult_21_C245_n622, B => 
                           mult_21_C245_n605, CI => mult_21_C245_n620, CO => 
                           mult_21_C245_n598, S => mult_21_C245_n599);
   mult_21_C245_U462 : ADFULD1 port map( A => mult_21_C245_n601, B => 
                           mult_21_C245_n603, CI => mult_21_C245_n618, CO => 
                           mult_21_C245_n596, S => mult_21_C245_n597);
   mult_21_C245_U461 : ADFULD1 port map( A => mult_21_C245_n616, B => 
                           mult_21_C245_n599, CI => mult_21_C245_n597, CO => 
                           mult_21_C245_n594, S => mult_21_C245_n595);
   mult_21_C245_U459 : ADFULD1 port map( A => mult_21_C245_n1289, B => 
                           mult_21_C245_n1179, CI => mult_21_C245_n1217, CO => 
                           mult_21_C245_n590, S => mult_21_C245_n591);
   mult_21_C245_U458 : ADFULD1 port map( A => mult_21_C245_n1263, B => 
                           mult_21_C245_n1149, CI => mult_21_C245_n1137, CO => 
                           mult_21_C245_n588, S => mult_21_C245_n589);
   mult_21_C245_U457 : ADFULD1 port map( A => mult_21_C245_n1163, B => 
                           mult_21_C245_n1239, CI => mult_21_C245_n1197, CO => 
                           mult_21_C245_n586, S => mult_21_C245_n587);
   mult_21_C245_U456 : ADFULD1 port map( A => mult_21_C245_n593, B => 
                           mult_21_C245_n612, CI => mult_21_C245_n610, CO => 
                           mult_21_C245_n584, S => mult_21_C245_n585);
   mult_21_C245_U455 : ADFULD1 port map( A => mult_21_C245_n606, B => 
                           mult_21_C245_n608, CI => mult_21_C245_n587, CO => 
                           mult_21_C245_n582, S => mult_21_C245_n583);
   mult_21_C245_U454 : ADFULD1 port map( A => mult_21_C245_n591, B => 
                           mult_21_C245_n589, CI => mult_21_C245_n604, CO => 
                           mult_21_C245_n580, S => mult_21_C245_n581);
   mult_21_C245_U453 : ADFULD1 port map( A => mult_21_C245_n585, B => 
                           mult_21_C245_n602, CI => mult_21_C245_n600, CO => 
                           mult_21_C245_n578, S => mult_21_C245_n579);
   mult_21_C245_U452 : ADFULD1 port map( A => mult_21_C245_n581, B => 
                           mult_21_C245_n583, CI => mult_21_C245_n598, CO => 
                           mult_21_C245_n576, S => mult_21_C245_n577);
   mult_21_C245_U451 : ADFULD1 port map( A => mult_21_C245_n596, B => 
                           mult_21_C245_n579, CI => mult_21_C245_n577, CO => 
                           mult_21_C245_n574, S => mult_21_C245_n575);
   mult_21_C245_U449 : ADFULD1 port map( A => mult_21_C245_n1136, B => 
                           mult_21_C245_n1346, CI => mult_21_C245_n1316, CO => 
                           mult_21_C245_n570, S => mult_21_C245_n571);
   mult_21_C245_U448 : ADFULD1 port map( A => mult_21_C245_n1288, B => 
                           mult_21_C245_n1178, CI => mult_21_C245_n1216, CO => 
                           mult_21_C245_n568, S => mult_21_C245_n569);
   mult_21_C245_U447 : ADFULD1 port map( A => mult_21_C245_n1148, B => 
                           mult_21_C245_n1262, CI => mult_21_C245_n1162, CO => 
                           mult_21_C245_n566, S => mult_21_C245_n567);
   mult_21_C245_U446 : ADFULD1 port map( A => mult_21_C245_n1196, B => 
                           mult_21_C245_n1238, CI => mult_21_C245_n592, CO => 
                           mult_21_C245_n564, S => mult_21_C245_n565);
   mult_21_C245_U445 : ADFULD1 port map( A => mult_21_C245_n590, B => 
                           mult_21_C245_n573, CI => mult_21_C245_n588, CO => 
                           mult_21_C245_n562, S => mult_21_C245_n563);
   mult_21_C245_U444 : ADFULD1 port map( A => mult_21_C245_n571, B => 
                           mult_21_C245_n586, CI => mult_21_C245_n567, CO => 
                           mult_21_C245_n560, S => mult_21_C245_n561);
   mult_21_C245_U443 : ADFULD1 port map( A => mult_21_C245_n565, B => 
                           mult_21_C245_n569, CI => mult_21_C245_n584, CO => 
                           mult_21_C245_n558, S => mult_21_C245_n559);
   mult_21_C245_U442 : ADFULD1 port map( A => mult_21_C245_n563, B => 
                           mult_21_C245_n582, CI => mult_21_C245_n580, CO => 
                           mult_21_C245_n556, S => mult_21_C245_n557);
   mult_21_C245_U441 : ADFULD1 port map( A => mult_21_C245_n559, B => 
                           mult_21_C245_n561, CI => mult_21_C245_n578, CO => 
                           mult_21_C245_n554, S => mult_21_C245_n555);
   mult_21_C245_U440 : ADFULD1 port map( A => mult_21_C245_n576, B => 
                           mult_21_C245_n557, CI => mult_21_C245_n555, CO => 
                           mult_21_C245_n552, S => mult_21_C245_n553);
   mult_21_C245_U438 : ADFULD1 port map( A => mult_21_C245_n1125, B => 
                           mult_21_C245_n1177, CI => mult_21_C245_n1215, CO => 
                           mult_21_C245_n548, S => mult_21_C245_n549);
   mult_21_C245_U437 : ADFULD1 port map( A => mult_21_C245_n1287, B => 
                           mult_21_C245_n1161, CI => mult_21_C245_n1261, CO => 
                           mult_21_C245_n546, S => mult_21_C245_n547);
   mult_21_C245_U436 : ADFULD1 port map( A => mult_21_C245_n1135, B => 
                           mult_21_C245_n1237, CI => mult_21_C245_n1147, CO => 
                           mult_21_C245_n544, S => mult_21_C245_n545);
   mult_21_C245_U435 : ADFULD1 port map( A => mult_21_C245_n572, B => 
                           mult_21_C245_n1195, CI => mult_21_C245_n551, CO => 
                           mult_21_C245_n542, S => mult_21_C245_n543);
   mult_21_C245_U434 : ADFULD1 port map( A => mult_21_C245_n566, B => 
                           mult_21_C245_n570, CI => mult_21_C245_n568, CO => 
                           mult_21_C245_n540, S => mult_21_C245_n541);
   mult_21_C245_U433 : ADFULD1 port map( A => mult_21_C245_n549, B => 
                           mult_21_C245_n564, CI => mult_21_C245_n547, CO => 
                           mult_21_C245_n538, S => mult_21_C245_n539);
   mult_21_C245_U432 : ADFULD1 port map( A => mult_21_C245_n562, B => 
                           mult_21_C245_n545, CI => mult_21_C245_n543, CO => 
                           mult_21_C245_n536, S => mult_21_C245_n537);
   mult_21_C245_U431 : ADFULD1 port map( A => mult_21_C245_n541, B => 
                           mult_21_C245_n560, CI => mult_21_C245_n558, CO => 
                           mult_21_C245_n534, S => mult_21_C245_n535);
   mult_21_C245_U430 : ADFULD1 port map( A => mult_21_C245_n556, B => 
                           mult_21_C245_n539, CI => mult_21_C245_n537, CO => 
                           mult_21_C245_n532, S => mult_21_C245_n533);
   mult_21_C245_U429 : ADFULD1 port map( A => mult_21_C245_n554, B => 
                           mult_21_C245_n535, CI => mult_21_C245_n533, CO => 
                           mult_21_C245_n530, S => mult_21_C245_n531);
   mult_21_C245_U427 : ADFULD1 port map( A => mult_21_C245_n1146, B => 
                           mult_21_C245_n1344, CI => mult_21_C245_n1314, CO => 
                           mult_21_C245_n526, S => mult_21_C245_n527);
   mult_21_C245_U426 : ADFULD1 port map( A => mult_21_C245_n1124, B => 
                           mult_21_C245_n1176, CI => mult_21_C245_n1214, CO => 
                           mult_21_C245_n524, S => mult_21_C245_n525);
   mult_21_C245_U425 : ADFULD1 port map( A => mult_21_C245_n1134, B => 
                           mult_21_C245_n1286, CI => mult_21_C245_n1160, CO => 
                           mult_21_C245_n522, S => mult_21_C245_n523);
   mult_21_C245_U424 : ADFULD1 port map( A => mult_21_C245_n1194, B => 
                           mult_21_C245_n1260, CI => mult_21_C245_n1236, CO => 
                           mult_21_C245_n520, S => mult_21_C245_n521);
   mult_21_C245_U423 : ADFULD1 port map( A => mult_21_C245_n529, B => 
                           mult_21_C245_n550, CI => mult_21_C245_n548, CO => 
                           mult_21_C245_n518, S => mult_21_C245_n519);
   mult_21_C245_U422 : ADFULD1 port map( A => mult_21_C245_n544, B => 
                           mult_21_C245_n546, CI => mult_21_C245_n527, CO => 
                           mult_21_C245_n516, S => mult_21_C245_n517);
   mult_21_C245_U421 : ADFULD1 port map( A => mult_21_C245_n525, B => 
                           mult_21_C245_n521, CI => mult_21_C245_n523, CO => 
                           mult_21_C245_n514, S => mult_21_C245_n515);
   mult_21_C245_U420 : ADFULD1 port map( A => mult_21_C245_n540, B => 
                           mult_21_C245_n542, CI => mult_21_C245_n519, CO => 
                           mult_21_C245_n512, S => mult_21_C245_n513);
   mult_21_C245_U419 : ADFULD1 port map( A => mult_21_C245_n517, B => 
                           mult_21_C245_n538, CI => mult_21_C245_n515, CO => 
                           mult_21_C245_n510, S => mult_21_C245_n511);
   mult_21_C245_U418 : ADFULD1 port map( A => mult_21_C245_n513, B => 
                           mult_21_C245_n536, CI => mult_21_C245_n534, CO => 
                           mult_21_C245_n508, S => mult_21_C245_n509);
   mult_21_C245_U417 : ADFULD1 port map( A => mult_21_C245_n532, B => 
                           mult_21_C245_n511, CI => mult_21_C245_n509, CO => 
                           mult_21_C245_n506, S => mult_21_C245_n507);
   mult_21_C245_U415 : ADFULD1 port map( A => mult_21_C245_n1115, B => 
                           mult_21_C245_n1175, CI => mult_21_C245_n1213, CO => 
                           mult_21_C245_n502, S => mult_21_C245_n503);
   mult_21_C245_U414 : ADFULD1 port map( A => mult_21_C245_n1123, B => 
                           mult_21_C245_n1145, CI => mult_21_C245_n1133, CO => 
                           mult_21_C245_n500, S => mult_21_C245_n501);
   mult_21_C245_U413 : ADFULD1 port map( A => mult_21_C245_n1159, B => 
                           mult_21_C245_n1285, CI => mult_21_C245_n1193, CO => 
                           mult_21_C245_n498, S => mult_21_C245_n499);
   mult_21_C245_U412 : ADFULD1 port map( A => mult_21_C245_n1235, B => 
                           mult_21_C245_n1259, CI => mult_21_C245_n528, CO => 
                           mult_21_C245_n496, S => mult_21_C245_n497);
   mult_21_C245_U411 : ADFULD1 port map( A => mult_21_C245_n526, B => 
                           mult_21_C245_n505, CI => mult_21_C245_n520, CO => 
                           mult_21_C245_n494, S => mult_21_C245_n495);
   mult_21_C245_U410 : ADFULD1 port map( A => mult_21_C245_n522, B => 
                           mult_21_C245_n524, CI => mult_21_C245_n499, CO => 
                           mult_21_C245_n492, S => mult_21_C245_n493);
   mult_21_C245_U409 : ADFULD1 port map( A => mult_21_C245_n501, B => 
                           mult_21_C245_n503, CI => mult_21_C245_n497, CO => 
                           mult_21_C245_n490, S => mult_21_C245_n491);
   mult_21_C245_U408 : ADFULD1 port map( A => mult_21_C245_n516, B => 
                           mult_21_C245_n518, CI => mult_21_C245_n495, CO => 
                           mult_21_C245_n488, S => mult_21_C245_n489);
   mult_21_C245_U407 : ADFULD1 port map( A => mult_21_C245_n493, B => 
                           mult_21_C245_n514, CI => mult_21_C245_n491, CO => 
                           mult_21_C245_n486, S => mult_21_C245_n487);
   mult_21_C245_U406 : ADFULD1 port map( A => mult_21_C245_n510, B => 
                           mult_21_C245_n512, CI => mult_21_C245_n489, CO => 
                           mult_21_C245_n484, S => mult_21_C245_n485);
   mult_21_C245_U405 : ADFULD1 port map( A => mult_21_C245_n508, B => 
                           mult_21_C245_n487, CI => mult_21_C245_n485, CO => 
                           mult_21_C245_n482, S => mult_21_C245_n483);
   mult_21_C245_U403 : ADFULD1 port map( A => mult_21_C245_n1114, B => 
                           mult_21_C245_n1342, CI => mult_21_C245_n1312, CO => 
                           mult_21_C245_n478, S => mult_21_C245_n479);
   mult_21_C245_U402 : ADFULD1 port map( A => mult_21_C245_n1284, B => 
                           mult_21_C245_n1174, CI => mult_21_C245_n1212, CO => 
                           mult_21_C245_n476, S => mult_21_C245_n477);
   mult_21_C245_U401 : ADFULD1 port map( A => mult_21_C245_n1258, B => 
                           mult_21_C245_n1132, CI => mult_21_C245_n1122, CO => 
                           mult_21_C245_n474, S => mult_21_C245_n475);
   mult_21_C245_U400 : ADFULD1 port map( A => mult_21_C245_n1144, B => 
                           mult_21_C245_n1234, CI => mult_21_C245_n1158, CO => 
                           mult_21_C245_n472, S => mult_21_C245_n473);
   mult_21_C245_U399 : ADFULD1 port map( A => mult_21_C245_n504, B => 
                           mult_21_C245_n1192, CI => mult_21_C245_n481, CO => 
                           mult_21_C245_n470, S => mult_21_C245_n471);
   mult_21_C245_U398 : ADFULD1 port map( A => mult_21_C245_n498, B => 
                           mult_21_C245_n502, CI => mult_21_C245_n496, CO => 
                           mult_21_C245_n468, S => mult_21_C245_n469);
   mult_21_C245_U397 : ADFULD1 port map( A => mult_21_C245_n479, B => 
                           mult_21_C245_n500, CI => mult_21_C245_n473, CO => 
                           mult_21_C245_n466, S => mult_21_C245_n467);
   mult_21_C245_U396 : ADFULD1 port map( A => mult_21_C245_n475, B => 
                           mult_21_C245_n477, CI => mult_21_C245_n471, CO => 
                           mult_21_C245_n464, S => mult_21_C245_n465);
   mult_21_C245_U395 : ADFULD1 port map( A => mult_21_C245_n492, B => 
                           mult_21_C245_n494, CI => mult_21_C245_n490, CO => 
                           mult_21_C245_n462, S => mult_21_C245_n463);
   mult_21_C245_U394 : ADFULD1 port map( A => mult_21_C245_n467, B => 
                           mult_21_C245_n469, CI => mult_21_C245_n465, CO => 
                           mult_21_C245_n460, S => mult_21_C245_n461);
   mult_21_C245_U393 : ADFULD1 port map( A => mult_21_C245_n486, B => 
                           mult_21_C245_n488, CI => mult_21_C245_n463, CO => 
                           mult_21_C245_n458, S => mult_21_C245_n459);
   mult_21_C245_U392 : ADFULD1 port map( A => mult_21_C245_n484, B => 
                           mult_21_C245_n461, CI => mult_21_C245_n459, CO => 
                           mult_21_C245_n456, S => mult_21_C245_n457);
   mult_21_C245_U390 : ADFULD1 port map( A => mult_21_C245_n1107, B => 
                           mult_21_C245_n1157, CI => mult_21_C245_n1211, CO => 
                           mult_21_C245_n452, S => mult_21_C245_n453);
   mult_21_C245_U389 : ADFULD1 port map( A => mult_21_C245_n1283, B => 
                           mult_21_C245_n1143, CI => mult_21_C245_n1257, CO => 
                           mult_21_C245_n450, S => mult_21_C245_n451);
   mult_21_C245_U388 : ADFULD1 port map( A => mult_21_C245_n1113, B => 
                           mult_21_C245_n1233, CI => mult_21_C245_n1121, CO => 
                           mult_21_C245_n448, S => mult_21_C245_n449);
   mult_21_C245_U387 : ADFULD1 port map( A => mult_21_C245_n1131, B => 
                           mult_21_C245_n1191, CI => mult_21_C245_n1173, CO => 
                           mult_21_C245_n446, S => mult_21_C245_n447);
   mult_21_C245_U386 : ADFULD1 port map( A => mult_21_C245_n455, B => 
                           mult_21_C245_n480, CI => mult_21_C245_n478, CO => 
                           mult_21_C245_n444, S => mult_21_C245_n445);
   mult_21_C245_U385 : ADFULD1 port map( A => mult_21_C245_n474, B => 
                           mult_21_C245_n472, CI => mult_21_C245_n476, CO => 
                           mult_21_C245_n442, S => mult_21_C245_n443);
   mult_21_C245_U384 : ADFULD1 port map( A => mult_21_C245_n453, B => 
                           mult_21_C245_n447, CI => mult_21_C245_n470, CO => 
                           mult_21_C245_n440, S => mult_21_C245_n441);
   mult_21_C245_U383 : ADFULD1 port map( A => mult_21_C245_n449, B => 
                           mult_21_C245_n451, CI => mult_21_C245_n468, CO => 
                           mult_21_C245_n438, S => mult_21_C245_n439);
   mult_21_C245_U382 : ADFULD1 port map( A => mult_21_C245_n466, B => 
                           mult_21_C245_n445, CI => mult_21_C245_n443, CO => 
                           mult_21_C245_n436, S => mult_21_C245_n437);
   mult_21_C245_U381 : ADFULD1 port map( A => mult_21_C245_n441, B => 
                           mult_21_C245_n464, CI => mult_21_C245_n462, CO => 
                           mult_21_C245_n434, S => mult_21_C245_n435);
   mult_21_C245_U380 : ADFULD1 port map( A => mult_21_C245_n437, B => 
                           mult_21_C245_n439, CI => mult_21_C245_n460, CO => 
                           mult_21_C245_n432, S => mult_21_C245_n433);
   mult_21_C245_U379 : ADFULD1 port map( A => mult_21_C245_n458, B => 
                           mult_21_C245_n435, CI => mult_21_C245_n433, CO => 
                           mult_21_C245_n430, S => mult_21_C245_n431);
   mult_21_C245_U377 : ADFULD1 port map( A => mult_21_C245_n1106, B => 
                           mult_21_C245_n1340, CI => mult_21_C245_n1310, CO => 
                           mult_21_C245_n426, S => mult_21_C245_n427);
   mult_21_C245_U376 : ADFULD1 port map( A => mult_21_C245_n1282, B => 
                           mult_21_C245_n1156, CI => mult_21_C245_n1210, CO => 
                           mult_21_C245_n424, S => mult_21_C245_n425);
   mult_21_C245_U375 : ADFULD1 port map( A => mult_21_C245_n1112, B => 
                           mult_21_C245_n1130, CI => mult_21_C245_n1120, CO => 
                           mult_21_C245_n422, S => mult_21_C245_n423);
   mult_21_C245_U374 : ADFULD1 port map( A => mult_21_C245_n1142, B => 
                           mult_21_C245_n1256, CI => mult_21_C245_n1172, CO => 
                           mult_21_C245_n420, S => mult_21_C245_n421);
   mult_21_C245_U373 : ADFULD1 port map( A => mult_21_C245_n1232, B => 
                           mult_21_C245_n1190, CI => mult_21_C245_n454, CO => 
                           mult_21_C245_n418, S => mult_21_C245_n419);
   mult_21_C245_U372 : ADFULD1 port map( A => mult_21_C245_n452, B => 
                           mult_21_C245_n429, CI => mult_21_C245_n450, CO => 
                           mult_21_C245_n416, S => mult_21_C245_n417);
   mult_21_C245_U371 : ADFULD1 port map( A => mult_21_C245_n448, B => 
                           mult_21_C245_n446, CI => mult_21_C245_n427, CO => 
                           mult_21_C245_n414, S => mult_21_C245_n415);
   mult_21_C245_U370 : ADFULD1 port map( A => mult_21_C245_n421, B => 
                           mult_21_C245_n423, CI => mult_21_C245_n425, CO => 
                           mult_21_C245_n412, S => mult_21_C245_n413);
   mult_21_C245_U369 : ADFULD1 port map( A => mult_21_C245_n444, B => 
                           mult_21_C245_n419, CI => mult_21_C245_n442, CO => 
                           mult_21_C245_n410, S => mult_21_C245_n411);
   mult_21_C245_U368 : ADFULD1 port map( A => mult_21_C245_n440, B => 
                           mult_21_C245_n417, CI => mult_21_C245_n415, CO => 
                           mult_21_C245_n408, S => mult_21_C245_n409);
   mult_21_C245_U367 : ADFULD1 port map( A => mult_21_C245_n438, B => 
                           mult_21_C245_n413, CI => mult_21_C245_n411, CO => 
                           mult_21_C245_n406, S => mult_21_C245_n407);
   mult_21_C245_U366 : ADFULD1 port map( A => mult_21_C245_n409, B => 
                           mult_21_C245_n436, CI => mult_21_C245_n434, CO => 
                           mult_21_C245_n404, S => mult_21_C245_n405);
   mult_21_C245_U365 : ADFULD1 port map( A => mult_21_C245_n432, B => 
                           mult_21_C245_n407, CI => mult_21_C245_n405, CO => 
                           mult_21_C245_n402, S => mult_21_C245_n403);
   mult_21_C245_U363 : ADFULD1 port map( A => mult_21_C245_n1281, B => 
                           mult_21_C245_n1155, CI => mult_21_C245_n1209, CO => 
                           mult_21_C245_n398, S => mult_21_C245_n399);
   mult_21_C245_U362 : ADFULD1 port map( A => mult_21_C245_n1255, B => 
                           mult_21_C245_n1119, CI => mult_21_C245_n1101, CO => 
                           mult_21_C245_n396, S => mult_21_C245_n397);
   mult_21_C245_U361 : ADFULD1 port map( A => mult_21_C245_n1231, B => 
                           mult_21_C245_n1111, CI => mult_21_C245_n1105, CO => 
                           mult_21_C245_n394, S => mult_21_C245_n395);
   mult_21_C245_U360 : ADFULD1 port map( A => mult_21_C245_n1129, B => 
                           mult_21_C245_n1189, CI => mult_21_C245_n1141, CO => 
                           mult_21_C245_n392, S => mult_21_C245_n393);
   mult_21_C245_U359 : ADFULD1 port map( A => mult_21_C245_n428, B => 
                           mult_21_C245_n1171, CI => mult_21_C245_n401, CO => 
                           mult_21_C245_n390, S => mult_21_C245_n391);
   mult_21_C245_U358 : ADFULD1 port map( A => mult_21_C245_n424, B => 
                           mult_21_C245_n426, CI => mult_21_C245_n420, CO => 
                           mult_21_C245_n388, S => mult_21_C245_n389);
   mult_21_C245_U357 : ADFULD1 port map( A => mult_21_C245_n418, B => 
                           mult_21_C245_n422, CI => mult_21_C245_n393, CO => 
                           mult_21_C245_n386, S => mult_21_C245_n387);
   mult_21_C245_U356 : ADFULD1 port map( A => mult_21_C245_n395, B => 
                           mult_21_C245_n397, CI => mult_21_C245_n399, CO => 
                           mult_21_C245_n384, S => mult_21_C245_n385);
   mult_21_C245_U355 : ADFULD1 port map( A => mult_21_C245_n391, B => 
                           mult_21_C245_n416, CI => mult_21_C245_n414, CO => 
                           mult_21_C245_n382, S => mult_21_C245_n383);
   mult_21_C245_U354 : ADFULD1 port map( A => mult_21_C245_n412, B => 
                           mult_21_C245_n389, CI => mult_21_C245_n387, CO => 
                           mult_21_C245_n380, S => mult_21_C245_n381);
   mult_21_C245_U353 : ADFULD1 port map( A => mult_21_C245_n410, B => 
                           mult_21_C245_n385, CI => mult_21_C245_n383, CO => 
                           mult_21_C245_n378, S => mult_21_C245_n379);
   mult_21_C245_U352 : ADFULD1 port map( A => mult_21_C245_n381, B => 
                           mult_21_C245_n408, CI => mult_21_C245_n406, CO => 
                           mult_21_C245_n376, S => mult_21_C245_n377);
   mult_21_C245_U351 : ADFULD1 port map( A => mult_21_C245_n404, B => 
                           mult_21_C245_n379, CI => mult_21_C245_n377, CO => 
                           mult_21_C245_n374, S => mult_21_C245_n375);
   mult_21_C245_U349 : ADFULD1 port map( A => mult_21_C245_n1100, B => 
                           mult_21_C245_n1338, CI => mult_21_C245_n1308, CO => 
                           mult_21_C245_n370, S => mult_21_C245_n371);
   mult_21_C245_U348 : ADFULD1 port map( A => mult_21_C245_n1280, B => 
                           mult_21_C245_n1154, CI => mult_21_C245_n1208, CO => 
                           mult_21_C245_n368, S => mult_21_C245_n369);
   mult_21_C245_U347 : ADFULD1 port map( A => mult_21_C245_n1254, B => 
                           mult_21_C245_n1128, CI => mult_21_C245_n1230, CO => 
                           mult_21_C245_n366, S => mult_21_C245_n367);
   mult_21_C245_U346 : ADFULD1 port map( A => mult_21_C245_n1104, B => 
                           mult_21_C245_n1188, CI => mult_21_C245_n1110, CO => 
                           mult_21_C245_n364, S => mult_21_C245_n365);
   mult_21_C245_U345 : ADFULD1 port map( A => mult_21_C245_n1170, B => 
                           mult_21_C245_n1118, CI => mult_21_C245_n1140, CO => 
                           mult_21_C245_n362, S => mult_21_C245_n363);
   mult_21_C245_U344 : ADFULD1 port map( A => mult_21_C245_n373, B => 
                           mult_21_C245_n400, CI => mult_21_C245_n392, CO => 
                           mult_21_C245_n360, S => mult_21_C245_n361);
   mult_21_C245_U343 : ADFULD1 port map( A => mult_21_C245_n398, B => 
                           mult_21_C245_n394, CI => mult_21_C245_n396, CO => 
                           mult_21_C245_n358, S => mult_21_C245_n359);
   mult_21_C245_U342 : ADFULD1 port map( A => mult_21_C245_n369, B => 
                           mult_21_C245_n371, CI => mult_21_C245_n367, CO => 
                           mult_21_C245_n356, S => mult_21_C245_n357);
   mult_21_C245_U341 : ADFULD1 port map( A => mult_21_C245_n365, B => 
                           mult_21_C245_n363, CI => mult_21_C245_n390, CO => 
                           mult_21_C245_n354, S => mult_21_C245_n355);
   mult_21_C245_U340 : ADFULD1 port map( A => mult_21_C245_n361, B => 
                           mult_21_C245_n388, CI => mult_21_C245_n386, CO => 
                           mult_21_C245_n352, S => mult_21_C245_n353);
   mult_21_C245_U339 : ADFULD1 port map( A => mult_21_C245_n359, B => 
                           mult_21_C245_n384, CI => mult_21_C245_n357, CO => 
                           mult_21_C245_n350, S => mult_21_C245_n351);
   mult_21_C245_U338 : ADFULD1 port map( A => mult_21_C245_n382, B => 
                           mult_21_C245_n355, CI => mult_21_C245_n380, CO => 
                           mult_21_C245_n348, S => mult_21_C245_n349);
   mult_21_C245_U337 : ADFULD1 port map( A => mult_21_C245_n351, B => 
                           mult_21_C245_n353, CI => mult_21_C245_n378, CO => 
                           mult_21_C245_n346, S => mult_21_C245_n347);
   mult_21_C245_U336 : ADFULD1 port map( A => mult_21_C245_n376, B => 
                           mult_21_C245_n349, CI => mult_21_C245_n347, CO => 
                           mult_21_C245_n344, S => mult_21_C245_n345);
   mult_21_C245_U334 : EXOR3D1 port map( A1 => mult_21_C245_n1097, A2 => 
                           mult_21_C245_n1279, A3 => mult_21_C245_n1207, Z => 
                           mult_21_C245_n342);
   mult_21_C245_U333 : EXOR3D1 port map( A1 => mult_21_C245_n1253, A2 => 
                           mult_21_C245_n1127, A3 => mult_21_C245_n1099, Z => 
                           mult_21_C245_n341);
   mult_21_C245_U332 : EXOR3D1 port map( A1 => mult_21_C245_n1103, A2 => 
                           mult_21_C245_n1117, A3 => mult_21_C245_n1109, Z => 
                           mult_21_C245_n340);
   mult_21_C245_U331 : EXOR3D1 port map( A1 => mult_21_C245_n1139, A2 => 
                           mult_21_C245_n1229, A3 => mult_21_C245_n1153, Z => 
                           mult_21_C245_n339);
   mult_21_C245_U330 : EXOR3D1 port map( A1 => mult_21_C245_n1187, A2 => 
                           mult_21_C245_n1169, A3 => mult_21_C245_n372, Z => 
                           mult_21_C245_n338);
   mult_21_C245_U329 : EXOR3D1 port map( A1 => mult_21_C245_n368, A2 => 
                           mult_21_C245_n370, A3 => mult_21_C245_n364, Z => 
                           mult_21_C245_n337);
   mult_21_C245_U328 : EXOR3D1 port map( A1 => mult_21_C245_n366, A2 => 
                           mult_21_C245_n343, A3 => mult_21_C245_n362, Z => 
                           mult_21_C245_n336);
   mult_21_C245_U327 : EXOR3D1 port map( A1 => mult_21_C245_n342, A2 => 
                           mult_21_C245_n338, A3 => mult_21_C245_n341, Z => 
                           mult_21_C245_n335);
   mult_21_C245_U326 : EXOR3D1 port map( A1 => mult_21_C245_n339, A2 => 
                           mult_21_C245_n340, A3 => mult_21_C245_n360, Z => 
                           mult_21_C245_n334);
   mult_21_C245_U325 : EXOR3D1 port map( A1 => mult_21_C245_n337, A2 => 
                           mult_21_C245_n358, A3 => mult_21_C245_n336, Z => 
                           mult_21_C245_n333);
   mult_21_C245_U324 : EXOR3D1 port map( A1 => mult_21_C245_n354, A2 => 
                           mult_21_C245_n356, A3 => mult_21_C245_n335, Z => 
                           mult_21_C245_n332);
   mult_21_C245_U323 : EXOR3D1 port map( A1 => mult_21_C245_n352, A2 => 
                           mult_21_C245_n334, A3 => mult_21_C245_n333, Z => 
                           mult_21_C245_n331);
   mult_21_C245_U322 : EXOR3D1 port map( A1 => mult_21_C245_n332, A2 => 
                           mult_21_C245_n350, A3 => mult_21_C245_n348, Z => 
                           mult_21_C245_n330);
   mult_21_C245_U321 : EXOR3D1 port map( A1 => mult_21_C245_n346, A2 => 
                           mult_21_C245_n331, A3 => mult_21_C245_n330, Z => 
                           mult_21_C245_n329);
   mult_21_C245_U313 : EXOR2D1 port map( A1 => mult_21_C245_n303, A2 => 
                           mult_21_C245_n305, Z => N3298);
   mult_21_C245_U305 : EXNOR2D1 port map( A1 => mult_21_C245_n176, A2 => 
                           mult_21_C245_n302, Z => N3299);
   mult_21_C245_U300 : OAI21D1 port map( A1 => mult_21_C245_n297, A2 => 
                           mult_21_C245_n295, B => mult_21_C245_n296, Z => 
                           mult_21_C245_n294);
   mult_21_C245_U299 : EXOR2D1 port map( A1 => mult_21_C245_n297, A2 => 
                           mult_21_C245_n175, Z => N3300);
   mult_21_C245_U291 : EXNOR2D1 port map( A1 => mult_21_C245_n174, A2 => 
                           mult_21_C245_n294, Z => N3301);
   mult_21_C245_U286 : OAI21D1 port map( A1 => mult_21_C245_n289, A2 => 
                           mult_21_C245_n287, B => mult_21_C245_n288, Z => 
                           mult_21_C245_n286);
   mult_21_C245_U284 : EXOR2D1 port map( A1 => mult_21_C245_n173, A2 => 
                           mult_21_C245_n289, Z => N3302);
   mult_21_C245_U279 : OAI21D1 port map( A1 => mult_21_C245_n285, A2 => 
                           mult_21_C245_n283, B => mult_21_C245_n284, Z => 
                           mult_21_C245_n282);
   mult_21_C245_U278 : EXOR2D1 port map( A1 => mult_21_C245_n172, A2 => 
                           mult_21_C245_n285, Z => N3303);
   mult_21_C245_U273 : OAI21D1 port map( A1 => mult_21_C245_n280, A2 => 
                           mult_21_C245_n284, B => mult_21_C245_n281, Z => 
                           mult_21_C245_n279);
   mult_21_C245_U271 : AOI21D1 port map( A1 => mult_21_C245_n278, A2 => 
                           mult_21_C245_n286, B => mult_21_C245_n279, Z => 
                           mult_21_C245_n277);
   mult_21_C245_U269 : EXNOR2D1 port map( A1 => mult_21_C245_n282, A2 => 
                           mult_21_C245_n171, Z => N3304);
   mult_21_C245_U262 : AOI21D1 port map( A1 => mult_21_C245_n276, A2 => 
                           mult_21_C245_n1527, B => mult_21_C245_n273, Z => 
                           mult_21_C245_n271);
   mult_21_C245_U261 : EXNOR2D1 port map( A1 => mult_21_C245_n276, A2 => 
                           mult_21_C245_n170, Z => N3305);
   mult_21_C245_U254 : AOI21D1 port map( A1 => mult_21_C245_n1524, A2 => 
                           mult_21_C245_n273, B => mult_21_C245_n268, Z => 
                           mult_21_C245_n266);
   mult_21_C245_U252 : OAI21D1 port map( A1 => mult_21_C245_n265, A2 => 
                           mult_21_C245_n277, B => mult_21_C245_n266, Z => 
                           mult_21_C245_n264);
   mult_21_C245_U250 : EXOR2D1 port map( A1 => mult_21_C245_n271, A2 => 
                           mult_21_C245_n169, Z => N3306);
   mult_21_C245_U245 : OAI21D1 port map( A1 => mult_21_C245_n263, A2 => 
                           mult_21_C245_n261, B => mult_21_C245_n262, Z => 
                           mult_21_C245_n260);
   mult_21_C245_U244 : EXOR2D1 port map( A1 => mult_21_C245_n263, A2 => 
                           mult_21_C245_n168, Z => N3307);
   mult_21_C245_U239 : OAI21D1 port map( A1 => mult_21_C245_n258, A2 => 
                           mult_21_C245_n262, B => mult_21_C245_n259, Z => 
                           mult_21_C245_n257);
   mult_21_C245_U237 : AOI21D1 port map( A1 => mult_21_C245_n256, A2 => 
                           mult_21_C245_n264, B => mult_21_C245_n257, Z => 
                           mult_21_C245_n255);
   mult_21_C245_U235 : EXNOR2D1 port map( A1 => mult_21_C245_n260, A2 => 
                           mult_21_C245_n167, Z => N3308);
   mult_21_C245_U228 : AOI21D1 port map( A1 => mult_21_C245_n254, A2 => 
                           mult_21_C245_n1529, B => mult_21_C245_n251, Z => 
                           mult_21_C245_n249);
   mult_21_C245_U227 : EXNOR2D1 port map( A1 => mult_21_C245_n254, A2 => 
                           mult_21_C245_n166, Z => N3309);
   mult_21_C245_U220 : AOI21D1 port map( A1 => mult_21_C245_n1530, A2 => 
                           mult_21_C245_n251, B => mult_21_C245_n246, Z => 
                           mult_21_C245_n244);
   mult_21_C245_U218 : OAI21D1 port map( A1 => mult_21_C245_n255, A2 => 
                           mult_21_C245_n243, B => mult_21_C245_n244, Z => 
                           mult_21_C245_n242);
   mult_21_C245_U216 : EXOR2D1 port map( A1 => mult_21_C245_n249, A2 => 
                           mult_21_C245_n165, Z => N3310);
   mult_21_C245_U211 : OAI21D1 port map( A1 => mult_21_C245_n241, A2 => 
                           mult_21_C245_n239, B => mult_21_C245_n240, Z => 
                           mult_21_C245_n238);
   mult_21_C245_U210 : EXOR2D1 port map( A1 => mult_21_C245_n241, A2 => 
                           mult_21_C245_n164, Z => N3311);
   mult_21_C245_U205 : OAI21D1 port map( A1 => mult_21_C245_n236, A2 => 
                           mult_21_C245_n240, B => mult_21_C245_n237, Z => 
                           mult_21_C245_n235);
   mult_21_C245_U203 : AOI21D1 port map( A1 => mult_21_C245_n242, A2 => 
                           mult_21_C245_n234, B => mult_21_C245_n235, Z => 
                           mult_21_C245_n233);
   mult_21_C245_U201 : EXNOR2D1 port map( A1 => mult_21_C245_n238, A2 => 
                           mult_21_C245_n163, Z => N3312);
   mult_21_C245_U194 : AOI21D1 port map( A1 => mult_21_C245_n232, A2 => 
                           mult_21_C245_n313, B => mult_21_C245_n229, Z => 
                           mult_21_C245_n227);
   mult_21_C245_U193 : EXNOR2D1 port map( A1 => mult_21_C245_n232, A2 => 
                           mult_21_C245_n162, Z => N3313);
   mult_21_C245_U188 : OAI21D1 port map( A1 => mult_21_C245_n225, A2 => 
                           mult_21_C245_n231, B => mult_21_C245_n226, Z => 
                           mult_21_C245_n224);
   mult_21_C245_U186 : AOI21D1 port map( A1 => mult_21_C245_n232, A2 => 
                           mult_21_C245_n223, B => mult_21_C245_n224, Z => 
                           mult_21_C245_n222);
   mult_21_C245_U185 : EXOR2D1 port map( A1 => mult_21_C245_n227, A2 => 
                           mult_21_C245_n161, Z => N3314);
   mult_21_C245_U178 : AOI21D1 port map( A1 => mult_21_C245_n224, A2 => 
                           mult_21_C245_n1528, B => mult_21_C245_n219, Z => 
                           mult_21_C245_n217);
   mult_21_C245_U176 : OAI21D1 port map( A1 => mult_21_C245_n233, A2 => 
                           mult_21_C245_n216, B => mult_21_C245_n217, Z => 
                           mult_21_C245_n215);
   mult_21_C245_U174 : EXOR2D1 port map( A1 => mult_21_C245_n222, A2 => 
                           mult_21_C245_n160, Z => N3315);
   mult_21_C245_U165 : OAI21D1 port map( A1 => mult_21_C245_n214, A2 => 
                           mult_21_C245_n208, B => mult_21_C245_n209, Z => 
                           mult_21_C245_n207);
   mult_21_C245_U164 : EXOR2D1 port map( A1 => mult_21_C245_n214, A2 => 
                           mult_21_C245_n159, Z => N3316);
   mult_21_C245_U157 : AOI21D1 port map( A1 => mult_21_C245_n1525, A2 => 
                           mult_21_C245_n211, B => mult_21_C245_n204, Z => 
                           mult_21_C245_n202);
   mult_21_C245_U155 : OAI21D1 port map( A1 => mult_21_C245_n214, A2 => 
                           mult_21_C245_n201, B => mult_21_C245_n202, Z => 
                           mult_21_C245_n200);
   mult_21_C245_U154 : EXNOR2D1 port map( A1 => mult_21_C245_n207, A2 => 
                           mult_21_C245_n158, Z => N3317);
   mult_21_C245_U147 : AOI21D1 port map( A1 => mult_21_C245_n200, A2 => 
                           mult_21_C245_n1526, B => mult_21_C245_n197, Z => 
                           mult_21_C245_n195);
   mult_21_C245_U146 : EXNOR2D1 port map( A1 => mult_21_C245_n200, A2 => 
                           mult_21_C245_n157, Z => N3318);
   mult_21_C245_U137 : OAI21D1 port map( A1 => mult_21_C245_n202, A2 => 
                           mult_21_C245_n189, B => mult_21_C245_n190, Z => 
                           mult_21_C245_n188);
   mult_21_C245_U134 : EXOR2D1 port map( A1 => mult_21_C245_n195, A2 => 
                           mult_21_C245_n156, Z => N3319);
   mult_21_C245_U132 : ADFULD1 port map( A => mult_21_C245_n531, B => 
                           mult_21_C245_n552, CI => mult_21_C245_n1521, CO => 
                           mult_21_C245_n185, S => N3320);
   mult_21_C245_U131 : ADFULD1 port map( A => mult_21_C245_n507, B => 
                           mult_21_C245_n530, CI => mult_21_C245_n185, CO => 
                           mult_21_C245_n184, S => N3321);
   mult_21_C245_U130 : ADFULD1 port map( A => mult_21_C245_n483, B => 
                           mult_21_C245_n506, CI => mult_21_C245_n184, CO => 
                           mult_21_C245_n183, S => N3322);
   mult_21_C245_U129 : ADFULD1 port map( A => mult_21_C245_n457, B => 
                           mult_21_C245_n482, CI => mult_21_C245_n183, CO => 
                           mult_21_C245_n182, S => N3323);
   mult_21_C245_U128 : ADFULD1 port map( A => mult_21_C245_n431, B => 
                           mult_21_C245_n456, CI => mult_21_C245_n182, CO => 
                           mult_21_C245_n181, S => N3324);
   mult_21_C245_U127 : ADFULD1 port map( A => mult_21_C245_n403, B => 
                           mult_21_C245_n430, CI => mult_21_C245_n181, CO => 
                           mult_21_C245_n180, S => N3325);
   mult_21_C245_U126 : ADFULD1 port map( A => mult_21_C245_n375, B => 
                           mult_21_C245_n402, CI => mult_21_C245_n180, CO => 
                           mult_21_C245_n179, S => N3326);
   mult_21_C245_U125 : ADFULD1 port map( A => mult_21_C245_n345, B => 
                           mult_21_C245_n374, CI => mult_21_C245_n179, CO => 
                           mult_21_C245_n178, S => N3327);
   mult_21_C247_U1403 : INVD1 port map( A => N3040, Z => mult_21_C247_n1066);
   mult_21_C247_U1402 : AO21D1 port map( A1 => N3038, A2 => N3039, B => 
                           mult_21_C247_n1066, Z => mult_21_C247_n105);
   mult_21_C247_U1401 : INVD1 port map( A => N3038, Z => mult_21_C247_n1067);
   mult_21_C247_U1400 : AO21D1 port map( A1 => N3036, A2 => N3037, B => 
                           mult_21_C247_n1067, Z => mult_21_C247_n101);
   mult_21_C247_U1399 : INVD1 port map( A => N3036, Z => mult_21_C247_n1068);
   mult_21_C247_U1398 : AO21D1 port map( A1 => N3034, A2 => N3035, B => 
                           mult_21_C247_n1068, Z => mult_21_C247_n96);
   mult_21_C247_U1397 : ADHALFDL port map( A => mult_21_C247_n1309, B => 
                           mult_21_C247_n1339, CO => mult_21_C247_n400, S => 
                           mult_21_C247_n401);
   mult_21_C247_U1396 : AO21D1 port map( A1 => N3032, A2 => N3033, B => 
                           mult_21_C247_n1069, Z => mult_21_C247_n91);
   mult_21_C247_U1395 : INVD1 port map( A => N3034, Z => mult_21_C247_n1069);
   mult_21_C247_U1394 : ADHALFDL port map( A => mult_21_C247_n1311, B => 
                           mult_21_C247_n1341, CO => mult_21_C247_n454, S => 
                           mult_21_C247_n455);
   mult_21_C247_U1393 : OAI21D1 port map( A1 => N3032, A2 => N3033, B => 
                           mult_21_C247_n1069, Z => mult_21_C247_n89);
   mult_21_C247_U1392 : ADHALFDL port map( A => mult_21_C247_n1313, B => 
                           mult_21_C247_n1343, CO => mult_21_C247_n504, S => 
                           mult_21_C247_n505);
   mult_21_C247_U1391 : AO21D1 port map( A1 => N3030, A2 => N3031, B => 
                           mult_21_C247_n1070, Z => mult_21_C247_n86);
   mult_21_C247_U1390 : INVD1 port map( A => N3032, Z => mult_21_C247_n1070);
   mult_21_C247_U1389 : OAI21D1 port map( A1 => N3030, A2 => N3031, B => 
                           mult_21_C247_n1070, Z => mult_21_C247_n84);
   mult_21_C247_U1388 : AO21D1 port map( A1 => N3028, A2 => N3029, B => 
                           mult_21_C247_n1071, Z => mult_21_C247_n81);
   mult_21_C247_U1387 : INVD1 port map( A => N3030, Z => mult_21_C247_n1071);
   mult_21_C247_U1386 : OAI21D1 port map( A1 => N3028, A2 => N3029, B => 
                           mult_21_C247_n1071, Z => mult_21_C247_n79);
   mult_21_C247_U1385 : EXNOR2D1 port map( A1 => N3030, A2 => N3031, Z => 
                           mult_21_C247_n88);
   mult_21_C247_U1384 : AO21D1 port map( A1 => N3026, A2 => N3027, B => 
                           mult_21_C247_n1072, Z => mult_21_C247_n76);
   mult_21_C247_U1383 : OAI21D1 port map( A1 => N3018, A2 => N3019, B => 
                           mult_21_C247_n1076, Z => mult_21_C247_n42);
   mult_21_C247_U1382 : INVD1 port map( A => N3028, Z => mult_21_C247_n1072);
   mult_21_C247_U1381 : OAI21D1 port map( A1 => N3026, A2 => N3027, B => 
                           mult_21_C247_n1072, Z => mult_21_C247_n73);
   mult_21_C247_U1380 : INVD1 port map( A => N3020, Z => mult_21_C247_n1076);
   mult_21_C247_U1379 : AO21D1 port map( A1 => N3018, A2 => N3019, B => 
                           mult_21_C247_n1076, Z => mult_21_C247_n45);
   mult_21_C247_U1378 : OAI21D1 port map( A1 => N3024, A2 => N3025, B => 
                           mult_21_C247_n1073, Z => mult_21_C247_n66);
   mult_21_C247_U1377 : INVD1 port map( A => N3026, Z => mult_21_C247_n1073);
   mult_21_C247_U1376 : OAI21D1 port map( A1 => N3022, A2 => N3023, B => 
                           mult_21_C247_n1074, Z => mult_21_C247_n58);
   mult_21_C247_U1375 : INVD1 port map( A => N3024, Z => mult_21_C247_n1074);
   mult_21_C247_U1374 : AO21D1 port map( A1 => N3024, A2 => N3025, B => 
                           mult_21_C247_n1073, Z => mult_21_C247_n69);
   mult_21_C247_U1373 : AO21D1 port map( A1 => N3022, A2 => N3023, B => 
                           mult_21_C247_n1074, Z => mult_21_C247_n61);
   mult_21_C247_U1372 : OAI21D1 port map( A1 => N3020, A2 => N3021, B => 
                           mult_21_C247_n1075, Z => mult_21_C247_n50);
   mult_21_C247_U1371 : AO21D1 port map( A1 => N3016, A2 => N3017, B => 
                           mult_21_C247_n1077, Z => mult_21_C247_n38);
   mult_21_C247_U1370 : AO21D1 port map( A1 => N3012, A2 => N3013, B => 
                           mult_21_C247_n1079, Z => mult_21_C247_n22);
   mult_21_C247_U1369 : ADHALFDL port map( A => mult_21_C247_n1315, B => 
                           mult_21_C247_n1345, CO => mult_21_C247_n550, S => 
                           mult_21_C247_n551);
   mult_21_C247_U1368 : INVD1 port map( A => N3022, Z => mult_21_C247_n1075);
   mult_21_C247_U1367 : AO21D1 port map( A1 => N3020, A2 => N3021, B => 
                           mult_21_C247_n1075, Z => mult_21_C247_n53);
   mult_21_C247_U1366 : INVD1 port map( A => N3009, Z => mult_21_C247_n8);
   mult_21_C247_U1365 : EXNOR2D1 port map( A1 => N3028, A2 => N3029, Z => 
                           mult_21_C247_n83);
   mult_21_C247_U1364 : AO21D1 port map( A1 => N3014, A2 => N3015, B => 
                           mult_21_C247_n1078, Z => mult_21_C247_n30);
   mult_21_C247_U1363 : AO21D1 port map( A1 => N3010, A2 => N3011, B => 
                           mult_21_C247_n1080, Z => mult_21_C247_n14);
   mult_21_C247_U1362 : EXNOR2D1 port map( A1 => N3026, A2 => N3027, Z => 
                           mult_21_C247_n78);
   mult_21_C247_U1361 : EXNOR2D1 port map( A1 => N3018, A2 => N3019, Z => 
                           mult_21_C247_n48);
   mult_21_C247_U1360 : INVD1 port map( A => n288, Z => mult_21_C247_n1557);
   mult_21_C247_U1359 : INVD1 port map( A => N3014, Z => mult_21_C247_n1079);
   mult_21_C247_U1358 : INVD1 port map( A => n287, Z => mult_21_C247_n1550);
   mult_21_C247_U1357 : EXNOR2D1 port map( A1 => N3024, A2 => N3025, Z => 
                           mult_21_C247_n71);
   mult_21_C247_U1356 : EXNOR2D1 port map( A1 => N3022, A2 => N3023, Z => 
                           mult_21_C247_n63);
   mult_21_C247_U1355 : INVD1 port map( A => n286, Z => mult_21_C247_n1552);
   mult_21_C247_U1354 : INVD1 port map( A => N3018, Z => mult_21_C247_n1077);
   mult_21_C247_U1353 : INVD1 port map( A => n285, Z => mult_21_C247_n1544);
   mult_21_C247_U1352 : INVD1 port map( A => n284, Z => mult_21_C247_n1555);
   mult_21_C247_U1351 : INVD1 port map( A => N3010, Z => mult_21_C247_n6);
   mult_21_C247_U1350 : NAN2D1 port map( A1 => N3009, A2 => mult_21_C247_n6, Z 
                           => mult_21_C247_n3);
   mult_21_C247_U1349 : INVD1 port map( A => n282, Z => mult_21_C247_n1548);
   mult_21_C247_U1348 : INVD1 port map( A => n280, Z => mult_21_C247_n1546);
   mult_21_C247_U1347 : INVD1 port map( A => N3016, Z => mult_21_C247_n1078);
   mult_21_C247_U1346 : EXNOR2D1 port map( A1 => N3020, A2 => N3021, Z => 
                           mult_21_C247_n56);
   mult_21_C247_U1345 : INVD1 port map( A => N3012, Z => mult_21_C247_n1080);
   mult_21_C247_U1344 : OA21D1 port map( A1 => N3014, A2 => N3015, B => 
                           mult_21_C247_n1078, Z => mult_21_C247_n1537);
   mult_21_C247_U1343 : ADHALFDL port map( A => mult_21_C247_n1325, B => 
                           mult_21_C247_n1355, CO => mult_21_C247_n720, S => 
                           mult_21_C247_n721);
   mult_21_C247_U1342 : ADHALFDL port map( A => mult_21_C247_n1321, B => 
                           mult_21_C247_n1351, CO => mult_21_C247_n664, S => 
                           mult_21_C247_n665);
   mult_21_C247_U1341 : ADHALFDL port map( A => mult_21_C247_n1319, B => 
                           mult_21_C247_n1349, CO => mult_21_C247_n630, S => 
                           mult_21_C247_n631);
   mult_21_C247_U1340 : ADHALFDL port map( A => mult_21_C247_n1327, B => 
                           mult_21_C247_n1357, CO => mult_21_C247_n742, S => 
                           mult_21_C247_n743);
   mult_21_C247_U1339 : ADHALFDL port map( A => mult_21_C247_n1317, B => 
                           mult_21_C247_n1347, CO => mult_21_C247_n592, S => 
                           mult_21_C247_n593);
   mult_21_C247_U1338 : EXOR2D1 port map( A1 => N3016, A2 => N3017, Z => 
                           mult_21_C247_n1536);
   mult_21_C247_U1337 : EXOR2D1 port map( A1 => N3012, A2 => N3013, Z => 
                           mult_21_C247_n1535);
   mult_21_C247_U1336 : EXOR2D1 port map( A1 => N3014, A2 => N3015, Z => 
                           mult_21_C247_n1534);
   mult_21_C247_U1335 : ADHALFDL port map( A => mult_21_C247_n1323, B => 
                           mult_21_C247_n1353, CO => mult_21_C247_n694, S => 
                           mult_21_C247_n695);
   mult_21_C247_U1334 : EXOR2D1 port map( A1 => N3010, A2 => N3011, Z => 
                           mult_21_C247_n1533);
   mult_21_C247_U1333 : ADHALFDL port map( A => mult_21_C247_n1098, B => 
                           mult_21_C247_n1081, CO => mult_21_C247_n372, S => 
                           mult_21_C247_n373);
   mult_21_C247_U1332 : EXOR2D1 port map( A1 => mult_21_C247_n1307, A2 => 
                           mult_21_C247_n1337, Z => mult_21_C247_n343);
   mult_21_C247_U1331 : ADHALFDL port map( A => mult_21_C247_n1102, B => 
                           mult_21_C247_n1082, CO => mult_21_C247_n428, S => 
                           mult_21_C247_n429);
   mult_21_C247_U1330 : ADHALFDL port map( A => mult_21_C247_n1108, B => 
                           mult_21_C247_n1083, CO => mult_21_C247_n480, S => 
                           mult_21_C247_n481);
   mult_21_C247_U1329 : ADHALFDL port map( A => mult_21_C247_n1116, B => 
                           mult_21_C247_n1084, CO => mult_21_C247_n528, S => 
                           mult_21_C247_n529);
   mult_21_C247_U1328 : ADHALFDL port map( A => mult_21_C247_n1126, B => 
                           mult_21_C247_n1085, CO => mult_21_C247_n572, S => 
                           mult_21_C247_n573);
   mult_21_C247_U1327 : INVD1 port map( A => mult_21_C247_n1367, Z => 
                           mult_21_C247_n303);
   mult_21_C247_U1326 : ADHALFDL port map( A => mult_21_C247_n1138, B => 
                           mult_21_C247_n1086, CO => mult_21_C247_n612, S => 
                           mult_21_C247_n613);
   mult_21_C247_U1325 : ADHALFDL port map( A => mult_21_C247_n1186, B => 
                           mult_21_C247_n1089, CO => mult_21_C247_n708, S => 
                           mult_21_C247_n709);
   mult_21_C247_U1324 : ADHALFDL port map( A => mult_21_C247_n1228, B => 
                           mult_21_C247_n1091, CO => mult_21_C247_n752, S => 
                           mult_21_C247_n753);
   mult_21_C247_U1323 : ADHALFDL port map( A => mult_21_C247_n1152, B => 
                           mult_21_C247_n1087, CO => mult_21_C247_n648, S => 
                           mult_21_C247_n649);
   mult_21_C247_U1322 : ADHALFDL port map( A => mult_21_C247_n1168, B => 
                           mult_21_C247_n1088, CO => mult_21_C247_n680, S => 
                           mult_21_C247_n681);
   mult_21_C247_U1321 : ADHALFDL port map( A => mult_21_C247_n1206, B => 
                           mult_21_C247_n1090, CO => mult_21_C247_n732, S => 
                           mult_21_C247_n733);
   mult_21_C247_U1320 : INVD1 port map( A => mult_21_C247_n1550, Z => 
                           mult_21_C247_n1549);
   mult_21_C247_U1319 : INVD1 port map( A => mult_21_C247_n1557, Z => 
                           mult_21_C247_n1556);
   mult_21_C247_U1318 : INVD1 port map( A => mult_21_C247_n1552, Z => 
                           mult_21_C247_n1551);
   mult_21_C247_U1317 : INVD1 port map( A => mult_21_C247_n1555, Z => 
                           mult_21_C247_n1554);
   mult_21_C247_U1316 : INVD1 port map( A => mult_21_C247_n1544, Z => 
                           mult_21_C247_n1543);
   mult_21_C247_U1315 : INVD1 port map( A => mult_21_C247_n1546, Z => 
                           mult_21_C247_n1545);
   mult_21_C247_U1314 : INVD1 port map( A => mult_21_C247_n1555, Z => 
                           mult_21_C247_n1553);
   mult_21_C247_U1313 : INVD1 port map( A => mult_21_C247_n1548, Z => 
                           mult_21_C247_n1547);
   mult_21_C247_U1312 : INVD1 port map( A => mult_21_C247_n1537, Z => 
                           mult_21_C247_n1540);
   mult_21_C247_U1311 : ADHALFDL port map( A => mult_21_C247_n1306, B => 
                           mult_21_C247_n1094, CO => mult_21_C247_n788, S => 
                           mult_21_C247_n789);
   mult_21_C247_U1310 : INVD1 port map( A => mult_21_C247_n1536, Z => 
                           mult_21_C247_n1538);
   mult_21_C247_U1309 : ADHALFDL port map( A => mult_21_C247_n1333, B => 
                           mult_21_C247_n1363, CO => mult_21_C247_n784, S => 
                           mult_21_C247_n785);
   mult_21_C247_U1308 : ADHALFDL port map( A => mult_21_C247_n1252, B => 
                           mult_21_C247_n1092, CO => mult_21_C247_n768, S => 
                           mult_21_C247_n769);
   mult_21_C247_U1307 : INVD1 port map( A => mult_21_C247_n1534, Z => 
                           mult_21_C247_n1539);
   mult_21_C247_U1306 : ADHALFDL port map( A => mult_21_C247_n1331, B => 
                           mult_21_C247_n1361, CO => mult_21_C247_n774, S => 
                           mult_21_C247_n775);
   mult_21_C247_U1305 : INVD1 port map( A => mult_21_C247_n1535, Z => 
                           mult_21_C247_n1541);
   mult_21_C247_U1304 : NOR2D1 port map( A1 => mult_21_C247_n1537, A2 => 
                           mult_21_C247_n30, Z => mult_21_C247_n1093);
   mult_21_C247_U1303 : ADHALFDL port map( A => mult_21_C247_n1336, B => 
                           mult_21_C247_n1095, CO => mult_21_C247_n792, S => 
                           mult_21_C247_n793);
   mult_21_C247_U1302 : ADHALFDL port map( A => mult_21_C247_n1335, B => 
                           mult_21_C247_n1365, CO => mult_21_C247_n790, S => 
                           mult_21_C247_n791);
   mult_21_C247_U1301 : INVD1 port map( A => mult_21_C247_n1533, Z => 
                           mult_21_C247_n1542);
   mult_21_C247_U1300 : ADHALFDL port map( A => mult_21_C247_n1329, B => 
                           mult_21_C247_n1359, CO => mult_21_C247_n760, S => 
                           mult_21_C247_n761);
   mult_21_C247_U1299 : NOR2D1 port map( A1 => mult_21_C247_n303, A2 => 
                           mult_21_C247_n305, Z => mult_21_C247_n302);
   mult_21_C247_U1298 : NAN2D1 port map( A1 => mult_21_C247_n1368, A2 => 
                           mult_21_C247_n1096, Z => mult_21_C247_n305);
   mult_21_C247_U1297 : NAN2D1 port map( A1 => mult_21_C247_n791, A2 => 
                           mult_21_C247_n792, Z => mult_21_C247_n296);
   mult_21_C247_U1296 : NAN2D1 port map( A1 => mult_21_C247_n783, A2 => 
                           mult_21_C247_n786, Z => mult_21_C247_n288);
   mult_21_C247_U1295 : NOR2D1 port map( A1 => mult_21_C247_n791, A2 => 
                           mult_21_C247_n792, Z => mult_21_C247_n295);
   mult_21_C247_U1294 : NOR2D1 port map( A1 => mult_21_C247_n783, A2 => 
                           mult_21_C247_n786, Z => mult_21_C247_n287);
   mult_21_C247_U1293 : NAN2D1 port map( A1 => mult_21_C247_n777, A2 => 
                           mult_21_C247_n782, Z => mult_21_C247_n284);
   mult_21_C247_U1292 : NAN2D1 port map( A1 => mult_21_C247_n793, A2 => 
                           mult_21_C247_n1366, Z => mult_21_C247_n301);
   mult_21_C247_U1291 : NAN2D1 port map( A1 => mult_21_C247_n787, A2 => 
                           mult_21_C247_n789, Z => mult_21_C247_n293);
   mult_21_C247_U1290 : NOR2D1 port map( A1 => mult_21_C247_n777, A2 => 
                           mult_21_C247_n782, Z => mult_21_C247_n283);
   mult_21_C247_U1289 : OR2D1 port map( A1 => mult_21_C247_n793, A2 => 
                           mult_21_C247_n1366, Z => mult_21_C247_n1532);
   mult_21_C247_U1288 : OR2D1 port map( A1 => mult_21_C247_n787, A2 => 
                           mult_21_C247_n789, Z => mult_21_C247_n1531);
   mult_21_C247_U1287 : EXOR2D1 port map( A1 => mult_21_C247_n329, A2 => 
                           mult_21_C247_n344, Z => mult_21_C247_n155);
   mult_21_C247_U1286 : EXOR2D1 port map( A1 => mult_21_C247_n178, A2 => 
                           mult_21_C247_n155, Z => N3360);
   mult_21_C247_U1285 : NAN2D1 port map( A1 => mult_21_C247_n1532, A2 => 
                           mult_21_C247_n301, Z => mult_21_C247_n176);
   mult_21_C247_U1284 : INVD1 port map( A => mult_21_C247_n295, Z => 
                           mult_21_C247_n326);
   mult_21_C247_U1283 : NAN2D1 port map( A1 => mult_21_C247_n326, A2 => 
                           mult_21_C247_n296, Z => mult_21_C247_n175);
   mult_21_C247_U1282 : NAN2D1 port map( A1 => mult_21_C247_n1531, A2 => 
                           mult_21_C247_n293, Z => mult_21_C247_n174);
   mult_21_C247_U1281 : INVD1 port map( A => mult_21_C247_n287, Z => 
                           mult_21_C247_n324);
   mult_21_C247_U1280 : NAN2D1 port map( A1 => mult_21_C247_n324, A2 => 
                           mult_21_C247_n288, Z => mult_21_C247_n173);
   mult_21_C247_U1279 : INVD1 port map( A => mult_21_C247_n283, Z => 
                           mult_21_C247_n323);
   mult_21_C247_U1278 : NAN2D1 port map( A1 => mult_21_C247_n323, A2 => 
                           mult_21_C247_n284, Z => mult_21_C247_n172);
   mult_21_C247_U1277 : INVD1 port map( A => mult_21_C247_n280, Z => 
                           mult_21_C247_n322);
   mult_21_C247_U1276 : NAN2D1 port map( A1 => mult_21_C247_n322, A2 => 
                           mult_21_C247_n281, Z => mult_21_C247_n171);
   mult_21_C247_U1275 : NAN2D1 port map( A1 => mult_21_C247_n697, A2 => 
                           mult_21_C247_n710, Z => mult_21_C247_n240);
   mult_21_C247_U1274 : NAN2D1 port map( A1 => mult_21_C247_n711, A2 => 
                           mult_21_C247_n722, Z => mult_21_C247_n248);
   mult_21_C247_U1273 : NAN2D1 port map( A1 => mult_21_C247_n633, A2 => 
                           mult_21_C247_n650, Z => mult_21_C247_n221);
   mult_21_C247_U1272 : NOR2D1 port map( A1 => mult_21_C247_n615, A2 => 
                           mult_21_C247_n632, Z => mult_21_C247_n208);
   mult_21_C247_U1271 : NOR2D1 port map( A1 => mult_21_C247_n697, A2 => 
                           mult_21_C247_n710, Z => mult_21_C247_n239);
   mult_21_C247_U1270 : NAN2D1 port map( A1 => mult_21_C247_n735, A2 => 
                           mult_21_C247_n744, Z => mult_21_C247_n259);
   mult_21_C247_U1269 : NAN2D1 port map( A1 => mult_21_C247_n615, A2 => 
                           mult_21_C247_n632, Z => mult_21_C247_n209);
   mult_21_C247_U1268 : NAN2D1 port map( A1 => mult_21_C247_n771, A2 => 
                           mult_21_C247_n776, Z => mult_21_C247_n281);
   mult_21_C247_U1267 : OR2D1 port map( A1 => mult_21_C247_n711, A2 => 
                           mult_21_C247_n722, Z => mult_21_C247_n1530);
   mult_21_C247_U1266 : OR2D1 port map( A1 => mult_21_C247_n723, A2 => 
                           mult_21_C247_n734, Z => mult_21_C247_n1529);
   mult_21_C247_U1265 : NAN2D1 port map( A1 => mult_21_C247_n745, A2 => 
                           mult_21_C247_n754, Z => mult_21_C247_n262);
   mult_21_C247_U1264 : OR2D1 port map( A1 => mult_21_C247_n633, A2 => 
                           mult_21_C247_n650, Z => mult_21_C247_n1528);
   mult_21_C247_U1263 : NAN2D1 port map( A1 => mult_21_C247_n595, A2 => 
                           mult_21_C247_n614, Z => mult_21_C247_n206);
   mult_21_C247_U1262 : OR2D1 port map( A1 => mult_21_C247_n763, A2 => 
                           mult_21_C247_n770, Z => mult_21_C247_n1527);
   mult_21_C247_U1261 : NAN2D1 port map( A1 => mult_21_C247_n651, A2 => 
                           mult_21_C247_n666, Z => mult_21_C247_n226);
   mult_21_C247_U1260 : NAN2D1 port map( A1 => mult_21_C247_n723, A2 => 
                           mult_21_C247_n734, Z => mult_21_C247_n253);
   mult_21_C247_U1259 : NAN2D1 port map( A1 => mult_21_C247_n575, A2 => 
                           mult_21_C247_n594, Z => mult_21_C247_n199);
   mult_21_C247_U1258 : OR2D1 port map( A1 => mult_21_C247_n575, A2 => 
                           mult_21_C247_n594, Z => mult_21_C247_n1526);
   mult_21_C247_U1257 : NAN2D1 port map( A1 => mult_21_C247_n763, A2 => 
                           mult_21_C247_n770, Z => mult_21_C247_n275);
   mult_21_C247_U1256 : NOR2D1 port map( A1 => mult_21_C247_n735, A2 => 
                           mult_21_C247_n744, Z => mult_21_C247_n258);
   mult_21_C247_U1255 : NOR2D1 port map( A1 => mult_21_C247_n745, A2 => 
                           mult_21_C247_n754, Z => mult_21_C247_n261);
   mult_21_C247_U1254 : NOR2D1 port map( A1 => mult_21_C247_n771, A2 => 
                           mult_21_C247_n776, Z => mult_21_C247_n280);
   mult_21_C247_U1253 : OR2D1 port map( A1 => mult_21_C247_n595, A2 => 
                           mult_21_C247_n614, Z => mult_21_C247_n1525);
   mult_21_C247_U1252 : OA21M20D1 port map( A1 => mult_21_C247_n1532, A2 => 
                           mult_21_C247_n302, B => mult_21_C247_n301, Z => 
                           mult_21_C247_n297);
   mult_21_C247_U1251 : NOR2D1 port map( A1 => mult_21_C247_n651, A2 => 
                           mult_21_C247_n666, Z => mult_21_C247_n225);
   mult_21_C247_U1250 : OA21M20D1 port map( A1 => mult_21_C247_n1531, A2 => 
                           mult_21_C247_n294, B => mult_21_C247_n293, Z => 
                           mult_21_C247_n289);
   mult_21_C247_U1249 : NOR2D1 port map( A1 => mult_21_C247_n280, A2 => 
                           mult_21_C247_n283, Z => mult_21_C247_n278);
   mult_21_C247_U1248 : NAN2D1 port map( A1 => mult_21_C247_n755, A2 => 
                           mult_21_C247_n762, Z => mult_21_C247_n270);
   mult_21_C247_U1247 : OR2D1 port map( A1 => mult_21_C247_n755, A2 => 
                           mult_21_C247_n762, Z => mult_21_C247_n1524);
   mult_21_C247_U1246 : INVD1 port map( A => mult_21_C247_n286, Z => 
                           mult_21_C247_n285);
   mult_21_C247_U1245 : NAN2D1 port map( A1 => mult_21_C247_n1527, A2 => 
                           mult_21_C247_n275, Z => mult_21_C247_n170);
   mult_21_C247_U1244 : NAN2D1 port map( A1 => mult_21_C247_n1524, A2 => 
                           mult_21_C247_n270, Z => mult_21_C247_n169);
   mult_21_C247_U1243 : INVD1 port map( A => mult_21_C247_n277, Z => 
                           mult_21_C247_n276);
   mult_21_C247_U1242 : INVD1 port map( A => mult_21_C247_n261, Z => 
                           mult_21_C247_n319);
   mult_21_C247_U1241 : NAN2D1 port map( A1 => mult_21_C247_n319, A2 => 
                           mult_21_C247_n262, Z => mult_21_C247_n168);
   mult_21_C247_U1240 : INVD1 port map( A => mult_21_C247_n258, Z => 
                           mult_21_C247_n318);
   mult_21_C247_U1239 : NAN2D1 port map( A1 => mult_21_C247_n318, A2 => 
                           mult_21_C247_n259, Z => mult_21_C247_n167);
   mult_21_C247_U1238 : NAN2D1 port map( A1 => mult_21_C247_n1529, A2 => 
                           mult_21_C247_n253, Z => mult_21_C247_n166);
   mult_21_C247_U1237 : INVD1 port map( A => mult_21_C247_n239, Z => 
                           mult_21_C247_n315);
   mult_21_C247_U1236 : NAN2D1 port map( A1 => mult_21_C247_n315, A2 => 
                           mult_21_C247_n240, Z => mult_21_C247_n164);
   mult_21_C247_U1235 : NAN2D1 port map( A1 => mult_21_C247_n1530, A2 => 
                           mult_21_C247_n248, Z => mult_21_C247_n165);
   mult_21_C247_U1234 : INVD1 port map( A => mult_21_C247_n236, Z => 
                           mult_21_C247_n314);
   mult_21_C247_U1233 : NAN2D1 port map( A1 => mult_21_C247_n314, A2 => 
                           mult_21_C247_n237, Z => mult_21_C247_n163);
   mult_21_C247_U1232 : NAN2D1 port map( A1 => mult_21_C247_n1528, A2 => 
                           mult_21_C247_n221, Z => mult_21_C247_n160);
   mult_21_C247_U1231 : INVD1 port map( A => mult_21_C247_n225, Z => 
                           mult_21_C247_n312);
   mult_21_C247_U1230 : NAN2D1 port map( A1 => mult_21_C247_n312, A2 => 
                           mult_21_C247_n226, Z => mult_21_C247_n161);
   mult_21_C247_U1229 : NAN2D1 port map( A1 => mult_21_C247_n310, A2 => 
                           mult_21_C247_n209, Z => mult_21_C247_n159);
   mult_21_C247_U1228 : NAN2D1 port map( A1 => mult_21_C247_n1525, A2 => 
                           mult_21_C247_n206, Z => mult_21_C247_n158);
   mult_21_C247_U1227 : NAN2D1 port map( A1 => mult_21_C247_n1526, A2 => 
                           mult_21_C247_n199, Z => mult_21_C247_n157);
   mult_21_C247_U1226 : NAN2D1 port map( A1 => mult_21_C247_n1523, A2 => 
                           mult_21_C247_n194, Z => mult_21_C247_n156);
   mult_21_C247_U1225 : NAN2D1 port map( A1 => mult_21_C247_n683, A2 => 
                           mult_21_C247_n696, Z => mult_21_C247_n237);
   mult_21_C247_U1224 : INVD1 port map( A => mult_21_C247_n208, Z => 
                           mult_21_C247_n310);
   mult_21_C247_U1223 : NOR2D1 port map( A1 => mult_21_C247_n667, A2 => 
                           mult_21_C247_n682, Z => mult_21_C247_n230);
   mult_21_C247_U1222 : NAN2D1 port map( A1 => mult_21_C247_n553, A2 => 
                           mult_21_C247_n574, Z => mult_21_C247_n194);
   mult_21_C247_U1221 : NOR2D1 port map( A1 => mult_21_C247_n683, A2 => 
                           mult_21_C247_n696, Z => mult_21_C247_n236);
   mult_21_C247_U1220 : NAN2D1 port map( A1 => mult_21_C247_n1525, A2 => 
                           mult_21_C247_n310, Z => mult_21_C247_n201);
   mult_21_C247_U1219 : NOR2D1 port map( A1 => mult_21_C247_n225, A2 => 
                           mult_21_C247_n230, Z => mult_21_C247_n223);
   mult_21_C247_U1218 : INVD1 port map( A => mult_21_C247_n253, Z => 
                           mult_21_C247_n251);
   mult_21_C247_U1217 : NAN2D1 port map( A1 => mult_21_C247_n667, A2 => 
                           mult_21_C247_n682, Z => mult_21_C247_n231);
   mult_21_C247_U1216 : INVD1 port map( A => mult_21_C247_n199, Z => 
                           mult_21_C247_n197);
   mult_21_C247_U1215 : NAN2D1 port map( A1 => mult_21_C247_n1523, A2 => 
                           mult_21_C247_n1526, Z => mult_21_C247_n189);
   mult_21_C247_U1214 : OR2D1 port map( A1 => mult_21_C247_n553, A2 => 
                           mult_21_C247_n574, Z => mult_21_C247_n1523);
   mult_21_C247_U1213 : INVD1 port map( A => mult_21_C247_n275, Z => 
                           mult_21_C247_n273);
   mult_21_C247_U1212 : INVD1 port map( A => mult_21_C247_n206, Z => 
                           mult_21_C247_n204);
   mult_21_C247_U1211 : INVD1 port map( A => mult_21_C247_n209, Z => 
                           mult_21_C247_n211);
   mult_21_C247_U1210 : NOR2D1 port map( A1 => mult_21_C247_n189, A2 => 
                           mult_21_C247_n201, Z => mult_21_C247_n187);
   mult_21_C247_U1209 : NOR2D1 port map( A1 => mult_21_C247_n236, A2 => 
                           mult_21_C247_n239, Z => mult_21_C247_n234);
   mult_21_C247_U1208 : NOR2D1 port map( A1 => mult_21_C247_n258, A2 => 
                           mult_21_C247_n261, Z => mult_21_C247_n256);
   mult_21_C247_U1207 : INVD1 port map( A => mult_21_C247_n270, Z => 
                           mult_21_C247_n268);
   mult_21_C247_U1206 : NAN2D1 port map( A1 => mult_21_C247_n1524, A2 => 
                           mult_21_C247_n1527, Z => mult_21_C247_n265);
   mult_21_C247_U1205 : INVD1 port map( A => mult_21_C247_n248, Z => 
                           mult_21_C247_n246);
   mult_21_C247_U1204 : NAN2D1 port map( A1 => mult_21_C247_n1530, A2 => 
                           mult_21_C247_n1529, Z => mult_21_C247_n243);
   mult_21_C247_U1203 : INVD1 port map( A => mult_21_C247_n221, Z => 
                           mult_21_C247_n219);
   mult_21_C247_U1202 : NAN2D1 port map( A1 => mult_21_C247_n223, A2 => 
                           mult_21_C247_n1528, Z => mult_21_C247_n216);
   mult_21_C247_U1201 : INVD1 port map( A => mult_21_C247_n264, Z => 
                           mult_21_C247_n263);
   mult_21_C247_U1200 : INVD1 port map( A => mult_21_C247_n231, Z => 
                           mult_21_C247_n229);
   mult_21_C247_U1199 : INVD1 port map( A => mult_21_C247_n230, Z => 
                           mult_21_C247_n313);
   mult_21_C247_U1198 : INVD1 port map( A => mult_21_C247_n255, Z => 
                           mult_21_C247_n254);
   mult_21_C247_U1197 : INVD1 port map( A => mult_21_C247_n242, Z => 
                           mult_21_C247_n241);
   mult_21_C247_U1196 : NAN2D1 port map( A1 => mult_21_C247_n313, A2 => 
                           mult_21_C247_n231, Z => mult_21_C247_n162);
   mult_21_C247_U1195 : INVD1 port map( A => mult_21_C247_n233, Z => 
                           mult_21_C247_n232);
   mult_21_C247_U1194 : INVD1 port map( A => mult_21_C247_n215, Z => 
                           mult_21_C247_n214);
   mult_21_C247_U1193 : OA21M20D1 port map( A1 => mult_21_C247_n1523, A2 => 
                           mult_21_C247_n197, B => mult_21_C247_n194, Z => 
                           mult_21_C247_n190);
   mult_21_C247_U1192 : OR2D1 port map( A1 => mult_21_C247_n1368, A2 => 
                           mult_21_C247_n1096, Z => mult_21_C247_n1522);
   mult_21_C247_U1191 : AO21D1 port map( A1 => mult_21_C247_n215, A2 => 
                           mult_21_C247_n187, B => mult_21_C247_n188, Z => 
                           mult_21_C247_n1521);
   mult_21_C247_U1190 : AND2D1 port map( A1 => mult_21_C247_n1522, A2 => 
                           mult_21_C247_n305, Z => N3329);
   mult_21_C247_U1189 : OAI21D1 port map( A1 => N3016, A2 => N3017, B => 
                           mult_21_C247_n1077, Z => mult_21_C247_n1519);
   mult_21_C247_U1188 : OAI21D1 port map( A1 => N3012, A2 => N3013, B => 
                           mult_21_C247_n1079, Z => mult_21_C247_n1518);
   mult_21_C247_U1187 : OAI21D1 port map( A1 => N3010, A2 => N3011, B => 
                           mult_21_C247_n1080, Z => mult_21_C247_n1517);
   mult_21_C247_U1186 : ADHALFDL port map( A => mult_21_C247_n1278, B => 
                           mult_21_C247_n1093, CO => mult_21_C247_n780, S => 
                           mult_21_C247_n781);
   mult_21_C247_U1135 : EXNOR2D1 port map( A1 => N3032, A2 => N3033, Z => 
                           mult_21_C247_n93);
   mult_21_C247_U1131 : EXNOR2D1 port map( A1 => N3034, A2 => N3035, Z => 
                           mult_21_C247_n98);
   mult_21_C247_U1129 : OAI21D1 port map( A1 => N3034, A2 => N3035, B => 
                           mult_21_C247_n1068, Z => mult_21_C247_n94);
   mult_21_C247_U1127 : EXNOR2D1 port map( A1 => N3036, A2 => N3037, Z => 
                           mult_21_C247_n103);
   mult_21_C247_U1125 : OAI21D1 port map( A1 => N3036, A2 => N3037, B => 
                           mult_21_C247_n1067, Z => mult_21_C247_n99);
   mult_21_C247_U1123 : EXNOR2D1 port map( A1 => N3038, A2 => N3039, Z => 
                           mult_21_C247_n106);
   mult_21_C247_U1121 : OAI21D1 port map( A1 => N3038, A2 => N3039, B => 
                           mult_21_C247_n1066, Z => mult_21_C247_n104);
   mult_21_C247_U1120 : NAN2M1D1 port map( A1 => mult_21_C247_n8, A2 => 
                           mult_21_C247_n1556, Z => mult_21_C247_n1065);
   mult_21_C247_U1119 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1065, Z => 
                           mult_21_C247_n1368);
   mult_21_C247_U1118 : MUXB2DL port map( A0 => n283, A1 => mult_21_C247_n1556,
                           SL => mult_21_C247_n8, Z => mult_21_C247_n1064);
   mult_21_C247_U1117 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1064, Z => 
                           mult_21_C247_n1367);
   mult_21_C247_U1116 : MUXB2DL port map( A0 => mult_21_C247_n1553, A1 => n283,
                           SL => mult_21_C247_n8, Z => mult_21_C247_n1063);
   mult_21_C247_U1115 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1063, Z => 
                           mult_21_C247_n1366);
   mult_21_C247_U1114 : MUXB2DL port map( A0 => n286, A1 => mult_21_C247_n1554,
                           SL => mult_21_C247_n8, Z => mult_21_C247_n1062);
   mult_21_C247_U1113 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1062, Z => 
                           mult_21_C247_n1365);
   mult_21_C247_U1112 : MUXB2DL port map( A0 => mult_21_C247_n1549, A1 => 
                           mult_21_C247_n1551, SL => mult_21_C247_n8, Z => 
                           mult_21_C247_n1061);
   mult_21_C247_U1111 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1061, Z => 
                           mult_21_C247_n1364);
   mult_21_C247_U1110 : MUXB2DL port map( A0 => n282, A1 => n287, SL => 
                           mult_21_C247_n8, Z => mult_21_C247_n1060);
   mult_21_C247_U1109 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1060, Z => 
                           mult_21_C247_n1363);
   mult_21_C247_U1108 : MUXB2DL port map( A0 => n278, A1 => mult_21_C247_n1547,
                           SL => mult_21_C247_n8, Z => mult_21_C247_n1059);
   mult_21_C247_U1107 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1059, Z => 
                           mult_21_C247_n1362);
   mult_21_C247_U1106 : MUXB2DL port map( A0 => n279, A1 => n278, SL => 
                           mult_21_C247_n8, Z => mult_21_C247_n1058);
   mult_21_C247_U1105 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1058, Z => 
                           mult_21_C247_n1361);
   mult_21_C247_U1104 : MUXB2DL port map( A0 => mult_21_C247_n1545, A1 => n279,
                           SL => mult_21_C247_n8, Z => mult_21_C247_n1057);
   mult_21_C247_U1103 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1057, Z => 
                           mult_21_C247_n1360);
   mult_21_C247_U1102 : MUXB2DL port map( A0 => n281, A1 => mult_21_C247_n1545,
                           SL => mult_21_C247_n8, Z => mult_21_C247_n1056);
   mult_21_C247_U1101 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1056, Z => 
                           mult_21_C247_n1359);
   mult_21_C247_U1100 : MUXB2DL port map( A0 => mult_21_C247_n1543, A1 => n281,
                           SL => mult_21_C247_n8, Z => mult_21_C247_n1055);
   mult_21_C247_U1099 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1055, Z => 
                           mult_21_C247_n1358);
   mult_21_C247_U1098 : MUXB2DL port map( A0 => n274, A1 => n285, SL => 
                           mult_21_C247_n8, Z => mult_21_C247_n1054);
   mult_21_C247_U1097 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1054, Z => 
                           mult_21_C247_n1357);
   mult_21_C247_U1096 : MUXB2DL port map( A0 => n271, A1 => n274, SL => 
                           mult_21_C247_n8, Z => mult_21_C247_n1053);
   mult_21_C247_U1095 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1053, Z => 
                           mult_21_C247_n1356);
   mult_21_C247_U1094 : MUXB2DL port map( A0 => n272, A1 => n271, SL => 
                           mult_21_C247_n8, Z => mult_21_C247_n1052);
   mult_21_C247_U1093 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1052, Z => 
                           mult_21_C247_n1355);
   mult_21_C247_U1092 : MUXB2DL port map( A0 => n273, A1 => n272, SL => 
                           mult_21_C247_n8, Z => mult_21_C247_n1051);
   mult_21_C247_U1091 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1051, Z => 
                           mult_21_C247_n1354);
   mult_21_C247_U1090 : MUXB2DL port map( A0 => n291, A1 => n273, SL => 
                           mult_21_C247_n8, Z => mult_21_C247_n1050);
   mult_21_C247_U1089 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1050, Z => 
                           mult_21_C247_n1353);
   mult_21_C247_U1088 : MUXB2DL port map( A0 => n292, A1 => n291, SL => 
                           mult_21_C247_n8, Z => mult_21_C247_n1049);
   mult_21_C247_U1087 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1049, Z => 
                           mult_21_C247_n1352);
   mult_21_C247_U1086 : MUXB2DL port map( A0 => n289, A1 => n292, SL => 
                           mult_21_C247_n8, Z => mult_21_C247_n1048);
   mult_21_C247_U1085 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1048, Z => 
                           mult_21_C247_n1351);
   mult_21_C247_U1084 : MUXB2DL port map( A0 => n290, A1 => n289, SL => 
                           mult_21_C247_n8, Z => mult_21_C247_n1047);
   mult_21_C247_U1083 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1047, Z => 
                           mult_21_C247_n1350);
   mult_21_C247_U1082 : MUXB2DL port map( A0 => n293, A1 => n290, SL => 
                           mult_21_C247_n8, Z => mult_21_C247_n1046);
   mult_21_C247_U1081 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1046, Z => 
                           mult_21_C247_n1349);
   mult_21_C247_U1080 : MUXB2DL port map( A0 => n294, A1 => n293, SL => 
                           mult_21_C247_n8, Z => mult_21_C247_n1045);
   mult_21_C247_U1079 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1045, Z => 
                           mult_21_C247_n1348);
   mult_21_C247_U1078 : MUXB2DL port map( A0 => n295, A1 => n294, SL => 
                           mult_21_C247_n8, Z => mult_21_C247_n1044);
   mult_21_C247_U1077 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1044, Z => 
                           mult_21_C247_n1347);
   mult_21_C247_U1076 : MUXB2DL port map( A0 => n296, A1 => n295, SL => 
                           mult_21_C247_n8, Z => mult_21_C247_n1043);
   mult_21_C247_U1075 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1043, Z => 
                           mult_21_C247_n1346);
   mult_21_C247_U1074 : MUXB2DL port map( A0 => n297, A1 => n296, SL => 
                           mult_21_C247_n8, Z => mult_21_C247_n1042);
   mult_21_C247_U1073 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1042, Z => 
                           mult_21_C247_n1345);
   mult_21_C247_U1072 : MUXB2DL port map( A0 => n298, A1 => n297, SL => 
                           mult_21_C247_n8, Z => mult_21_C247_n1041);
   mult_21_C247_U1071 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1041, Z => 
                           mult_21_C247_n1344);
   mult_21_C247_U1070 : MUXB2DL port map( A0 => n299, A1 => n298, SL => 
                           mult_21_C247_n8, Z => mult_21_C247_n1040);
   mult_21_C247_U1069 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1040, Z => 
                           mult_21_C247_n1343);
   mult_21_C247_U1068 : MUXB2DL port map( A0 => n302, A1 => n299, SL => 
                           mult_21_C247_n8, Z => mult_21_C247_n1039);
   mult_21_C247_U1067 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1039, Z => 
                           mult_21_C247_n1342);
   mult_21_C247_U1066 : MUXB2DL port map( A0 => n303, A1 => n302, SL => 
                           mult_21_C247_n8, Z => mult_21_C247_n1038);
   mult_21_C247_U1065 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1038, Z => 
                           mult_21_C247_n1341);
   mult_21_C247_U1064 : MUXB2DL port map( A0 => n305, A1 => n303, SL => 
                           mult_21_C247_n8, Z => mult_21_C247_n1037);
   mult_21_C247_U1063 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1037, Z => 
                           mult_21_C247_n1340);
   mult_21_C247_U1062 : MUXB2DL port map( A0 => n310, A1 => n305, SL => 
                           mult_21_C247_n8, Z => mult_21_C247_n1036);
   mult_21_C247_U1061 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1036, Z => 
                           mult_21_C247_n1339);
   mult_21_C247_U1060 : MUXB2DL port map( A0 => n311, A1 => n310, SL => 
                           mult_21_C247_n8, Z => mult_21_C247_n1035);
   mult_21_C247_U1059 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1035, Z => 
                           mult_21_C247_n1338);
   mult_21_C247_U1058 : MUXB2DL port map( A0 => n312, A1 => n311, SL => 
                           mult_21_C247_n8, Z => mult_21_C247_n1034);
   mult_21_C247_U1057 : MUXB2DL port map( A0 => mult_21_C247_n3, A1 => 
                           mult_21_C247_n6, SL => mult_21_C247_n1034, Z => 
                           mult_21_C247_n1337);
   mult_21_C247_U1056 : NOR2M1D1 port map( A1 => mult_21_C247_n3, A2 => 
                           mult_21_C247_n6, Z => mult_21_C247_n1096);
   mult_21_C247_U1055 : NAN2M1D1 port map( A1 => mult_21_C247_n1542, A2 => n288
                           , Z => mult_21_C247_n1033);
   mult_21_C247_U1054 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1033, Z => 
                           mult_21_C247_n1336);
   mult_21_C247_U1053 : MUXB2DL port map( A0 => n283, A1 => mult_21_C247_n1556,
                           SL => mult_21_C247_n1542, Z => mult_21_C247_n1032);
   mult_21_C247_U1052 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1032, Z => 
                           mult_21_C247_n1335);
   mult_21_C247_U1051 : MUXB2DL port map( A0 => mult_21_C247_n1553, A1 => n283,
                           SL => mult_21_C247_n1542, Z => mult_21_C247_n1031);
   mult_21_C247_U1050 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1031, Z => 
                           mult_21_C247_n1334);
   mult_21_C247_U1049 : MUXB2DL port map( A0 => n286, A1 => mult_21_C247_n1554,
                           SL => mult_21_C247_n1542, Z => mult_21_C247_n1030);
   mult_21_C247_U1048 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1030, Z => 
                           mult_21_C247_n1333);
   mult_21_C247_U1047 : MUXB2DL port map( A0 => mult_21_C247_n1549, A1 => 
                           mult_21_C247_n1551, SL => mult_21_C247_n1542, Z => 
                           mult_21_C247_n1029);
   mult_21_C247_U1046 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1029, Z => 
                           mult_21_C247_n1332);
   mult_21_C247_U1045 : MUXB2DL port map( A0 => n282, A1 => n287, SL => 
                           mult_21_C247_n1542, Z => mult_21_C247_n1028);
   mult_21_C247_U1044 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1028, Z => 
                           mult_21_C247_n1331);
   mult_21_C247_U1043 : MUXB2DL port map( A0 => n278, A1 => mult_21_C247_n1547,
                           SL => mult_21_C247_n1542, Z => mult_21_C247_n1027);
   mult_21_C247_U1042 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1027, Z => 
                           mult_21_C247_n1330);
   mult_21_C247_U1041 : MUXB2DL port map( A0 => n279, A1 => n278, SL => 
                           mult_21_C247_n1542, Z => mult_21_C247_n1026);
   mult_21_C247_U1040 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1026, Z => 
                           mult_21_C247_n1329);
   mult_21_C247_U1039 : MUXB2DL port map( A0 => mult_21_C247_n1545, A1 => n279,
                           SL => mult_21_C247_n1542, Z => mult_21_C247_n1025);
   mult_21_C247_U1038 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1025, Z => 
                           mult_21_C247_n1328);
   mult_21_C247_U1037 : MUXB2DL port map( A0 => n281, A1 => n280, SL => 
                           mult_21_C247_n1542, Z => mult_21_C247_n1024);
   mult_21_C247_U1036 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1024, Z => 
                           mult_21_C247_n1327);
   mult_21_C247_U1035 : MUXB2DL port map( A0 => mult_21_C247_n1543, A1 => n281,
                           SL => mult_21_C247_n1542, Z => mult_21_C247_n1023);
   mult_21_C247_U1034 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1023, Z => 
                           mult_21_C247_n1326);
   mult_21_C247_U1033 : MUXB2DL port map( A0 => n274, A1 => n285, SL => 
                           mult_21_C247_n1542, Z => mult_21_C247_n1022);
   mult_21_C247_U1032 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1022, Z => 
                           mult_21_C247_n1325);
   mult_21_C247_U1031 : MUXB2DL port map( A0 => n271, A1 => n274, SL => 
                           mult_21_C247_n1542, Z => mult_21_C247_n1021);
   mult_21_C247_U1030 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1021, Z => 
                           mult_21_C247_n1324);
   mult_21_C247_U1029 : MUXB2DL port map( A0 => n272, A1 => n271, SL => 
                           mult_21_C247_n1542, Z => mult_21_C247_n1020);
   mult_21_C247_U1028 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1020, Z => 
                           mult_21_C247_n1323);
   mult_21_C247_U1027 : MUXB2DL port map( A0 => n273, A1 => n272, SL => 
                           mult_21_C247_n1542, Z => mult_21_C247_n1019);
   mult_21_C247_U1026 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1019, Z => 
                           mult_21_C247_n1322);
   mult_21_C247_U1025 : MUXB2DL port map( A0 => n291, A1 => n273, SL => 
                           mult_21_C247_n1542, Z => mult_21_C247_n1018);
   mult_21_C247_U1024 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1018, Z => 
                           mult_21_C247_n1321);
   mult_21_C247_U1023 : MUXB2DL port map( A0 => n292, A1 => n291, SL => 
                           mult_21_C247_n1542, Z => mult_21_C247_n1017);
   mult_21_C247_U1022 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1017, Z => 
                           mult_21_C247_n1320);
   mult_21_C247_U1021 : MUXB2DL port map( A0 => n289, A1 => n292, SL => 
                           mult_21_C247_n1542, Z => mult_21_C247_n1016);
   mult_21_C247_U1020 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1016, Z => 
                           mult_21_C247_n1319);
   mult_21_C247_U1019 : MUXB2DL port map( A0 => n290, A1 => n289, SL => 
                           mult_21_C247_n1542, Z => mult_21_C247_n1015);
   mult_21_C247_U1018 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1015, Z => 
                           mult_21_C247_n1318);
   mult_21_C247_U1017 : MUXB2DL port map( A0 => n293, A1 => n290, SL => 
                           mult_21_C247_n1542, Z => mult_21_C247_n1014);
   mult_21_C247_U1016 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1014, Z => 
                           mult_21_C247_n1317);
   mult_21_C247_U1015 : MUXB2DL port map( A0 => n294, A1 => n293, SL => 
                           mult_21_C247_n1542, Z => mult_21_C247_n1013);
   mult_21_C247_U1014 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1013, Z => 
                           mult_21_C247_n1316);
   mult_21_C247_U1013 : MUXB2DL port map( A0 => n295, A1 => n294, SL => 
                           mult_21_C247_n1542, Z => mult_21_C247_n1012);
   mult_21_C247_U1012 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1012, Z => 
                           mult_21_C247_n1315);
   mult_21_C247_U1011 : MUXB2DL port map( A0 => n296, A1 => n295, SL => 
                           mult_21_C247_n1542, Z => mult_21_C247_n1011);
   mult_21_C247_U1010 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1011, Z => 
                           mult_21_C247_n1314);
   mult_21_C247_U1009 : MUXB2DL port map( A0 => n297, A1 => n296, SL => 
                           mult_21_C247_n1542, Z => mult_21_C247_n1010);
   mult_21_C247_U1008 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1010, Z => 
                           mult_21_C247_n1313);
   mult_21_C247_U1007 : MUXB2DL port map( A0 => n298, A1 => n297, SL => 
                           mult_21_C247_n1542, Z => mult_21_C247_n1009);
   mult_21_C247_U1006 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1009, Z => 
                           mult_21_C247_n1312);
   mult_21_C247_U1005 : MUXB2DL port map( A0 => n299, A1 => n298, SL => 
                           mult_21_C247_n1542, Z => mult_21_C247_n1008);
   mult_21_C247_U1004 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1008, Z => 
                           mult_21_C247_n1311);
   mult_21_C247_U1003 : MUXB2DL port map( A0 => n302, A1 => n299, SL => 
                           mult_21_C247_n1542, Z => mult_21_C247_n1007);
   mult_21_C247_U1002 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1007, Z => 
                           mult_21_C247_n1310);
   mult_21_C247_U1001 : MUXB2DL port map( A0 => n303, A1 => n302, SL => 
                           mult_21_C247_n1542, Z => mult_21_C247_n1006);
   mult_21_C247_U1000 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1006, Z => 
                           mult_21_C247_n1309);
   mult_21_C247_U999 : MUXB2DL port map( A0 => n305, A1 => n303, SL => 
                           mult_21_C247_n1542, Z => mult_21_C247_n1005);
   mult_21_C247_U998 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1005, Z => 
                           mult_21_C247_n1308);
   mult_21_C247_U997 : MUXB2DL port map( A0 => n310, A1 => n305, SL => 
                           mult_21_C247_n1542, Z => mult_21_C247_n1004);
   mult_21_C247_U996 : MUXB2DL port map( A0 => mult_21_C247_n1517, A1 => 
                           mult_21_C247_n14, SL => mult_21_C247_n1004, Z => 
                           mult_21_C247_n1307);
   mult_21_C247_U995 : NOR2M1D1 port map( A1 => mult_21_C247_n1517, A2 => 
                           mult_21_C247_n14, Z => mult_21_C247_n1095);
   mult_21_C247_U994 : NAN2M1D1 port map( A1 => mult_21_C247_n1541, A2 => n288,
                           Z => mult_21_C247_n1003);
   mult_21_C247_U993 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n1003, Z => 
                           mult_21_C247_n1306);
   mult_21_C247_U992 : MUXB2DL port map( A0 => n283, A1 => mult_21_C247_n1556, 
                           SL => mult_21_C247_n1541, Z => mult_21_C247_n1002);
   mult_21_C247_U991 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n1002, Z => 
                           mult_21_C247_n1305);
   mult_21_C247_U990 : MUXB2DL port map( A0 => mult_21_C247_n1553, A1 => n283, 
                           SL => mult_21_C247_n1541, Z => mult_21_C247_n1001);
   mult_21_C247_U989 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n1001, Z => 
                           mult_21_C247_n1304);
   mult_21_C247_U988 : MUXB2DL port map( A0 => n286, A1 => mult_21_C247_n1554, 
                           SL => mult_21_C247_n1541, Z => mult_21_C247_n1000);
   mult_21_C247_U987 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n1000, Z => 
                           mult_21_C247_n1303);
   mult_21_C247_U986 : MUXB2DL port map( A0 => mult_21_C247_n1549, A1 => 
                           mult_21_C247_n1551, SL => mult_21_C247_n1541, Z => 
                           mult_21_C247_n999);
   mult_21_C247_U985 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n999, Z => 
                           mult_21_C247_n1302);
   mult_21_C247_U984 : MUXB2DL port map( A0 => n282, A1 => n287, SL => 
                           mult_21_C247_n1541, Z => mult_21_C247_n998);
   mult_21_C247_U983 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n998, Z => 
                           mult_21_C247_n1301);
   mult_21_C247_U982 : MUXB2DL port map( A0 => n278, A1 => mult_21_C247_n1547, 
                           SL => mult_21_C247_n1541, Z => mult_21_C247_n997);
   mult_21_C247_U981 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n997, Z => 
                           mult_21_C247_n1300);
   mult_21_C247_U980 : MUXB2DL port map( A0 => n279, A1 => n278, SL => 
                           mult_21_C247_n1541, Z => mult_21_C247_n996);
   mult_21_C247_U979 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n996, Z => 
                           mult_21_C247_n1299);
   mult_21_C247_U978 : MUXB2DL port map( A0 => mult_21_C247_n1545, A1 => n279, 
                           SL => mult_21_C247_n1541, Z => mult_21_C247_n995);
   mult_21_C247_U977 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n995, Z => 
                           mult_21_C247_n1298);
   mult_21_C247_U976 : MUXB2DL port map( A0 => n281, A1 => n280, SL => 
                           mult_21_C247_n1541, Z => mult_21_C247_n994);
   mult_21_C247_U975 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n994, Z => 
                           mult_21_C247_n1297);
   mult_21_C247_U974 : MUXB2DL port map( A0 => mult_21_C247_n1543, A1 => n281, 
                           SL => mult_21_C247_n1541, Z => mult_21_C247_n993);
   mult_21_C247_U973 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n993, Z => 
                           mult_21_C247_n1296);
   mult_21_C247_U972 : MUXB2DL port map( A0 => n274, A1 => mult_21_C247_n1543, 
                           SL => mult_21_C247_n1541, Z => mult_21_C247_n992);
   mult_21_C247_U971 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n992, Z => 
                           mult_21_C247_n1295);
   mult_21_C247_U970 : MUXB2DL port map( A0 => n271, A1 => n274, SL => 
                           mult_21_C247_n1541, Z => mult_21_C247_n991);
   mult_21_C247_U969 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n991, Z => 
                           mult_21_C247_n1294);
   mult_21_C247_U968 : MUXB2DL port map( A0 => n272, A1 => n271, SL => 
                           mult_21_C247_n1541, Z => mult_21_C247_n990);
   mult_21_C247_U967 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n990, Z => 
                           mult_21_C247_n1293);
   mult_21_C247_U966 : MUXB2DL port map( A0 => n273, A1 => n272, SL => 
                           mult_21_C247_n1541, Z => mult_21_C247_n989);
   mult_21_C247_U965 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n989, Z => 
                           mult_21_C247_n1292);
   mult_21_C247_U964 : MUXB2DL port map( A0 => n291, A1 => n273, SL => 
                           mult_21_C247_n1541, Z => mult_21_C247_n988);
   mult_21_C247_U963 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n988, Z => 
                           mult_21_C247_n1291);
   mult_21_C247_U962 : MUXB2DL port map( A0 => n292, A1 => n291, SL => 
                           mult_21_C247_n1541, Z => mult_21_C247_n987);
   mult_21_C247_U961 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n987, Z => 
                           mult_21_C247_n1290);
   mult_21_C247_U960 : MUXB2DL port map( A0 => n289, A1 => n292, SL => 
                           mult_21_C247_n1541, Z => mult_21_C247_n986);
   mult_21_C247_U959 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n986, Z => 
                           mult_21_C247_n1289);
   mult_21_C247_U958 : MUXB2DL port map( A0 => n290, A1 => n289, SL => 
                           mult_21_C247_n1541, Z => mult_21_C247_n985);
   mult_21_C247_U957 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n985, Z => 
                           mult_21_C247_n1288);
   mult_21_C247_U956 : MUXB2DL port map( A0 => n293, A1 => n290, SL => 
                           mult_21_C247_n1541, Z => mult_21_C247_n984);
   mult_21_C247_U955 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n984, Z => 
                           mult_21_C247_n1287);
   mult_21_C247_U954 : MUXB2DL port map( A0 => n294, A1 => n293, SL => 
                           mult_21_C247_n1541, Z => mult_21_C247_n983);
   mult_21_C247_U953 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n983, Z => 
                           mult_21_C247_n1286);
   mult_21_C247_U952 : MUXB2DL port map( A0 => n295, A1 => n294, SL => 
                           mult_21_C247_n1541, Z => mult_21_C247_n982);
   mult_21_C247_U951 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n982, Z => 
                           mult_21_C247_n1285);
   mult_21_C247_U950 : MUXB2DL port map( A0 => n296, A1 => n295, SL => 
                           mult_21_C247_n1541, Z => mult_21_C247_n981);
   mult_21_C247_U949 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n981, Z => 
                           mult_21_C247_n1284);
   mult_21_C247_U948 : MUXB2DL port map( A0 => n297, A1 => n296, SL => 
                           mult_21_C247_n1541, Z => mult_21_C247_n980);
   mult_21_C247_U947 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n980, Z => 
                           mult_21_C247_n1283);
   mult_21_C247_U946 : MUXB2DL port map( A0 => n298, A1 => n297, SL => 
                           mult_21_C247_n1541, Z => mult_21_C247_n979);
   mult_21_C247_U945 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n979, Z => 
                           mult_21_C247_n1282);
   mult_21_C247_U944 : MUXB2DL port map( A0 => n299, A1 => n298, SL => 
                           mult_21_C247_n1541, Z => mult_21_C247_n978);
   mult_21_C247_U943 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n978, Z => 
                           mult_21_C247_n1281);
   mult_21_C247_U942 : MUXB2DL port map( A0 => n302, A1 => n299, SL => 
                           mult_21_C247_n1541, Z => mult_21_C247_n977);
   mult_21_C247_U941 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n977, Z => 
                           mult_21_C247_n1280);
   mult_21_C247_U940 : MUXB2DL port map( A0 => n303, A1 => n302, SL => 
                           mult_21_C247_n1541, Z => mult_21_C247_n976);
   mult_21_C247_U939 : MUXB2DL port map( A0 => mult_21_C247_n1518, A1 => 
                           mult_21_C247_n22, SL => mult_21_C247_n976, Z => 
                           mult_21_C247_n1279);
   mult_21_C247_U938 : NOR2M1D1 port map( A1 => mult_21_C247_n1518, A2 => 
                           mult_21_C247_n22, Z => mult_21_C247_n1094);
   mult_21_C247_U937 : NAN2M1D1 port map( A1 => mult_21_C247_n1539, A2 => n288,
                           Z => mult_21_C247_n975);
   mult_21_C247_U936 : MUXB2DL port map( A0 => mult_21_C247_n1540, A1 => 
                           mult_21_C247_n30, SL => mult_21_C247_n975, Z => 
                           mult_21_C247_n1278);
   mult_21_C247_U935 : MUXB2DL port map( A0 => n283, A1 => n288, SL => 
                           mult_21_C247_n1539, Z => mult_21_C247_n974);
   mult_21_C247_U934 : MUXB2DL port map( A0 => mult_21_C247_n1540, A1 => 
                           mult_21_C247_n30, SL => mult_21_C247_n974, Z => 
                           mult_21_C247_n1277);
   mult_21_C247_U933 : MUXB2DL port map( A0 => mult_21_C247_n1553, A1 => n283, 
                           SL => mult_21_C247_n1539, Z => mult_21_C247_n973);
   mult_21_C247_U932 : MUXB2DL port map( A0 => mult_21_C247_n1540, A1 => 
                           mult_21_C247_n30, SL => mult_21_C247_n973, Z => 
                           mult_21_C247_n1276);
   mult_21_C247_U931 : MUXB2DL port map( A0 => n286, A1 => mult_21_C247_n1553, 
                           SL => mult_21_C247_n1539, Z => mult_21_C247_n972);
   mult_21_C247_U930 : MUXB2DL port map( A0 => mult_21_C247_n1540, A1 => 
                           mult_21_C247_n30, SL => mult_21_C247_n972, Z => 
                           mult_21_C247_n1275);
   mult_21_C247_U929 : MUXB2DL port map( A0 => mult_21_C247_n1549, A1 => n286, 
                           SL => mult_21_C247_n1539, Z => mult_21_C247_n971);
   mult_21_C247_U928 : MUXB2DL port map( A0 => mult_21_C247_n1540, A1 => 
                           mult_21_C247_n30, SL => mult_21_C247_n971, Z => 
                           mult_21_C247_n1274);
   mult_21_C247_U927 : MUXB2DL port map( A0 => n282, A1 => mult_21_C247_n1549, 
                           SL => mult_21_C247_n1539, Z => mult_21_C247_n970);
   mult_21_C247_U926 : MUXB2DL port map( A0 => mult_21_C247_n1540, A1 => 
                           mult_21_C247_n30, SL => mult_21_C247_n970, Z => 
                           mult_21_C247_n1273);
   mult_21_C247_U925 : MUXB2DL port map( A0 => n278, A1 => mult_21_C247_n1547, 
                           SL => mult_21_C247_n1539, Z => mult_21_C247_n969);
   mult_21_C247_U924 : MUXB2DL port map( A0 => mult_21_C247_n1540, A1 => 
                           mult_21_C247_n30, SL => mult_21_C247_n969, Z => 
                           mult_21_C247_n1272);
   mult_21_C247_U923 : MUXB2DL port map( A0 => n279, A1 => n278, SL => 
                           mult_21_C247_n1539, Z => mult_21_C247_n968);
   mult_21_C247_U922 : MUXB2DL port map( A0 => mult_21_C247_n1540, A1 => 
                           mult_21_C247_n30, SL => mult_21_C247_n968, Z => 
                           mult_21_C247_n1271);
   mult_21_C247_U921 : MUXB2DL port map( A0 => mult_21_C247_n1545, A1 => n279, 
                           SL => mult_21_C247_n1539, Z => mult_21_C247_n967);
   mult_21_C247_U920 : MUXB2DL port map( A0 => mult_21_C247_n1540, A1 => 
                           mult_21_C247_n30, SL => mult_21_C247_n967, Z => 
                           mult_21_C247_n1270);
   mult_21_C247_U919 : MUXB2DL port map( A0 => n281, A1 => n280, SL => 
                           mult_21_C247_n1539, Z => mult_21_C247_n966);
   mult_21_C247_U918 : MUXB2DL port map( A0 => mult_21_C247_n1540, A1 => 
                           mult_21_C247_n30, SL => mult_21_C247_n966, Z => 
                           mult_21_C247_n1269);
   mult_21_C247_U917 : MUXB2DL port map( A0 => mult_21_C247_n1543, A1 => n281, 
                           SL => mult_21_C247_n1539, Z => mult_21_C247_n965);
   mult_21_C247_U916 : MUXB2DL port map( A0 => mult_21_C247_n1540, A1 => 
                           mult_21_C247_n30, SL => mult_21_C247_n965, Z => 
                           mult_21_C247_n1268);
   mult_21_C247_U915 : MUXB2DL port map( A0 => n274, A1 => n285, SL => 
                           mult_21_C247_n1539, Z => mult_21_C247_n964);
   mult_21_C247_U914 : MUXB2DL port map( A0 => mult_21_C247_n1540, A1 => 
                           mult_21_C247_n30, SL => mult_21_C247_n964, Z => 
                           mult_21_C247_n1267);
   mult_21_C247_U913 : MUXB2DL port map( A0 => n271, A1 => n274, SL => 
                           mult_21_C247_n1539, Z => mult_21_C247_n963);
   mult_21_C247_U912 : MUXB2DL port map( A0 => mult_21_C247_n1540, A1 => 
                           mult_21_C247_n30, SL => mult_21_C247_n963, Z => 
                           mult_21_C247_n1266);
   mult_21_C247_U911 : MUXB2DL port map( A0 => n272, A1 => n271, SL => 
                           mult_21_C247_n1539, Z => mult_21_C247_n962);
   mult_21_C247_U910 : MUXB2DL port map( A0 => mult_21_C247_n1540, A1 => 
                           mult_21_C247_n30, SL => mult_21_C247_n962, Z => 
                           mult_21_C247_n1265);
   mult_21_C247_U909 : MUXB2DL port map( A0 => n273, A1 => n272, SL => 
                           mult_21_C247_n1539, Z => mult_21_C247_n961);
   mult_21_C247_U908 : MUXB2DL port map( A0 => mult_21_C247_n1540, A1 => 
                           mult_21_C247_n30, SL => mult_21_C247_n961, Z => 
                           mult_21_C247_n1264);
   mult_21_C247_U907 : MUXB2DL port map( A0 => n291, A1 => n273, SL => 
                           mult_21_C247_n1539, Z => mult_21_C247_n960);
   mult_21_C247_U906 : MUXB2DL port map( A0 => mult_21_C247_n1540, A1 => 
                           mult_21_C247_n30, SL => mult_21_C247_n960, Z => 
                           mult_21_C247_n1263);
   mult_21_C247_U905 : MUXB2DL port map( A0 => n292, A1 => n291, SL => 
                           mult_21_C247_n1539, Z => mult_21_C247_n959);
   mult_21_C247_U904 : MUXB2DL port map( A0 => mult_21_C247_n1540, A1 => 
                           mult_21_C247_n30, SL => mult_21_C247_n959, Z => 
                           mult_21_C247_n1262);
   mult_21_C247_U903 : MUXB2DL port map( A0 => n289, A1 => n292, SL => 
                           mult_21_C247_n1539, Z => mult_21_C247_n958);
   mult_21_C247_U902 : MUXB2DL port map( A0 => mult_21_C247_n1540, A1 => 
                           mult_21_C247_n30, SL => mult_21_C247_n958, Z => 
                           mult_21_C247_n1261);
   mult_21_C247_U901 : MUXB2DL port map( A0 => n290, A1 => n289, SL => 
                           mult_21_C247_n1539, Z => mult_21_C247_n957);
   mult_21_C247_U900 : MUXB2DL port map( A0 => mult_21_C247_n1540, A1 => 
                           mult_21_C247_n30, SL => mult_21_C247_n957, Z => 
                           mult_21_C247_n1260);
   mult_21_C247_U899 : MUXB2DL port map( A0 => n293, A1 => n290, SL => 
                           mult_21_C247_n1539, Z => mult_21_C247_n956);
   mult_21_C247_U898 : MUXB2DL port map( A0 => mult_21_C247_n1540, A1 => 
                           mult_21_C247_n30, SL => mult_21_C247_n956, Z => 
                           mult_21_C247_n1259);
   mult_21_C247_U897 : MUXB2DL port map( A0 => n294, A1 => n293, SL => 
                           mult_21_C247_n1539, Z => mult_21_C247_n955);
   mult_21_C247_U896 : MUXB2DL port map( A0 => mult_21_C247_n1540, A1 => 
                           mult_21_C247_n30, SL => mult_21_C247_n955, Z => 
                           mult_21_C247_n1258);
   mult_21_C247_U895 : MUXB2DL port map( A0 => n295, A1 => n294, SL => 
                           mult_21_C247_n1539, Z => mult_21_C247_n954);
   mult_21_C247_U894 : MUXB2DL port map( A0 => mult_21_C247_n1540, A1 => 
                           mult_21_C247_n30, SL => mult_21_C247_n954, Z => 
                           mult_21_C247_n1257);
   mult_21_C247_U893 : MUXB2DL port map( A0 => n296, A1 => n295, SL => 
                           mult_21_C247_n1539, Z => mult_21_C247_n953);
   mult_21_C247_U892 : MUXB2DL port map( A0 => mult_21_C247_n1540, A1 => 
                           mult_21_C247_n30, SL => mult_21_C247_n953, Z => 
                           mult_21_C247_n1256);
   mult_21_C247_U891 : MUXB2DL port map( A0 => n297, A1 => n296, SL => 
                           mult_21_C247_n1539, Z => mult_21_C247_n952);
   mult_21_C247_U890 : MUXB2DL port map( A0 => mult_21_C247_n1540, A1 => 
                           mult_21_C247_n30, SL => mult_21_C247_n952, Z => 
                           mult_21_C247_n1255);
   mult_21_C247_U889 : MUXB2DL port map( A0 => n298, A1 => n297, SL => 
                           mult_21_C247_n1539, Z => mult_21_C247_n951);
   mult_21_C247_U888 : MUXB2DL port map( A0 => mult_21_C247_n1540, A1 => 
                           mult_21_C247_n30, SL => mult_21_C247_n951, Z => 
                           mult_21_C247_n1254);
   mult_21_C247_U887 : MUXB2DL port map( A0 => n299, A1 => n298, SL => 
                           mult_21_C247_n1539, Z => mult_21_C247_n950);
   mult_21_C247_U886 : MUXB2DL port map( A0 => mult_21_C247_n1540, A1 => 
                           mult_21_C247_n30, SL => mult_21_C247_n950, Z => 
                           mult_21_C247_n1253);
   mult_21_C247_U884 : NAN2M1D1 port map( A1 => mult_21_C247_n1538, A2 => n288,
                           Z => mult_21_C247_n949);
   mult_21_C247_U883 : MUXB2DL port map( A0 => mult_21_C247_n1519, A1 => 
                           mult_21_C247_n38, SL => mult_21_C247_n949, Z => 
                           mult_21_C247_n1252);
   mult_21_C247_U882 : MUXB2DL port map( A0 => n283, A1 => n288, SL => 
                           mult_21_C247_n1538, Z => mult_21_C247_n948);
   mult_21_C247_U881 : MUXB2DL port map( A0 => mult_21_C247_n1519, A1 => 
                           mult_21_C247_n38, SL => mult_21_C247_n948, Z => 
                           mult_21_C247_n1251);
   mult_21_C247_U880 : MUXB2DL port map( A0 => mult_21_C247_n1553, A1 => n283, 
                           SL => mult_21_C247_n1538, Z => mult_21_C247_n947);
   mult_21_C247_U879 : MUXB2DL port map( A0 => mult_21_C247_n1519, A1 => 
                           mult_21_C247_n38, SL => mult_21_C247_n947, Z => 
                           mult_21_C247_n1250);
   mult_21_C247_U878 : MUXB2DL port map( A0 => n286, A1 => mult_21_C247_n1553, 
                           SL => mult_21_C247_n1538, Z => mult_21_C247_n946);
   mult_21_C247_U877 : MUXB2DL port map( A0 => mult_21_C247_n1519, A1 => 
                           mult_21_C247_n38, SL => mult_21_C247_n946, Z => 
                           mult_21_C247_n1249);
   mult_21_C247_U876 : MUXB2DL port map( A0 => mult_21_C247_n1549, A1 => n286, 
                           SL => mult_21_C247_n1538, Z => mult_21_C247_n945);
   mult_21_C247_U875 : MUXB2DL port map( A0 => mult_21_C247_n1519, A1 => 
                           mult_21_C247_n38, SL => mult_21_C247_n945, Z => 
                           mult_21_C247_n1248);
   mult_21_C247_U874 : MUXB2DL port map( A0 => n282, A1 => n287, SL => 
                           mult_21_C247_n1538, Z => mult_21_C247_n944);
   mult_21_C247_U873 : MUXB2DL port map( A0 => mult_21_C247_n1519, A1 => 
                           mult_21_C247_n38, SL => mult_21_C247_n944, Z => 
                           mult_21_C247_n1247);
   mult_21_C247_U872 : MUXB2DL port map( A0 => n278, A1 => mult_21_C247_n1547, 
                           SL => mult_21_C247_n1538, Z => mult_21_C247_n943);
   mult_21_C247_U871 : MUXB2DL port map( A0 => mult_21_C247_n1519, A1 => 
                           mult_21_C247_n38, SL => mult_21_C247_n943, Z => 
                           mult_21_C247_n1246);
   mult_21_C247_U870 : MUXB2DL port map( A0 => n279, A1 => n278, SL => 
                           mult_21_C247_n1538, Z => mult_21_C247_n942);
   mult_21_C247_U869 : MUXB2DL port map( A0 => mult_21_C247_n1519, A1 => 
                           mult_21_C247_n38, SL => mult_21_C247_n942, Z => 
                           mult_21_C247_n1245);
   mult_21_C247_U868 : MUXB2DL port map( A0 => mult_21_C247_n1545, A1 => n279, 
                           SL => mult_21_C247_n1538, Z => mult_21_C247_n941);
   mult_21_C247_U867 : MUXB2DL port map( A0 => mult_21_C247_n1519, A1 => 
                           mult_21_C247_n38, SL => mult_21_C247_n941, Z => 
                           mult_21_C247_n1244);
   mult_21_C247_U866 : MUXB2DL port map( A0 => n281, A1 => n280, SL => 
                           mult_21_C247_n1538, Z => mult_21_C247_n940);
   mult_21_C247_U865 : MUXB2DL port map( A0 => mult_21_C247_n1519, A1 => 
                           mult_21_C247_n38, SL => mult_21_C247_n940, Z => 
                           mult_21_C247_n1243);
   mult_21_C247_U864 : MUXB2DL port map( A0 => mult_21_C247_n1543, A1 => n281, 
                           SL => mult_21_C247_n1538, Z => mult_21_C247_n939);
   mult_21_C247_U863 : MUXB2DL port map( A0 => mult_21_C247_n1519, A1 => 
                           mult_21_C247_n38, SL => mult_21_C247_n939, Z => 
                           mult_21_C247_n1242);
   mult_21_C247_U862 : MUXB2DL port map( A0 => n274, A1 => mult_21_C247_n1543, 
                           SL => mult_21_C247_n1538, Z => mult_21_C247_n938);
   mult_21_C247_U861 : MUXB2DL port map( A0 => mult_21_C247_n1519, A1 => 
                           mult_21_C247_n38, SL => mult_21_C247_n938, Z => 
                           mult_21_C247_n1241);
   mult_21_C247_U860 : MUXB2DL port map( A0 => n271, A1 => n274, SL => 
                           mult_21_C247_n1538, Z => mult_21_C247_n937);
   mult_21_C247_U859 : MUXB2DL port map( A0 => mult_21_C247_n1519, A1 => 
                           mult_21_C247_n38, SL => mult_21_C247_n937, Z => 
                           mult_21_C247_n1240);
   mult_21_C247_U858 : MUXB2DL port map( A0 => n272, A1 => n271, SL => 
                           mult_21_C247_n1538, Z => mult_21_C247_n936);
   mult_21_C247_U857 : MUXB2DL port map( A0 => mult_21_C247_n1519, A1 => 
                           mult_21_C247_n38, SL => mult_21_C247_n936, Z => 
                           mult_21_C247_n1239);
   mult_21_C247_U856 : MUXB2DL port map( A0 => n273, A1 => n272, SL => 
                           mult_21_C247_n1538, Z => mult_21_C247_n935);
   mult_21_C247_U855 : MUXB2DL port map( A0 => mult_21_C247_n1519, A1 => 
                           mult_21_C247_n38, SL => mult_21_C247_n935, Z => 
                           mult_21_C247_n1238);
   mult_21_C247_U854 : MUXB2DL port map( A0 => n291, A1 => n273, SL => 
                           mult_21_C247_n1538, Z => mult_21_C247_n934);
   mult_21_C247_U853 : MUXB2DL port map( A0 => mult_21_C247_n1519, A1 => 
                           mult_21_C247_n38, SL => mult_21_C247_n934, Z => 
                           mult_21_C247_n1237);
   mult_21_C247_U852 : MUXB2DL port map( A0 => n292, A1 => n291, SL => 
                           mult_21_C247_n1538, Z => mult_21_C247_n933);
   mult_21_C247_U851 : MUXB2DL port map( A0 => mult_21_C247_n1519, A1 => 
                           mult_21_C247_n38, SL => mult_21_C247_n933, Z => 
                           mult_21_C247_n1236);
   mult_21_C247_U850 : MUXB2DL port map( A0 => n289, A1 => n292, SL => 
                           mult_21_C247_n1538, Z => mult_21_C247_n932);
   mult_21_C247_U849 : MUXB2DL port map( A0 => mult_21_C247_n1519, A1 => 
                           mult_21_C247_n38, SL => mult_21_C247_n932, Z => 
                           mult_21_C247_n1235);
   mult_21_C247_U848 : MUXB2DL port map( A0 => n290, A1 => n289, SL => 
                           mult_21_C247_n1538, Z => mult_21_C247_n931);
   mult_21_C247_U847 : MUXB2DL port map( A0 => mult_21_C247_n1519, A1 => 
                           mult_21_C247_n38, SL => mult_21_C247_n931, Z => 
                           mult_21_C247_n1234);
   mult_21_C247_U846 : MUXB2DL port map( A0 => n293, A1 => n290, SL => 
                           mult_21_C247_n1538, Z => mult_21_C247_n930);
   mult_21_C247_U845 : MUXB2DL port map( A0 => mult_21_C247_n1519, A1 => 
                           mult_21_C247_n38, SL => mult_21_C247_n930, Z => 
                           mult_21_C247_n1233);
   mult_21_C247_U844 : MUXB2DL port map( A0 => n294, A1 => n293, SL => 
                           mult_21_C247_n1538, Z => mult_21_C247_n929);
   mult_21_C247_U843 : MUXB2DL port map( A0 => mult_21_C247_n1519, A1 => 
                           mult_21_C247_n38, SL => mult_21_C247_n929, Z => 
                           mult_21_C247_n1232);
   mult_21_C247_U842 : MUXB2DL port map( A0 => n295, A1 => n294, SL => 
                           mult_21_C247_n1538, Z => mult_21_C247_n928);
   mult_21_C247_U841 : MUXB2DL port map( A0 => mult_21_C247_n1519, A1 => 
                           mult_21_C247_n38, SL => mult_21_C247_n928, Z => 
                           mult_21_C247_n1231);
   mult_21_C247_U840 : MUXB2DL port map( A0 => n296, A1 => n295, SL => 
                           mult_21_C247_n1538, Z => mult_21_C247_n927);
   mult_21_C247_U839 : MUXB2DL port map( A0 => mult_21_C247_n1519, A1 => 
                           mult_21_C247_n38, SL => mult_21_C247_n927, Z => 
                           mult_21_C247_n1230);
   mult_21_C247_U838 : MUXB2DL port map( A0 => n297, A1 => n296, SL => 
                           mult_21_C247_n1538, Z => mult_21_C247_n926);
   mult_21_C247_U837 : MUXB2DL port map( A0 => mult_21_C247_n1519, A1 => 
                           mult_21_C247_n38, SL => mult_21_C247_n926, Z => 
                           mult_21_C247_n1229);
   mult_21_C247_U836 : NOR2M1D1 port map( A1 => mult_21_C247_n1519, A2 => 
                           mult_21_C247_n38, Z => mult_21_C247_n1092);
   mult_21_C247_U835 : NAN2M1D1 port map( A1 => mult_21_C247_n48, A2 => n288, Z
                           => mult_21_C247_n925);
   mult_21_C247_U834 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n45, SL => mult_21_C247_n925, Z => 
                           mult_21_C247_n1228);
   mult_21_C247_U833 : MUXB2DL port map( A0 => n283, A1 => n288, SL => 
                           mult_21_C247_n48, Z => mult_21_C247_n924);
   mult_21_C247_U832 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n45, SL => mult_21_C247_n924, Z => 
                           mult_21_C247_n1227);
   mult_21_C247_U831 : MUXB2DL port map( A0 => mult_21_C247_n1553, A1 => n283, 
                           SL => mult_21_C247_n48, Z => mult_21_C247_n923);
   mult_21_C247_U830 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n45, SL => mult_21_C247_n923, Z => 
                           mult_21_C247_n1226);
   mult_21_C247_U829 : MUXB2DL port map( A0 => n286, A1 => mult_21_C247_n1554, 
                           SL => mult_21_C247_n48, Z => mult_21_C247_n922);
   mult_21_C247_U828 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n45, SL => mult_21_C247_n922, Z => 
                           mult_21_C247_n1225);
   mult_21_C247_U827 : MUXB2DL port map( A0 => mult_21_C247_n1549, A1 => n286, 
                           SL => mult_21_C247_n48, Z => mult_21_C247_n921);
   mult_21_C247_U826 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n45, SL => mult_21_C247_n921, Z => 
                           mult_21_C247_n1224);
   mult_21_C247_U825 : MUXB2DL port map( A0 => n282, A1 => mult_21_C247_n1549, 
                           SL => mult_21_C247_n48, Z => mult_21_C247_n920);
   mult_21_C247_U824 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n45, SL => mult_21_C247_n920, Z => 
                           mult_21_C247_n1223);
   mult_21_C247_U823 : MUXB2DL port map( A0 => n278, A1 => mult_21_C247_n1547, 
                           SL => mult_21_C247_n48, Z => mult_21_C247_n919);
   mult_21_C247_U822 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n45, SL => mult_21_C247_n919, Z => 
                           mult_21_C247_n1222);
   mult_21_C247_U821 : MUXB2DL port map( A0 => n279, A1 => n278, SL => 
                           mult_21_C247_n48, Z => mult_21_C247_n918);
   mult_21_C247_U820 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n45, SL => mult_21_C247_n918, Z => 
                           mult_21_C247_n1221);
   mult_21_C247_U819 : MUXB2DL port map( A0 => mult_21_C247_n1545, A1 => n279, 
                           SL => mult_21_C247_n48, Z => mult_21_C247_n917);
   mult_21_C247_U818 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n45, SL => mult_21_C247_n917, Z => 
                           mult_21_C247_n1220);
   mult_21_C247_U817 : MUXB2DL port map( A0 => n281, A1 => mult_21_C247_n1545, 
                           SL => mult_21_C247_n48, Z => mult_21_C247_n916);
   mult_21_C247_U816 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n45, SL => mult_21_C247_n916, Z => 
                           mult_21_C247_n1219);
   mult_21_C247_U815 : MUXB2DL port map( A0 => mult_21_C247_n1543, A1 => n281, 
                           SL => mult_21_C247_n48, Z => mult_21_C247_n915);
   mult_21_C247_U814 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n45, SL => mult_21_C247_n915, Z => 
                           mult_21_C247_n1218);
   mult_21_C247_U813 : MUXB2DL port map( A0 => n274, A1 => n285, SL => 
                           mult_21_C247_n48, Z => mult_21_C247_n914);
   mult_21_C247_U812 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n45, SL => mult_21_C247_n914, Z => 
                           mult_21_C247_n1217);
   mult_21_C247_U811 : MUXB2DL port map( A0 => n271, A1 => n274, SL => 
                           mult_21_C247_n48, Z => mult_21_C247_n913);
   mult_21_C247_U810 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n45, SL => mult_21_C247_n913, Z => 
                           mult_21_C247_n1216);
   mult_21_C247_U809 : MUXB2DL port map( A0 => n272, A1 => n271, SL => 
                           mult_21_C247_n48, Z => mult_21_C247_n912);
   mult_21_C247_U808 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n45, SL => mult_21_C247_n912, Z => 
                           mult_21_C247_n1215);
   mult_21_C247_U807 : MUXB2DL port map( A0 => n273, A1 => n272, SL => 
                           mult_21_C247_n48, Z => mult_21_C247_n911);
   mult_21_C247_U806 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n45, SL => mult_21_C247_n911, Z => 
                           mult_21_C247_n1214);
   mult_21_C247_U805 : MUXB2DL port map( A0 => n291, A1 => n273, SL => 
                           mult_21_C247_n48, Z => mult_21_C247_n910);
   mult_21_C247_U804 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n45, SL => mult_21_C247_n910, Z => 
                           mult_21_C247_n1213);
   mult_21_C247_U803 : MUXB2DL port map( A0 => n292, A1 => n291, SL => 
                           mult_21_C247_n48, Z => mult_21_C247_n909);
   mult_21_C247_U802 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n45, SL => mult_21_C247_n909, Z => 
                           mult_21_C247_n1212);
   mult_21_C247_U801 : MUXB2DL port map( A0 => n289, A1 => n292, SL => 
                           mult_21_C247_n48, Z => mult_21_C247_n908);
   mult_21_C247_U800 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n45, SL => mult_21_C247_n908, Z => 
                           mult_21_C247_n1211);
   mult_21_C247_U799 : MUXB2DL port map( A0 => n290, A1 => n289, SL => 
                           mult_21_C247_n48, Z => mult_21_C247_n907);
   mult_21_C247_U798 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n45, SL => mult_21_C247_n907, Z => 
                           mult_21_C247_n1210);
   mult_21_C247_U797 : MUXB2DL port map( A0 => n293, A1 => n290, SL => 
                           mult_21_C247_n48, Z => mult_21_C247_n906);
   mult_21_C247_U796 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n45, SL => mult_21_C247_n906, Z => 
                           mult_21_C247_n1209);
   mult_21_C247_U795 : MUXB2DL port map( A0 => n294, A1 => n293, SL => 
                           mult_21_C247_n48, Z => mult_21_C247_n905);
   mult_21_C247_U794 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n45, SL => mult_21_C247_n905, Z => 
                           mult_21_C247_n1208);
   mult_21_C247_U793 : MUXB2DL port map( A0 => n295, A1 => n294, SL => 
                           mult_21_C247_n48, Z => mult_21_C247_n904);
   mult_21_C247_U792 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n45, SL => mult_21_C247_n904, Z => 
                           mult_21_C247_n1207);
   mult_21_C247_U791 : NOR2M1D1 port map( A1 => mult_21_C247_n42, A2 => 
                           mult_21_C247_n45, Z => mult_21_C247_n1091);
   mult_21_C247_U790 : NAN2M1D1 port map( A1 => mult_21_C247_n56, A2 => 
                           mult_21_C247_n1556, Z => mult_21_C247_n903);
   mult_21_C247_U789 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n53, SL => mult_21_C247_n903, Z => 
                           mult_21_C247_n1206);
   mult_21_C247_U788 : MUXB2DL port map( A0 => n283, A1 => n288, SL => 
                           mult_21_C247_n56, Z => mult_21_C247_n902);
   mult_21_C247_U787 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n53, SL => mult_21_C247_n902, Z => 
                           mult_21_C247_n1205);
   mult_21_C247_U786 : MUXB2DL port map( A0 => mult_21_C247_n1553, A1 => n283, 
                           SL => mult_21_C247_n56, Z => mult_21_C247_n901);
   mult_21_C247_U785 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n53, SL => mult_21_C247_n901, Z => 
                           mult_21_C247_n1204);
   mult_21_C247_U784 : MUXB2DL port map( A0 => mult_21_C247_n1551, A1 => 
                           mult_21_C247_n1553, SL => mult_21_C247_n56, Z => 
                           mult_21_C247_n900);
   mult_21_C247_U783 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n53, SL => mult_21_C247_n900, Z => 
                           mult_21_C247_n1203);
   mult_21_C247_U782 : MUXB2DL port map( A0 => mult_21_C247_n1549, A1 => 
                           mult_21_C247_n1551, SL => mult_21_C247_n56, Z => 
                           mult_21_C247_n899);
   mult_21_C247_U781 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n53, SL => mult_21_C247_n899, Z => 
                           mult_21_C247_n1202);
   mult_21_C247_U780 : MUXB2DL port map( A0 => n282, A1 => mult_21_C247_n1549, 
                           SL => mult_21_C247_n56, Z => mult_21_C247_n898);
   mult_21_C247_U779 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n53, SL => mult_21_C247_n898, Z => 
                           mult_21_C247_n1201);
   mult_21_C247_U778 : MUXB2DL port map( A0 => n278, A1 => mult_21_C247_n1547, 
                           SL => mult_21_C247_n56, Z => mult_21_C247_n897);
   mult_21_C247_U777 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n53, SL => mult_21_C247_n897, Z => 
                           mult_21_C247_n1200);
   mult_21_C247_U776 : MUXB2DL port map( A0 => n279, A1 => n278, SL => 
                           mult_21_C247_n56, Z => mult_21_C247_n896);
   mult_21_C247_U775 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n53, SL => mult_21_C247_n896, Z => 
                           mult_21_C247_n1199);
   mult_21_C247_U774 : MUXB2DL port map( A0 => mult_21_C247_n1545, A1 => n279, 
                           SL => mult_21_C247_n56, Z => mult_21_C247_n895);
   mult_21_C247_U773 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n53, SL => mult_21_C247_n895, Z => 
                           mult_21_C247_n1198);
   mult_21_C247_U772 : MUXB2DL port map( A0 => n281, A1 => n280, SL => 
                           mult_21_C247_n56, Z => mult_21_C247_n894);
   mult_21_C247_U771 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n53, SL => mult_21_C247_n894, Z => 
                           mult_21_C247_n1197);
   mult_21_C247_U770 : MUXB2DL port map( A0 => mult_21_C247_n1543, A1 => n281, 
                           SL => mult_21_C247_n56, Z => mult_21_C247_n893);
   mult_21_C247_U769 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n53, SL => mult_21_C247_n893, Z => 
                           mult_21_C247_n1196);
   mult_21_C247_U768 : MUXB2DL port map( A0 => n274, A1 => n285, SL => 
                           mult_21_C247_n56, Z => mult_21_C247_n892);
   mult_21_C247_U767 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n53, SL => mult_21_C247_n892, Z => 
                           mult_21_C247_n1195);
   mult_21_C247_U766 : MUXB2DL port map( A0 => n271, A1 => n274, SL => 
                           mult_21_C247_n56, Z => mult_21_C247_n891);
   mult_21_C247_U765 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n53, SL => mult_21_C247_n891, Z => 
                           mult_21_C247_n1194);
   mult_21_C247_U764 : MUXB2DL port map( A0 => n272, A1 => n271, SL => 
                           mult_21_C247_n56, Z => mult_21_C247_n890);
   mult_21_C247_U763 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n53, SL => mult_21_C247_n890, Z => 
                           mult_21_C247_n1193);
   mult_21_C247_U762 : MUXB2DL port map( A0 => n273, A1 => n272, SL => 
                           mult_21_C247_n56, Z => mult_21_C247_n889);
   mult_21_C247_U761 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n53, SL => mult_21_C247_n889, Z => 
                           mult_21_C247_n1192);
   mult_21_C247_U760 : MUXB2DL port map( A0 => n291, A1 => n273, SL => 
                           mult_21_C247_n56, Z => mult_21_C247_n888);
   mult_21_C247_U759 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n53, SL => mult_21_C247_n888, Z => 
                           mult_21_C247_n1191);
   mult_21_C247_U758 : MUXB2DL port map( A0 => n292, A1 => n291, SL => 
                           mult_21_C247_n56, Z => mult_21_C247_n887);
   mult_21_C247_U757 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n53, SL => mult_21_C247_n887, Z => 
                           mult_21_C247_n1190);
   mult_21_C247_U756 : MUXB2DL port map( A0 => n289, A1 => n292, SL => 
                           mult_21_C247_n56, Z => mult_21_C247_n886);
   mult_21_C247_U755 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n53, SL => mult_21_C247_n886, Z => 
                           mult_21_C247_n1189);
   mult_21_C247_U754 : MUXB2DL port map( A0 => n290, A1 => n289, SL => 
                           mult_21_C247_n56, Z => mult_21_C247_n885);
   mult_21_C247_U753 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n53, SL => mult_21_C247_n885, Z => 
                           mult_21_C247_n1188);
   mult_21_C247_U752 : MUXB2DL port map( A0 => n293, A1 => n290, SL => 
                           mult_21_C247_n56, Z => mult_21_C247_n884);
   mult_21_C247_U751 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n53, SL => mult_21_C247_n884, Z => 
                           mult_21_C247_n1187);
   mult_21_C247_U750 : NOR2M1D1 port map( A1 => mult_21_C247_n50, A2 => 
                           mult_21_C247_n53, Z => mult_21_C247_n1090);
   mult_21_C247_U749 : NAN2M1D1 port map( A1 => mult_21_C247_n63, A2 => n288, Z
                           => mult_21_C247_n883);
   mult_21_C247_U748 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n61, SL => mult_21_C247_n883, Z => 
                           mult_21_C247_n1186);
   mult_21_C247_U747 : MUXB2DL port map( A0 => n283, A1 => mult_21_C247_n1556, 
                           SL => mult_21_C247_n63, Z => mult_21_C247_n882);
   mult_21_C247_U746 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n61, SL => mult_21_C247_n882, Z => 
                           mult_21_C247_n1185);
   mult_21_C247_U745 : MUXB2DL port map( A0 => mult_21_C247_n1553, A1 => n283, 
                           SL => mult_21_C247_n63, Z => mult_21_C247_n881);
   mult_21_C247_U744 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n61, SL => mult_21_C247_n881, Z => 
                           mult_21_C247_n1184);
   mult_21_C247_U743 : MUXB2DL port map( A0 => n286, A1 => mult_21_C247_n1554, 
                           SL => mult_21_C247_n63, Z => mult_21_C247_n880);
   mult_21_C247_U742 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n61, SL => mult_21_C247_n880, Z => 
                           mult_21_C247_n1183);
   mult_21_C247_U741 : MUXB2DL port map( A0 => mult_21_C247_n1549, A1 => 
                           mult_21_C247_n1551, SL => mult_21_C247_n63, Z => 
                           mult_21_C247_n879);
   mult_21_C247_U740 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n61, SL => mult_21_C247_n879, Z => 
                           mult_21_C247_n1182);
   mult_21_C247_U739 : MUXB2DL port map( A0 => mult_21_C247_n1547, A1 => n287, 
                           SL => mult_21_C247_n63, Z => mult_21_C247_n878);
   mult_21_C247_U738 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n61, SL => mult_21_C247_n878, Z => 
                           mult_21_C247_n1181);
   mult_21_C247_U737 : MUXB2DL port map( A0 => n278, A1 => mult_21_C247_n1547, 
                           SL => mult_21_C247_n63, Z => mult_21_C247_n877);
   mult_21_C247_U736 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n61, SL => mult_21_C247_n877, Z => 
                           mult_21_C247_n1180);
   mult_21_C247_U735 : MUXB2DL port map( A0 => n279, A1 => n278, SL => 
                           mult_21_C247_n63, Z => mult_21_C247_n876);
   mult_21_C247_U734 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n61, SL => mult_21_C247_n876, Z => 
                           mult_21_C247_n1179);
   mult_21_C247_U733 : MUXB2DL port map( A0 => mult_21_C247_n1545, A1 => n279, 
                           SL => mult_21_C247_n63, Z => mult_21_C247_n875);
   mult_21_C247_U732 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n61, SL => mult_21_C247_n875, Z => 
                           mult_21_C247_n1178);
   mult_21_C247_U731 : MUXB2DL port map( A0 => n281, A1 => mult_21_C247_n1545, 
                           SL => mult_21_C247_n63, Z => mult_21_C247_n874);
   mult_21_C247_U730 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n61, SL => mult_21_C247_n874, Z => 
                           mult_21_C247_n1177);
   mult_21_C247_U729 : MUXB2DL port map( A0 => mult_21_C247_n1543, A1 => n281, 
                           SL => mult_21_C247_n63, Z => mult_21_C247_n873);
   mult_21_C247_U728 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n61, SL => mult_21_C247_n873, Z => 
                           mult_21_C247_n1176);
   mult_21_C247_U727 : MUXB2DL port map( A0 => n274, A1 => mult_21_C247_n1543, 
                           SL => mult_21_C247_n63, Z => mult_21_C247_n872);
   mult_21_C247_U726 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n61, SL => mult_21_C247_n872, Z => 
                           mult_21_C247_n1175);
   mult_21_C247_U725 : MUXB2DL port map( A0 => n271, A1 => n274, SL => 
                           mult_21_C247_n63, Z => mult_21_C247_n871);
   mult_21_C247_U724 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n61, SL => mult_21_C247_n871, Z => 
                           mult_21_C247_n1174);
   mult_21_C247_U723 : MUXB2DL port map( A0 => n272, A1 => n271, SL => 
                           mult_21_C247_n63, Z => mult_21_C247_n870);
   mult_21_C247_U722 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n61, SL => mult_21_C247_n870, Z => 
                           mult_21_C247_n1173);
   mult_21_C247_U721 : MUXB2DL port map( A0 => n273, A1 => n272, SL => 
                           mult_21_C247_n63, Z => mult_21_C247_n869);
   mult_21_C247_U720 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n61, SL => mult_21_C247_n869, Z => 
                           mult_21_C247_n1172);
   mult_21_C247_U719 : MUXB2DL port map( A0 => n291, A1 => n273, SL => 
                           mult_21_C247_n63, Z => mult_21_C247_n868);
   mult_21_C247_U718 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n61, SL => mult_21_C247_n868, Z => 
                           mult_21_C247_n1171);
   mult_21_C247_U717 : MUXB2DL port map( A0 => n292, A1 => n291, SL => 
                           mult_21_C247_n63, Z => mult_21_C247_n867);
   mult_21_C247_U716 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n61, SL => mult_21_C247_n867, Z => 
                           mult_21_C247_n1170);
   mult_21_C247_U715 : MUXB2DL port map( A0 => n289, A1 => n292, SL => 
                           mult_21_C247_n63, Z => mult_21_C247_n866);
   mult_21_C247_U714 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n61, SL => mult_21_C247_n866, Z => 
                           mult_21_C247_n1169);
   mult_21_C247_U713 : NOR2M1D1 port map( A1 => mult_21_C247_n58, A2 => 
                           mult_21_C247_n61, Z => mult_21_C247_n1089);
   mult_21_C247_U712 : NAN2M1D1 port map( A1 => mult_21_C247_n71, A2 => 
                           mult_21_C247_n1556, Z => mult_21_C247_n865);
   mult_21_C247_U711 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n69, SL => mult_21_C247_n865, Z => 
                           mult_21_C247_n1168);
   mult_21_C247_U710 : MUXB2DL port map( A0 => n283, A1 => mult_21_C247_n1556, 
                           SL => mult_21_C247_n71, Z => mult_21_C247_n864);
   mult_21_C247_U709 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n69, SL => mult_21_C247_n864, Z => 
                           mult_21_C247_n1167);
   mult_21_C247_U708 : MUXB2DL port map( A0 => mult_21_C247_n1553, A1 => n283, 
                           SL => mult_21_C247_n71, Z => mult_21_C247_n863);
   mult_21_C247_U707 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n69, SL => mult_21_C247_n863, Z => 
                           mult_21_C247_n1166);
   mult_21_C247_U706 : MUXB2DL port map( A0 => mult_21_C247_n1551, A1 => 
                           mult_21_C247_n1554, SL => mult_21_C247_n71, Z => 
                           mult_21_C247_n862);
   mult_21_C247_U705 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n69, SL => mult_21_C247_n862, Z => 
                           mult_21_C247_n1165);
   mult_21_C247_U704 : MUXB2DL port map( A0 => n287, A1 => mult_21_C247_n1551, 
                           SL => mult_21_C247_n71, Z => mult_21_C247_n861);
   mult_21_C247_U703 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n69, SL => mult_21_C247_n861, Z => 
                           mult_21_C247_n1164);
   mult_21_C247_U702 : MUXB2DL port map( A0 => mult_21_C247_n1547, A1 => 
                           mult_21_C247_n1549, SL => mult_21_C247_n71, Z => 
                           mult_21_C247_n860);
   mult_21_C247_U701 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n69, SL => mult_21_C247_n860, Z => 
                           mult_21_C247_n1163);
   mult_21_C247_U700 : MUXB2DL port map( A0 => n278, A1 => mult_21_C247_n1547, 
                           SL => mult_21_C247_n71, Z => mult_21_C247_n859);
   mult_21_C247_U699 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n69, SL => mult_21_C247_n859, Z => 
                           mult_21_C247_n1162);
   mult_21_C247_U698 : MUXB2DL port map( A0 => n279, A1 => n278, SL => 
                           mult_21_C247_n71, Z => mult_21_C247_n858);
   mult_21_C247_U697 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n69, SL => mult_21_C247_n858, Z => 
                           mult_21_C247_n1161);
   mult_21_C247_U696 : MUXB2DL port map( A0 => mult_21_C247_n1545, A1 => n279, 
                           SL => mult_21_C247_n71, Z => mult_21_C247_n857);
   mult_21_C247_U695 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n69, SL => mult_21_C247_n857, Z => 
                           mult_21_C247_n1160);
   mult_21_C247_U694 : MUXB2DL port map( A0 => n281, A1 => n280, SL => 
                           mult_21_C247_n71, Z => mult_21_C247_n856);
   mult_21_C247_U693 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n69, SL => mult_21_C247_n856, Z => 
                           mult_21_C247_n1159);
   mult_21_C247_U692 : MUXB2DL port map( A0 => mult_21_C247_n1543, A1 => n281, 
                           SL => mult_21_C247_n71, Z => mult_21_C247_n855);
   mult_21_C247_U691 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n69, SL => mult_21_C247_n855, Z => 
                           mult_21_C247_n1158);
   mult_21_C247_U690 : MUXB2DL port map( A0 => n274, A1 => n285, SL => 
                           mult_21_C247_n71, Z => mult_21_C247_n854);
   mult_21_C247_U689 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n69, SL => mult_21_C247_n854, Z => 
                           mult_21_C247_n1157);
   mult_21_C247_U688 : MUXB2DL port map( A0 => n271, A1 => n274, SL => 
                           mult_21_C247_n71, Z => mult_21_C247_n853);
   mult_21_C247_U687 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n69, SL => mult_21_C247_n853, Z => 
                           mult_21_C247_n1156);
   mult_21_C247_U686 : MUXB2DL port map( A0 => n272, A1 => n271, SL => 
                           mult_21_C247_n71, Z => mult_21_C247_n852);
   mult_21_C247_U685 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n69, SL => mult_21_C247_n852, Z => 
                           mult_21_C247_n1155);
   mult_21_C247_U684 : MUXB2DL port map( A0 => n273, A1 => n272, SL => 
                           mult_21_C247_n71, Z => mult_21_C247_n851);
   mult_21_C247_U683 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n69, SL => mult_21_C247_n851, Z => 
                           mult_21_C247_n1154);
   mult_21_C247_U682 : MUXB2DL port map( A0 => n291, A1 => n273, SL => 
                           mult_21_C247_n71, Z => mult_21_C247_n850);
   mult_21_C247_U681 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n69, SL => mult_21_C247_n850, Z => 
                           mult_21_C247_n1153);
   mult_21_C247_U680 : NOR2M1D1 port map( A1 => mult_21_C247_n66, A2 => 
                           mult_21_C247_n69, Z => mult_21_C247_n1088);
   mult_21_C247_U679 : NAN2M1D1 port map( A1 => mult_21_C247_n78, A2 => 
                           mult_21_C247_n1556, Z => mult_21_C247_n849);
   mult_21_C247_U678 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n76, SL => mult_21_C247_n849, Z => 
                           mult_21_C247_n1152);
   mult_21_C247_U677 : MUXB2DL port map( A0 => n283, A1 => mult_21_C247_n1556, 
                           SL => mult_21_C247_n78, Z => mult_21_C247_n848);
   mult_21_C247_U676 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n76, SL => mult_21_C247_n848, Z => 
                           mult_21_C247_n1151);
   mult_21_C247_U675 : MUXB2DL port map( A0 => mult_21_C247_n1554, A1 => n283, 
                           SL => mult_21_C247_n78, Z => mult_21_C247_n847);
   mult_21_C247_U674 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n76, SL => mult_21_C247_n847, Z => 
                           mult_21_C247_n1150);
   mult_21_C247_U673 : MUXB2DL port map( A0 => mult_21_C247_n1551, A1 => 
                           mult_21_C247_n1554, SL => mult_21_C247_n78, Z => 
                           mult_21_C247_n846);
   mult_21_C247_U672 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n76, SL => mult_21_C247_n846, Z => 
                           mult_21_C247_n1149);
   mult_21_C247_U671 : MUXB2DL port map( A0 => mult_21_C247_n1549, A1 => 
                           mult_21_C247_n1551, SL => mult_21_C247_n78, Z => 
                           mult_21_C247_n845);
   mult_21_C247_U670 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n76, SL => mult_21_C247_n845, Z => 
                           mult_21_C247_n1148);
   mult_21_C247_U669 : MUXB2DL port map( A0 => n282, A1 => n287, SL => 
                           mult_21_C247_n78, Z => mult_21_C247_n844);
   mult_21_C247_U668 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n76, SL => mult_21_C247_n844, Z => 
                           mult_21_C247_n1147);
   mult_21_C247_U667 : MUXB2DL port map( A0 => n278, A1 => mult_21_C247_n1547, 
                           SL => mult_21_C247_n78, Z => mult_21_C247_n843);
   mult_21_C247_U666 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n76, SL => mult_21_C247_n843, Z => 
                           mult_21_C247_n1146);
   mult_21_C247_U665 : MUXB2DL port map( A0 => n279, A1 => n278, SL => 
                           mult_21_C247_n78, Z => mult_21_C247_n842);
   mult_21_C247_U664 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n76, SL => mult_21_C247_n842, Z => 
                           mult_21_C247_n1145);
   mult_21_C247_U663 : MUXB2DL port map( A0 => mult_21_C247_n1545, A1 => n279, 
                           SL => mult_21_C247_n78, Z => mult_21_C247_n841);
   mult_21_C247_U662 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n76, SL => mult_21_C247_n841, Z => 
                           mult_21_C247_n1144);
   mult_21_C247_U661 : MUXB2DL port map( A0 => n281, A1 => n280, SL => 
                           mult_21_C247_n78, Z => mult_21_C247_n840);
   mult_21_C247_U660 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n76, SL => mult_21_C247_n840, Z => 
                           mult_21_C247_n1143);
   mult_21_C247_U659 : MUXB2DL port map( A0 => mult_21_C247_n1543, A1 => n281, 
                           SL => mult_21_C247_n78, Z => mult_21_C247_n839);
   mult_21_C247_U658 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n76, SL => mult_21_C247_n839, Z => 
                           mult_21_C247_n1142);
   mult_21_C247_U657 : MUXB2DL port map( A0 => n274, A1 => mult_21_C247_n1543, 
                           SL => mult_21_C247_n78, Z => mult_21_C247_n838);
   mult_21_C247_U656 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n76, SL => mult_21_C247_n838, Z => 
                           mult_21_C247_n1141);
   mult_21_C247_U655 : MUXB2DL port map( A0 => n271, A1 => n274, SL => 
                           mult_21_C247_n78, Z => mult_21_C247_n837);
   mult_21_C247_U654 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n76, SL => mult_21_C247_n837, Z => 
                           mult_21_C247_n1140);
   mult_21_C247_U653 : MUXB2DL port map( A0 => n272, A1 => n271, SL => 
                           mult_21_C247_n78, Z => mult_21_C247_n836);
   mult_21_C247_U652 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n76, SL => mult_21_C247_n836, Z => 
                           mult_21_C247_n1139);
   mult_21_C247_U651 : NOR2M1D1 port map( A1 => mult_21_C247_n73, A2 => 
                           mult_21_C247_n76, Z => mult_21_C247_n1087);
   mult_21_C247_U650 : NAN2M1D1 port map( A1 => mult_21_C247_n83, A2 => n288, Z
                           => mult_21_C247_n835);
   mult_21_C247_U649 : MUXB2DL port map( A0 => mult_21_C247_n79, A1 => 
                           mult_21_C247_n81, SL => mult_21_C247_n835, Z => 
                           mult_21_C247_n1138);
   mult_21_C247_U648 : MUXB2DL port map( A0 => n283, A1 => mult_21_C247_n1556, 
                           SL => mult_21_C247_n83, Z => mult_21_C247_n834);
   mult_21_C247_U647 : MUXB2DL port map( A0 => mult_21_C247_n79, A1 => 
                           mult_21_C247_n81, SL => mult_21_C247_n834, Z => 
                           mult_21_C247_n1137);
   mult_21_C247_U646 : MUXB2DL port map( A0 => mult_21_C247_n1554, A1 => n283, 
                           SL => mult_21_C247_n83, Z => mult_21_C247_n833);
   mult_21_C247_U645 : MUXB2DL port map( A0 => mult_21_C247_n79, A1 => 
                           mult_21_C247_n81, SL => mult_21_C247_n833, Z => 
                           mult_21_C247_n1136);
   mult_21_C247_U644 : MUXB2DL port map( A0 => mult_21_C247_n1551, A1 => 
                           mult_21_C247_n1554, SL => mult_21_C247_n83, Z => 
                           mult_21_C247_n832);
   mult_21_C247_U643 : MUXB2DL port map( A0 => mult_21_C247_n79, A1 => 
                           mult_21_C247_n81, SL => mult_21_C247_n832, Z => 
                           mult_21_C247_n1135);
   mult_21_C247_U642 : MUXB2DL port map( A0 => mult_21_C247_n1549, A1 => 
                           mult_21_C247_n1551, SL => mult_21_C247_n83, Z => 
                           mult_21_C247_n831);
   mult_21_C247_U641 : MUXB2DL port map( A0 => mult_21_C247_n79, A1 => 
                           mult_21_C247_n81, SL => mult_21_C247_n831, Z => 
                           mult_21_C247_n1134);
   mult_21_C247_U640 : MUXB2DL port map( A0 => n282, A1 => n287, SL => 
                           mult_21_C247_n83, Z => mult_21_C247_n830);
   mult_21_C247_U639 : MUXB2DL port map( A0 => mult_21_C247_n79, A1 => 
                           mult_21_C247_n81, SL => mult_21_C247_n830, Z => 
                           mult_21_C247_n1133);
   mult_21_C247_U638 : MUXB2DL port map( A0 => n278, A1 => mult_21_C247_n1547, 
                           SL => mult_21_C247_n83, Z => mult_21_C247_n829);
   mult_21_C247_U637 : MUXB2DL port map( A0 => mult_21_C247_n79, A1 => 
                           mult_21_C247_n81, SL => mult_21_C247_n829, Z => 
                           mult_21_C247_n1132);
   mult_21_C247_U636 : MUXB2DL port map( A0 => n279, A1 => n278, SL => 
                           mult_21_C247_n83, Z => mult_21_C247_n828);
   mult_21_C247_U635 : MUXB2DL port map( A0 => mult_21_C247_n79, A1 => 
                           mult_21_C247_n81, SL => mult_21_C247_n828, Z => 
                           mult_21_C247_n1131);
   mult_21_C247_U634 : MUXB2DL port map( A0 => mult_21_C247_n1545, A1 => n279, 
                           SL => mult_21_C247_n83, Z => mult_21_C247_n827);
   mult_21_C247_U633 : MUXB2DL port map( A0 => mult_21_C247_n79, A1 => 
                           mult_21_C247_n81, SL => mult_21_C247_n827, Z => 
                           mult_21_C247_n1130);
   mult_21_C247_U632 : MUXB2DL port map( A0 => n281, A1 => n280, SL => 
                           mult_21_C247_n83, Z => mult_21_C247_n826);
   mult_21_C247_U631 : MUXB2DL port map( A0 => mult_21_C247_n79, A1 => 
                           mult_21_C247_n81, SL => mult_21_C247_n826, Z => 
                           mult_21_C247_n1129);
   mult_21_C247_U630 : MUXB2DL port map( A0 => mult_21_C247_n1543, A1 => n281, 
                           SL => mult_21_C247_n83, Z => mult_21_C247_n825);
   mult_21_C247_U629 : MUXB2DL port map( A0 => mult_21_C247_n79, A1 => 
                           mult_21_C247_n81, SL => mult_21_C247_n825, Z => 
                           mult_21_C247_n1128);
   mult_21_C247_U628 : MUXB2DL port map( A0 => n274, A1 => n285, SL => 
                           mult_21_C247_n83, Z => mult_21_C247_n824);
   mult_21_C247_U627 : MUXB2DL port map( A0 => mult_21_C247_n79, A1 => 
                           mult_21_C247_n81, SL => mult_21_C247_n824, Z => 
                           mult_21_C247_n1127);
   mult_21_C247_U626 : NOR2M1D1 port map( A1 => mult_21_C247_n79, A2 => 
                           mult_21_C247_n81, Z => mult_21_C247_n1086);
   mult_21_C247_U625 : NAN2M1D1 port map( A1 => mult_21_C247_n88, A2 => 
                           mult_21_C247_n1556, Z => mult_21_C247_n823);
   mult_21_C247_U624 : MUXB2DL port map( A0 => mult_21_C247_n84, A1 => 
                           mult_21_C247_n86, SL => mult_21_C247_n823, Z => 
                           mult_21_C247_n1126);
   mult_21_C247_U623 : MUXB2DL port map( A0 => n283, A1 => mult_21_C247_n1556, 
                           SL => mult_21_C247_n88, Z => mult_21_C247_n822);
   mult_21_C247_U622 : MUXB2DL port map( A0 => mult_21_C247_n84, A1 => 
                           mult_21_C247_n86, SL => mult_21_C247_n822, Z => 
                           mult_21_C247_n1125);
   mult_21_C247_U621 : MUXB2DL port map( A0 => mult_21_C247_n1553, A1 => n283, 
                           SL => mult_21_C247_n88, Z => mult_21_C247_n821);
   mult_21_C247_U620 : MUXB2DL port map( A0 => mult_21_C247_n84, A1 => 
                           mult_21_C247_n86, SL => mult_21_C247_n821, Z => 
                           mult_21_C247_n1124);
   mult_21_C247_U619 : MUXB2DL port map( A0 => n286, A1 => mult_21_C247_n1554, 
                           SL => mult_21_C247_n88, Z => mult_21_C247_n820);
   mult_21_C247_U618 : MUXB2DL port map( A0 => mult_21_C247_n84, A1 => 
                           mult_21_C247_n86, SL => mult_21_C247_n820, Z => 
                           mult_21_C247_n1123);
   mult_21_C247_U617 : MUXB2DL port map( A0 => mult_21_C247_n1549, A1 => 
                           mult_21_C247_n1551, SL => mult_21_C247_n88, Z => 
                           mult_21_C247_n819);
   mult_21_C247_U616 : MUXB2DL port map( A0 => mult_21_C247_n84, A1 => 
                           mult_21_C247_n86, SL => mult_21_C247_n819, Z => 
                           mult_21_C247_n1122);
   mult_21_C247_U615 : MUXB2DL port map( A0 => n282, A1 => n287, SL => 
                           mult_21_C247_n88, Z => mult_21_C247_n818);
   mult_21_C247_U614 : MUXB2DL port map( A0 => mult_21_C247_n84, A1 => 
                           mult_21_C247_n86, SL => mult_21_C247_n818, Z => 
                           mult_21_C247_n1121);
   mult_21_C247_U613 : MUXB2DL port map( A0 => n278, A1 => mult_21_C247_n1547, 
                           SL => mult_21_C247_n88, Z => mult_21_C247_n817);
   mult_21_C247_U612 : MUXB2DL port map( A0 => mult_21_C247_n84, A1 => 
                           mult_21_C247_n86, SL => mult_21_C247_n817, Z => 
                           mult_21_C247_n1120);
   mult_21_C247_U611 : MUXB2DL port map( A0 => n279, A1 => n278, SL => 
                           mult_21_C247_n88, Z => mult_21_C247_n816);
   mult_21_C247_U610 : MUXB2DL port map( A0 => mult_21_C247_n84, A1 => 
                           mult_21_C247_n86, SL => mult_21_C247_n816, Z => 
                           mult_21_C247_n1119);
   mult_21_C247_U609 : MUXB2DL port map( A0 => mult_21_C247_n1545, A1 => n279, 
                           SL => mult_21_C247_n88, Z => mult_21_C247_n815);
   mult_21_C247_U608 : MUXB2DL port map( A0 => mult_21_C247_n84, A1 => 
                           mult_21_C247_n86, SL => mult_21_C247_n815, Z => 
                           mult_21_C247_n1118);
   mult_21_C247_U607 : MUXB2DL port map( A0 => n281, A1 => n280, SL => 
                           mult_21_C247_n88, Z => mult_21_C247_n814);
   mult_21_C247_U606 : MUXB2DL port map( A0 => mult_21_C247_n84, A1 => 
                           mult_21_C247_n86, SL => mult_21_C247_n814, Z => 
                           mult_21_C247_n1117);
   mult_21_C247_U605 : NOR2M1D1 port map( A1 => mult_21_C247_n84, A2 => 
                           mult_21_C247_n86, Z => mult_21_C247_n1085);
   mult_21_C247_U604 : NAN2M1D1 port map( A1 => mult_21_C247_n93, A2 => 
                           mult_21_C247_n1556, Z => mult_21_C247_n813);
   mult_21_C247_U603 : MUXB2DL port map( A0 => mult_21_C247_n89, A1 => 
                           mult_21_C247_n91, SL => mult_21_C247_n813, Z => 
                           mult_21_C247_n1116);
   mult_21_C247_U602 : MUXB2DL port map( A0 => n283, A1 => mult_21_C247_n1556, 
                           SL => mult_21_C247_n93, Z => mult_21_C247_n812);
   mult_21_C247_U601 : MUXB2DL port map( A0 => mult_21_C247_n89, A1 => 
                           mult_21_C247_n91, SL => mult_21_C247_n812, Z => 
                           mult_21_C247_n1115);
   mult_21_C247_U600 : MUXB2DL port map( A0 => mult_21_C247_n1553, A1 => n283, 
                           SL => mult_21_C247_n93, Z => mult_21_C247_n811);
   mult_21_C247_U599 : MUXB2DL port map( A0 => mult_21_C247_n89, A1 => 
                           mult_21_C247_n91, SL => mult_21_C247_n811, Z => 
                           mult_21_C247_n1114);
   mult_21_C247_U598 : MUXB2DL port map( A0 => n286, A1 => mult_21_C247_n1554, 
                           SL => mult_21_C247_n93, Z => mult_21_C247_n810);
   mult_21_C247_U597 : MUXB2DL port map( A0 => mult_21_C247_n89, A1 => 
                           mult_21_C247_n91, SL => mult_21_C247_n810, Z => 
                           mult_21_C247_n1113);
   mult_21_C247_U596 : MUXB2DL port map( A0 => mult_21_C247_n1549, A1 => 
                           mult_21_C247_n1551, SL => mult_21_C247_n93, Z => 
                           mult_21_C247_n809);
   mult_21_C247_U595 : MUXB2DL port map( A0 => mult_21_C247_n89, A1 => 
                           mult_21_C247_n91, SL => mult_21_C247_n809, Z => 
                           mult_21_C247_n1112);
   mult_21_C247_U594 : MUXB2DL port map( A0 => n282, A1 => n287, SL => 
                           mult_21_C247_n93, Z => mult_21_C247_n808);
   mult_21_C247_U593 : MUXB2DL port map( A0 => mult_21_C247_n89, A1 => 
                           mult_21_C247_n91, SL => mult_21_C247_n808, Z => 
                           mult_21_C247_n1111);
   mult_21_C247_U592 : MUXB2DL port map( A0 => n278, A1 => mult_21_C247_n1547, 
                           SL => mult_21_C247_n93, Z => mult_21_C247_n807);
   mult_21_C247_U591 : MUXB2DL port map( A0 => mult_21_C247_n89, A1 => 
                           mult_21_C247_n91, SL => mult_21_C247_n807, Z => 
                           mult_21_C247_n1110);
   mult_21_C247_U590 : MUXB2DL port map( A0 => n279, A1 => n278, SL => 
                           mult_21_C247_n93, Z => mult_21_C247_n806);
   mult_21_C247_U589 : MUXB2DL port map( A0 => mult_21_C247_n89, A1 => 
                           mult_21_C247_n91, SL => mult_21_C247_n806, Z => 
                           mult_21_C247_n1109);
   mult_21_C247_U588 : NOR2M1D1 port map( A1 => mult_21_C247_n89, A2 => 
                           mult_21_C247_n91, Z => mult_21_C247_n1084);
   mult_21_C247_U587 : NAN2M1D1 port map( A1 => mult_21_C247_n98, A2 => n288, Z
                           => mult_21_C247_n805);
   mult_21_C247_U586 : MUXB2DL port map( A0 => mult_21_C247_n94, A1 => 
                           mult_21_C247_n96, SL => mult_21_C247_n805, Z => 
                           mult_21_C247_n1108);
   mult_21_C247_U585 : MUXB2DL port map( A0 => n283, A1 => mult_21_C247_n1556, 
                           SL => mult_21_C247_n98, Z => mult_21_C247_n804);
   mult_21_C247_U584 : MUXB2DL port map( A0 => mult_21_C247_n94, A1 => 
                           mult_21_C247_n96, SL => mult_21_C247_n804, Z => 
                           mult_21_C247_n1107);
   mult_21_C247_U583 : MUXB2DL port map( A0 => mult_21_C247_n1553, A1 => n283, 
                           SL => mult_21_C247_n98, Z => mult_21_C247_n803);
   mult_21_C247_U582 : MUXB2DL port map( A0 => mult_21_C247_n94, A1 => 
                           mult_21_C247_n96, SL => mult_21_C247_n803, Z => 
                           mult_21_C247_n1106);
   mult_21_C247_U581 : MUXB2DL port map( A0 => n286, A1 => mult_21_C247_n1554, 
                           SL => mult_21_C247_n98, Z => mult_21_C247_n802);
   mult_21_C247_U580 : MUXB2DL port map( A0 => mult_21_C247_n94, A1 => 
                           mult_21_C247_n96, SL => mult_21_C247_n802, Z => 
                           mult_21_C247_n1105);
   mult_21_C247_U579 : MUXB2DL port map( A0 => mult_21_C247_n1549, A1 => 
                           mult_21_C247_n1551, SL => mult_21_C247_n98, Z => 
                           mult_21_C247_n801);
   mult_21_C247_U578 : MUXB2DL port map( A0 => mult_21_C247_n94, A1 => 
                           mult_21_C247_n96, SL => mult_21_C247_n801, Z => 
                           mult_21_C247_n1104);
   mult_21_C247_U577 : MUXB2DL port map( A0 => n282, A1 => n287, SL => 
                           mult_21_C247_n98, Z => mult_21_C247_n800);
   mult_21_C247_U576 : MUXB2DL port map( A0 => mult_21_C247_n94, A1 => 
                           mult_21_C247_n96, SL => mult_21_C247_n800, Z => 
                           mult_21_C247_n1103);
   mult_21_C247_U575 : NOR2M1D1 port map( A1 => mult_21_C247_n94, A2 => 
                           mult_21_C247_n96, Z => mult_21_C247_n1083);
   mult_21_C247_U574 : NAN2M1D1 port map( A1 => mult_21_C247_n103, A2 => n288, 
                           Z => mult_21_C247_n799);
   mult_21_C247_U573 : MUXB2DL port map( A0 => mult_21_C247_n99, A1 => 
                           mult_21_C247_n101, SL => mult_21_C247_n799, Z => 
                           mult_21_C247_n1102);
   mult_21_C247_U572 : MUXB2DL port map( A0 => n283, A1 => mult_21_C247_n1556, 
                           SL => mult_21_C247_n103, Z => mult_21_C247_n798);
   mult_21_C247_U571 : MUXB2DL port map( A0 => mult_21_C247_n99, A1 => 
                           mult_21_C247_n101, SL => mult_21_C247_n798, Z => 
                           mult_21_C247_n1101);
   mult_21_C247_U570 : MUXB2DL port map( A0 => mult_21_C247_n1553, A1 => n283, 
                           SL => mult_21_C247_n103, Z => mult_21_C247_n797);
   mult_21_C247_U569 : MUXB2DL port map( A0 => mult_21_C247_n99, A1 => 
                           mult_21_C247_n101, SL => mult_21_C247_n797, Z => 
                           mult_21_C247_n1100);
   mult_21_C247_U568 : MUXB2DL port map( A0 => n286, A1 => mult_21_C247_n1554, 
                           SL => mult_21_C247_n103, Z => mult_21_C247_n796);
   mult_21_C247_U567 : MUXB2DL port map( A0 => mult_21_C247_n99, A1 => 
                           mult_21_C247_n101, SL => mult_21_C247_n796, Z => 
                           mult_21_C247_n1099);
   mult_21_C247_U566 : NOR2M1D1 port map( A1 => mult_21_C247_n99, A2 => 
                           mult_21_C247_n101, Z => mult_21_C247_n1082);
   mult_21_C247_U565 : NAN2M1D1 port map( A1 => mult_21_C247_n106, A2 => n288, 
                           Z => mult_21_C247_n795);
   mult_21_C247_U564 : MUXB2DL port map( A0 => mult_21_C247_n104, A1 => 
                           mult_21_C247_n105, SL => mult_21_C247_n795, Z => 
                           mult_21_C247_n1098);
   mult_21_C247_U563 : MUXB2DL port map( A0 => n283, A1 => mult_21_C247_n1556, 
                           SL => mult_21_C247_n106, Z => mult_21_C247_n794);
   mult_21_C247_U562 : MUXB2DL port map( A0 => mult_21_C247_n104, A1 => 
                           mult_21_C247_n105, SL => mult_21_C247_n794, Z => 
                           mult_21_C247_n1097);
   mult_21_C247_U561 : NOR2M1D1 port map( A1 => mult_21_C247_n104, A2 => 
                           mult_21_C247_n105, Z => mult_21_C247_n1081);
   mult_21_C247_U557 : ADFULD1 port map( A => mult_21_C247_n1334, B => 
                           mult_21_C247_n1364, CI => mult_21_C247_n790, CO => 
                           mult_21_C247_n786, S => mult_21_C247_n787);
   mult_21_C247_U555 : ADFULD1 port map( A => mult_21_C247_n788, B => 
                           mult_21_C247_n1305, CI => mult_21_C247_n785, CO => 
                           mult_21_C247_n782, S => mult_21_C247_n783);
   mult_21_C247_U553 : ADFULD1 port map( A => mult_21_C247_n1304, B => 
                           mult_21_C247_n1362, CI => mult_21_C247_n1332, CO => 
                           mult_21_C247_n778, S => mult_21_C247_n779);
   mult_21_C247_U552 : ADFULD1 port map( A => mult_21_C247_n781, B => 
                           mult_21_C247_n784, CI => mult_21_C247_n779, CO => 
                           mult_21_C247_n776, S => mult_21_C247_n777);
   mult_21_C247_U550 : ADFULD1 port map( A => mult_21_C247_n1277, B => 
                           mult_21_C247_n1303, CI => mult_21_C247_n780, CO => 
                           mult_21_C247_n772, S => mult_21_C247_n773);
   mult_21_C247_U549 : ADFULD1 port map( A => mult_21_C247_n778, B => 
                           mult_21_C247_n775, CI => mult_21_C247_n773, CO => 
                           mult_21_C247_n770, S => mult_21_C247_n771);
   mult_21_C247_U547 : ADFULD1 port map( A => mult_21_C247_n1276, B => 
                           mult_21_C247_n1360, CI => mult_21_C247_n1330, CO => 
                           mult_21_C247_n766, S => mult_21_C247_n767);
   mult_21_C247_U546 : ADFULD1 port map( A => mult_21_C247_n774, B => 
                           mult_21_C247_n1302, CI => mult_21_C247_n769, CO => 
                           mult_21_C247_n764, S => mult_21_C247_n765);
   mult_21_C247_U545 : ADFULD1 port map( A => mult_21_C247_n767, B => 
                           mult_21_C247_n772, CI => mult_21_C247_n765, CO => 
                           mult_21_C247_n762, S => mult_21_C247_n763);
   mult_21_C247_U543 : ADFULD1 port map( A => mult_21_C247_n1275, B => 
                           mult_21_C247_n1301, CI => mult_21_C247_n1251, CO => 
                           mult_21_C247_n758, S => mult_21_C247_n759);
   mult_21_C247_U542 : ADFULD1 port map( A => mult_21_C247_n761, B => 
                           mult_21_C247_n768, CI => mult_21_C247_n766, CO => 
                           mult_21_C247_n756, S => mult_21_C247_n757);
   mult_21_C247_U541 : ADFULD1 port map( A => mult_21_C247_n764, B => 
                           mult_21_C247_n759, CI => mult_21_C247_n757, CO => 
                           mult_21_C247_n754, S => mult_21_C247_n755);
   mult_21_C247_U539 : ADFULD1 port map( A => mult_21_C247_n1250, B => 
                           mult_21_C247_n1358, CI => mult_21_C247_n1328, CO => 
                           mult_21_C247_n750, S => mult_21_C247_n751);
   mult_21_C247_U538 : ADFULD1 port map( A => mult_21_C247_n1274, B => 
                           mult_21_C247_n1300, CI => mult_21_C247_n760, CO => 
                           mult_21_C247_n748, S => mult_21_C247_n749);
   mult_21_C247_U537 : ADFULD1 port map( A => mult_21_C247_n758, B => 
                           mult_21_C247_n753, CI => mult_21_C247_n751, CO => 
                           mult_21_C247_n746, S => mult_21_C247_n747);
   mult_21_C247_U536 : ADFULD1 port map( A => mult_21_C247_n756, B => 
                           mult_21_C247_n749, CI => mult_21_C247_n747, CO => 
                           mult_21_C247_n744, S => mult_21_C247_n745);
   mult_21_C247_U534 : ADFULD1 port map( A => mult_21_C247_n1273, B => 
                           mult_21_C247_n1249, CI => mult_21_C247_n1227, CO => 
                           mult_21_C247_n740, S => mult_21_C247_n741);
   mult_21_C247_U533 : ADFULD1 port map( A => mult_21_C247_n752, B => 
                           mult_21_C247_n1299, CI => mult_21_C247_n743, CO => 
                           mult_21_C247_n738, S => mult_21_C247_n739);
   mult_21_C247_U532 : ADFULD1 port map( A => mult_21_C247_n748, B => 
                           mult_21_C247_n750, CI => mult_21_C247_n741, CO => 
                           mult_21_C247_n736, S => mult_21_C247_n737);
   mult_21_C247_U531 : ADFULD1 port map( A => mult_21_C247_n746, B => 
                           mult_21_C247_n739, CI => mult_21_C247_n737, CO => 
                           mult_21_C247_n734, S => mult_21_C247_n735);
   mult_21_C247_U529 : ADFULD1 port map( A => mult_21_C247_n1248, B => 
                           mult_21_C247_n1356, CI => mult_21_C247_n1326, CO => 
                           mult_21_C247_n730, S => mult_21_C247_n731);
   mult_21_C247_U528 : ADFULD1 port map( A => mult_21_C247_n1272, B => 
                           mult_21_C247_n1298, CI => mult_21_C247_n1226, CO => 
                           mult_21_C247_n728, S => mult_21_C247_n729);
   mult_21_C247_U527 : ADFULD1 port map( A => mult_21_C247_n733, B => 
                           mult_21_C247_n742, CI => mult_21_C247_n740, CO => 
                           mult_21_C247_n726, S => mult_21_C247_n727);
   mult_21_C247_U526 : ADFULD1 port map( A => mult_21_C247_n729, B => 
                           mult_21_C247_n731, CI => mult_21_C247_n738, CO => 
                           mult_21_C247_n724, S => mult_21_C247_n725);
   mult_21_C247_U525 : ADFULD1 port map( A => mult_21_C247_n736, B => 
                           mult_21_C247_n727, CI => mult_21_C247_n725, CO => 
                           mult_21_C247_n722, S => mult_21_C247_n723);
   mult_21_C247_U523 : ADFULD1 port map( A => mult_21_C247_n1205, B => 
                           mult_21_C247_n1297, CI => mult_21_C247_n1225, CO => 
                           mult_21_C247_n718, S => mult_21_C247_n719);
   mult_21_C247_U522 : ADFULD1 port map( A => mult_21_C247_n1247, B => 
                           mult_21_C247_n1271, CI => mult_21_C247_n732, CO => 
                           mult_21_C247_n716, S => mult_21_C247_n717);
   mult_21_C247_U521 : ADFULD1 port map( A => mult_21_C247_n730, B => 
                           mult_21_C247_n721, CI => mult_21_C247_n728, CO => 
                           mult_21_C247_n714, S => mult_21_C247_n715);
   mult_21_C247_U520 : ADFULD1 port map( A => mult_21_C247_n717, B => 
                           mult_21_C247_n719, CI => mult_21_C247_n726, CO => 
                           mult_21_C247_n712, S => mult_21_C247_n713);
   mult_21_C247_U519 : ADFULD1 port map( A => mult_21_C247_n724, B => 
                           mult_21_C247_n715, CI => mult_21_C247_n713, CO => 
                           mult_21_C247_n710, S => mult_21_C247_n711);
   mult_21_C247_U517 : ADFULD1 port map( A => mult_21_C247_n1204, B => 
                           mult_21_C247_n1354, CI => mult_21_C247_n1324, CO => 
                           mult_21_C247_n706, S => mult_21_C247_n707);
   mult_21_C247_U516 : ADFULD1 port map( A => mult_21_C247_n1246, B => 
                           mult_21_C247_n1296, CI => mult_21_C247_n1224, CO => 
                           mult_21_C247_n704, S => mult_21_C247_n705);
   mult_21_C247_U515 : ADFULD1 port map( A => mult_21_C247_n720, B => 
                           mult_21_C247_n1270, CI => mult_21_C247_n709, CO => 
                           mult_21_C247_n702, S => mult_21_C247_n703);
   mult_21_C247_U514 : ADFULD1 port map( A => mult_21_C247_n716, B => 
                           mult_21_C247_n718, CI => mult_21_C247_n707, CO => 
                           mult_21_C247_n700, S => mult_21_C247_n701);
   mult_21_C247_U513 : ADFULD1 port map( A => mult_21_C247_n703, B => 
                           mult_21_C247_n705, CI => mult_21_C247_n714, CO => 
                           mult_21_C247_n698, S => mult_21_C247_n699);
   mult_21_C247_U512 : ADFULD1 port map( A => mult_21_C247_n712, B => 
                           mult_21_C247_n701, CI => mult_21_C247_n699, CO => 
                           mult_21_C247_n696, S => mult_21_C247_n697);
   mult_21_C247_U510 : ADFULD1 port map( A => mult_21_C247_n1185, B => 
                           mult_21_C247_n1269, CI => mult_21_C247_n1223, CO => 
                           mult_21_C247_n692, S => mult_21_C247_n693);
   mult_21_C247_U509 : ADFULD1 port map( A => mult_21_C247_n1203, B => 
                           mult_21_C247_n1295, CI => mult_21_C247_n1245, CO => 
                           mult_21_C247_n690, S => mult_21_C247_n691);
   mult_21_C247_U508 : ADFULD1 port map( A => mult_21_C247_n695, B => 
                           mult_21_C247_n708, CI => mult_21_C247_n706, CO => 
                           mult_21_C247_n688, S => mult_21_C247_n689);
   mult_21_C247_U507 : ADFULD1 port map( A => mult_21_C247_n691, B => 
                           mult_21_C247_n704, CI => mult_21_C247_n693, CO => 
                           mult_21_C247_n686, S => mult_21_C247_n687);
   mult_21_C247_U506 : ADFULD1 port map( A => mult_21_C247_n700, B => 
                           mult_21_C247_n702, CI => mult_21_C247_n689, CO => 
                           mult_21_C247_n684, S => mult_21_C247_n685);
   mult_21_C247_U505 : ADFULD1 port map( A => mult_21_C247_n698, B => 
                           mult_21_C247_n687, CI => mult_21_C247_n685, CO => 
                           mult_21_C247_n682, S => mult_21_C247_n683);
   mult_21_C247_U503 : ADFULD1 port map( A => mult_21_C247_n1202, B => 
                           mult_21_C247_n1352, CI => mult_21_C247_n1322, CO => 
                           mult_21_C247_n678, S => mult_21_C247_n679);
   mult_21_C247_U502 : ADFULD1 port map( A => mult_21_C247_n1184, B => 
                           mult_21_C247_n1268, CI => mult_21_C247_n1222, CO => 
                           mult_21_C247_n676, S => mult_21_C247_n677);
   mult_21_C247_U501 : ADFULD1 port map( A => mult_21_C247_n1244, B => 
                           mult_21_C247_n1294, CI => mult_21_C247_n694, CO => 
                           mult_21_C247_n674, S => mult_21_C247_n675);
   mult_21_C247_U500 : ADFULD1 port map( A => mult_21_C247_n692, B => 
                           mult_21_C247_n681, CI => mult_21_C247_n690, CO => 
                           mult_21_C247_n672, S => mult_21_C247_n673);
   mult_21_C247_U499 : ADFULD1 port map( A => mult_21_C247_n677, B => 
                           mult_21_C247_n679, CI => mult_21_C247_n675, CO => 
                           mult_21_C247_n670, S => mult_21_C247_n671);
   mult_21_C247_U498 : ADFULD1 port map( A => mult_21_C247_n686, B => 
                           mult_21_C247_n688, CI => mult_21_C247_n673, CO => 
                           mult_21_C247_n668, S => mult_21_C247_n669);
   mult_21_C247_U497 : ADFULD1 port map( A => mult_21_C247_n684, B => 
                           mult_21_C247_n671, CI => mult_21_C247_n669, CO => 
                           mult_21_C247_n666, S => mult_21_C247_n667);
   mult_21_C247_U495 : ADFULD1 port map( A => mult_21_C247_n1167, B => 
                           mult_21_C247_n1201, CI => mult_21_C247_n1221, CO => 
                           mult_21_C247_n662, S => mult_21_C247_n663);
   mult_21_C247_U494 : ADFULD1 port map( A => mult_21_C247_n1243, B => 
                           mult_21_C247_n1183, CI => mult_21_C247_n1267, CO => 
                           mult_21_C247_n660, S => mult_21_C247_n661);
   mult_21_C247_U493 : ADFULD1 port map( A => mult_21_C247_n680, B => 
                           mult_21_C247_n1293, CI => mult_21_C247_n665, CO => 
                           mult_21_C247_n658, S => mult_21_C247_n659);
   mult_21_C247_U492 : ADFULD1 port map( A => mult_21_C247_n676, B => 
                           mult_21_C247_n678, CI => mult_21_C247_n674, CO => 
                           mult_21_C247_n656, S => mult_21_C247_n657);
   mult_21_C247_U491 : ADFULD1 port map( A => mult_21_C247_n663, B => 
                           mult_21_C247_n661, CI => mult_21_C247_n672, CO => 
                           mult_21_C247_n654, S => mult_21_C247_n655);
   mult_21_C247_U490 : ADFULD1 port map( A => mult_21_C247_n670, B => 
                           mult_21_C247_n659, CI => mult_21_C247_n657, CO => 
                           mult_21_C247_n652, S => mult_21_C247_n653);
   mult_21_C247_U489 : ADFULD1 port map( A => mult_21_C247_n668, B => 
                           mult_21_C247_n655, CI => mult_21_C247_n653, CO => 
                           mult_21_C247_n650, S => mult_21_C247_n651);
   mult_21_C247_U487 : ADFULD1 port map( A => mult_21_C247_n1200, B => 
                           mult_21_C247_n1350, CI => mult_21_C247_n1320, CO => 
                           mult_21_C247_n646, S => mult_21_C247_n647);
   mult_21_C247_U486 : ADFULD1 port map( A => mult_21_C247_n1166, B => 
                           mult_21_C247_n1266, CI => mult_21_C247_n1220, CO => 
                           mult_21_C247_n644, S => mult_21_C247_n645);
   mult_21_C247_U485 : ADFULD1 port map( A => mult_21_C247_n1182, B => 
                           mult_21_C247_n1292, CI => mult_21_C247_n1242, CO => 
                           mult_21_C247_n642, S => mult_21_C247_n643);
   mult_21_C247_U484 : ADFULD1 port map( A => mult_21_C247_n649, B => 
                           mult_21_C247_n664, CI => mult_21_C247_n662, CO => 
                           mult_21_C247_n640, S => mult_21_C247_n641);
   mult_21_C247_U483 : ADFULD1 port map( A => mult_21_C247_n647, B => 
                           mult_21_C247_n660, CI => mult_21_C247_n643, CO => 
                           mult_21_C247_n638, S => mult_21_C247_n639);
   mult_21_C247_U482 : ADFULD1 port map( A => mult_21_C247_n658, B => 
                           mult_21_C247_n645, CI => mult_21_C247_n656, CO => 
                           mult_21_C247_n636, S => mult_21_C247_n637);
   mult_21_C247_U481 : ADFULD1 port map( A => mult_21_C247_n639, B => 
                           mult_21_C247_n641, CI => mult_21_C247_n654, CO => 
                           mult_21_C247_n634, S => mult_21_C247_n635);
   mult_21_C247_U480 : ADFULD1 port map( A => mult_21_C247_n652, B => 
                           mult_21_C247_n637, CI => mult_21_C247_n635, CO => 
                           mult_21_C247_n632, S => mult_21_C247_n633);
   mult_21_C247_U478 : ADFULD1 port map( A => mult_21_C247_n1151, B => 
                           mult_21_C247_n1199, CI => mult_21_C247_n1219, CO => 
                           mult_21_C247_n628, S => mult_21_C247_n629);
   mult_21_C247_U477 : ADFULD1 port map( A => mult_21_C247_n1291, B => 
                           mult_21_C247_n1181, CI => mult_21_C247_n1165, CO => 
                           mult_21_C247_n626, S => mult_21_C247_n627);
   mult_21_C247_U476 : ADFULD1 port map( A => mult_21_C247_n1241, B => 
                           mult_21_C247_n1265, CI => mult_21_C247_n648, CO => 
                           mult_21_C247_n624, S => mult_21_C247_n625);
   mult_21_C247_U475 : ADFULD1 port map( A => mult_21_C247_n646, B => 
                           mult_21_C247_n631, CI => mult_21_C247_n642, CO => 
                           mult_21_C247_n622, S => mult_21_C247_n623);
   mult_21_C247_U474 : ADFULD1 port map( A => mult_21_C247_n627, B => 
                           mult_21_C247_n644, CI => mult_21_C247_n629, CO => 
                           mult_21_C247_n620, S => mult_21_C247_n621);
   mult_21_C247_U473 : ADFULD1 port map( A => mult_21_C247_n640, B => 
                           mult_21_C247_n625, CI => mult_21_C247_n638, CO => 
                           mult_21_C247_n618, S => mult_21_C247_n619);
   mult_21_C247_U472 : ADFULD1 port map( A => mult_21_C247_n621, B => 
                           mult_21_C247_n623, CI => mult_21_C247_n636, CO => 
                           mult_21_C247_n616, S => mult_21_C247_n617);
   mult_21_C247_U471 : ADFULD1 port map( A => mult_21_C247_n634, B => 
                           mult_21_C247_n619, CI => mult_21_C247_n617, CO => 
                           mult_21_C247_n614, S => mult_21_C247_n615);
   mult_21_C247_U469 : ADFULD1 port map( A => mult_21_C247_n1164, B => 
                           mult_21_C247_n1348, CI => mult_21_C247_n1318, CO => 
                           mult_21_C247_n610, S => mult_21_C247_n611);
   mult_21_C247_U468 : ADFULD1 port map( A => mult_21_C247_n1290, B => 
                           mult_21_C247_n1198, CI => mult_21_C247_n1218, CO => 
                           mult_21_C247_n608, S => mult_21_C247_n609);
   mult_21_C247_U467 : ADFULD1 port map( A => mult_21_C247_n1150, B => 
                           mult_21_C247_n1264, CI => mult_21_C247_n1180, CO => 
                           mult_21_C247_n606, S => mult_21_C247_n607);
   mult_21_C247_U466 : ADFULD1 port map( A => mult_21_C247_n630, B => 
                           mult_21_C247_n1240, CI => mult_21_C247_n613, CO => 
                           mult_21_C247_n604, S => mult_21_C247_n605);
   mult_21_C247_U465 : ADFULD1 port map( A => mult_21_C247_n626, B => 
                           mult_21_C247_n628, CI => mult_21_C247_n624, CO => 
                           mult_21_C247_n602, S => mult_21_C247_n603);
   mult_21_C247_U464 : ADFULD1 port map( A => mult_21_C247_n609, B => 
                           mult_21_C247_n611, CI => mult_21_C247_n607, CO => 
                           mult_21_C247_n600, S => mult_21_C247_n601);
   mult_21_C247_U463 : ADFULD1 port map( A => mult_21_C247_n622, B => 
                           mult_21_C247_n605, CI => mult_21_C247_n620, CO => 
                           mult_21_C247_n598, S => mult_21_C247_n599);
   mult_21_C247_U462 : ADFULD1 port map( A => mult_21_C247_n601, B => 
                           mult_21_C247_n603, CI => mult_21_C247_n618, CO => 
                           mult_21_C247_n596, S => mult_21_C247_n597);
   mult_21_C247_U461 : ADFULD1 port map( A => mult_21_C247_n616, B => 
                           mult_21_C247_n599, CI => mult_21_C247_n597, CO => 
                           mult_21_C247_n594, S => mult_21_C247_n595);
   mult_21_C247_U459 : ADFULD1 port map( A => mult_21_C247_n1137, B => 
                           mult_21_C247_n1179, CI => mult_21_C247_n1217, CO => 
                           mult_21_C247_n590, S => mult_21_C247_n591);
   mult_21_C247_U458 : ADFULD1 port map( A => mult_21_C247_n1289, B => 
                           mult_21_C247_n1163, CI => mult_21_C247_n1149, CO => 
                           mult_21_C247_n588, S => mult_21_C247_n589);
   mult_21_C247_U457 : ADFULD1 port map( A => mult_21_C247_n1197, B => 
                           mult_21_C247_n1263, CI => mult_21_C247_n1239, CO => 
                           mult_21_C247_n586, S => mult_21_C247_n587);
   mult_21_C247_U456 : ADFULD1 port map( A => mult_21_C247_n593, B => 
                           mult_21_C247_n612, CI => mult_21_C247_n610, CO => 
                           mult_21_C247_n584, S => mult_21_C247_n585);
   mult_21_C247_U455 : ADFULD1 port map( A => mult_21_C247_n606, B => 
                           mult_21_C247_n608, CI => mult_21_C247_n587, CO => 
                           mult_21_C247_n582, S => mult_21_C247_n583);
   mult_21_C247_U454 : ADFULD1 port map( A => mult_21_C247_n591, B => 
                           mult_21_C247_n589, CI => mult_21_C247_n604, CO => 
                           mult_21_C247_n580, S => mult_21_C247_n581);
   mult_21_C247_U453 : ADFULD1 port map( A => mult_21_C247_n585, B => 
                           mult_21_C247_n602, CI => mult_21_C247_n600, CO => 
                           mult_21_C247_n578, S => mult_21_C247_n579);
   mult_21_C247_U452 : ADFULD1 port map( A => mult_21_C247_n581, B => 
                           mult_21_C247_n583, CI => mult_21_C247_n598, CO => 
                           mult_21_C247_n576, S => mult_21_C247_n577);
   mult_21_C247_U451 : ADFULD1 port map( A => mult_21_C247_n596, B => 
                           mult_21_C247_n579, CI => mult_21_C247_n577, CO => 
                           mult_21_C247_n574, S => mult_21_C247_n575);
   mult_21_C247_U449 : ADFULD1 port map( A => mult_21_C247_n1136, B => 
                           mult_21_C247_n1346, CI => mult_21_C247_n1316, CO => 
                           mult_21_C247_n570, S => mult_21_C247_n571);
   mult_21_C247_U448 : ADFULD1 port map( A => mult_21_C247_n1288, B => 
                           mult_21_C247_n1178, CI => mult_21_C247_n1216, CO => 
                           mult_21_C247_n568, S => mult_21_C247_n569);
   mult_21_C247_U447 : ADFULD1 port map( A => mult_21_C247_n1148, B => 
                           mult_21_C247_n1262, CI => mult_21_C247_n1162, CO => 
                           mult_21_C247_n566, S => mult_21_C247_n567);
   mult_21_C247_U446 : ADFULD1 port map( A => mult_21_C247_n1196, B => 
                           mult_21_C247_n1238, CI => mult_21_C247_n592, CO => 
                           mult_21_C247_n564, S => mult_21_C247_n565);
   mult_21_C247_U445 : ADFULD1 port map( A => mult_21_C247_n590, B => 
                           mult_21_C247_n573, CI => mult_21_C247_n588, CO => 
                           mult_21_C247_n562, S => mult_21_C247_n563);
   mult_21_C247_U444 : ADFULD1 port map( A => mult_21_C247_n571, B => 
                           mult_21_C247_n586, CI => mult_21_C247_n567, CO => 
                           mult_21_C247_n560, S => mult_21_C247_n561);
   mult_21_C247_U443 : ADFULD1 port map( A => mult_21_C247_n565, B => 
                           mult_21_C247_n569, CI => mult_21_C247_n584, CO => 
                           mult_21_C247_n558, S => mult_21_C247_n559);
   mult_21_C247_U442 : ADFULD1 port map( A => mult_21_C247_n563, B => 
                           mult_21_C247_n582, CI => mult_21_C247_n580, CO => 
                           mult_21_C247_n556, S => mult_21_C247_n557);
   mult_21_C247_U441 : ADFULD1 port map( A => mult_21_C247_n559, B => 
                           mult_21_C247_n561, CI => mult_21_C247_n578, CO => 
                           mult_21_C247_n554, S => mult_21_C247_n555);
   mult_21_C247_U440 : ADFULD1 port map( A => mult_21_C247_n576, B => 
                           mult_21_C247_n557, CI => mult_21_C247_n555, CO => 
                           mult_21_C247_n552, S => mult_21_C247_n553);
   mult_21_C247_U438 : ADFULD1 port map( A => mult_21_C247_n1125, B => 
                           mult_21_C247_n1177, CI => mult_21_C247_n1215, CO => 
                           mult_21_C247_n548, S => mult_21_C247_n549);
   mult_21_C247_U437 : ADFULD1 port map( A => mult_21_C247_n1287, B => 
                           mult_21_C247_n1161, CI => mult_21_C247_n1261, CO => 
                           mult_21_C247_n546, S => mult_21_C247_n547);
   mult_21_C247_U436 : ADFULD1 port map( A => mult_21_C247_n1135, B => 
                           mult_21_C247_n1237, CI => mult_21_C247_n1147, CO => 
                           mult_21_C247_n544, S => mult_21_C247_n545);
   mult_21_C247_U435 : ADFULD1 port map( A => mult_21_C247_n572, B => 
                           mult_21_C247_n1195, CI => mult_21_C247_n551, CO => 
                           mult_21_C247_n542, S => mult_21_C247_n543);
   mult_21_C247_U434 : ADFULD1 port map( A => mult_21_C247_n566, B => 
                           mult_21_C247_n570, CI => mult_21_C247_n568, CO => 
                           mult_21_C247_n540, S => mult_21_C247_n541);
   mult_21_C247_U433 : ADFULD1 port map( A => mult_21_C247_n549, B => 
                           mult_21_C247_n564, CI => mult_21_C247_n547, CO => 
                           mult_21_C247_n538, S => mult_21_C247_n539);
   mult_21_C247_U432 : ADFULD1 port map( A => mult_21_C247_n562, B => 
                           mult_21_C247_n545, CI => mult_21_C247_n543, CO => 
                           mult_21_C247_n536, S => mult_21_C247_n537);
   mult_21_C247_U431 : ADFULD1 port map( A => mult_21_C247_n541, B => 
                           mult_21_C247_n560, CI => mult_21_C247_n558, CO => 
                           mult_21_C247_n534, S => mult_21_C247_n535);
   mult_21_C247_U430 : ADFULD1 port map( A => mult_21_C247_n556, B => 
                           mult_21_C247_n539, CI => mult_21_C247_n537, CO => 
                           mult_21_C247_n532, S => mult_21_C247_n533);
   mult_21_C247_U429 : ADFULD1 port map( A => mult_21_C247_n554, B => 
                           mult_21_C247_n535, CI => mult_21_C247_n533, CO => 
                           mult_21_C247_n530, S => mult_21_C247_n531);
   mult_21_C247_U427 : ADFULD1 port map( A => mult_21_C247_n1146, B => 
                           mult_21_C247_n1344, CI => mult_21_C247_n1314, CO => 
                           mult_21_C247_n526, S => mult_21_C247_n527);
   mult_21_C247_U426 : ADFULD1 port map( A => mult_21_C247_n1124, B => 
                           mult_21_C247_n1176, CI => mult_21_C247_n1214, CO => 
                           mult_21_C247_n524, S => mult_21_C247_n525);
   mult_21_C247_U425 : ADFULD1 port map( A => mult_21_C247_n1134, B => 
                           mult_21_C247_n1286, CI => mult_21_C247_n1160, CO => 
                           mult_21_C247_n522, S => mult_21_C247_n523);
   mult_21_C247_U424 : ADFULD1 port map( A => mult_21_C247_n1194, B => 
                           mult_21_C247_n1260, CI => mult_21_C247_n1236, CO => 
                           mult_21_C247_n520, S => mult_21_C247_n521);
   mult_21_C247_U423 : ADFULD1 port map( A => mult_21_C247_n529, B => 
                           mult_21_C247_n550, CI => mult_21_C247_n548, CO => 
                           mult_21_C247_n518, S => mult_21_C247_n519);
   mult_21_C247_U422 : ADFULD1 port map( A => mult_21_C247_n544, B => 
                           mult_21_C247_n546, CI => mult_21_C247_n527, CO => 
                           mult_21_C247_n516, S => mult_21_C247_n517);
   mult_21_C247_U421 : ADFULD1 port map( A => mult_21_C247_n525, B => 
                           mult_21_C247_n521, CI => mult_21_C247_n523, CO => 
                           mult_21_C247_n514, S => mult_21_C247_n515);
   mult_21_C247_U420 : ADFULD1 port map( A => mult_21_C247_n540, B => 
                           mult_21_C247_n542, CI => mult_21_C247_n519, CO => 
                           mult_21_C247_n512, S => mult_21_C247_n513);
   mult_21_C247_U419 : ADFULD1 port map( A => mult_21_C247_n517, B => 
                           mult_21_C247_n538, CI => mult_21_C247_n515, CO => 
                           mult_21_C247_n510, S => mult_21_C247_n511);
   mult_21_C247_U418 : ADFULD1 port map( A => mult_21_C247_n513, B => 
                           mult_21_C247_n536, CI => mult_21_C247_n534, CO => 
                           mult_21_C247_n508, S => mult_21_C247_n509);
   mult_21_C247_U417 : ADFULD1 port map( A => mult_21_C247_n532, B => 
                           mult_21_C247_n511, CI => mult_21_C247_n509, CO => 
                           mult_21_C247_n506, S => mult_21_C247_n507);
   mult_21_C247_U415 : ADFULD1 port map( A => mult_21_C247_n1115, B => 
                           mult_21_C247_n1175, CI => mult_21_C247_n1213, CO => 
                           mult_21_C247_n502, S => mult_21_C247_n503);
   mult_21_C247_U414 : ADFULD1 port map( A => mult_21_C247_n1123, B => 
                           mult_21_C247_n1145, CI => mult_21_C247_n1133, CO => 
                           mult_21_C247_n500, S => mult_21_C247_n501);
   mult_21_C247_U413 : ADFULD1 port map( A => mult_21_C247_n1159, B => 
                           mult_21_C247_n1285, CI => mult_21_C247_n1193, CO => 
                           mult_21_C247_n498, S => mult_21_C247_n499);
   mult_21_C247_U412 : ADFULD1 port map( A => mult_21_C247_n1235, B => 
                           mult_21_C247_n1259, CI => mult_21_C247_n528, CO => 
                           mult_21_C247_n496, S => mult_21_C247_n497);
   mult_21_C247_U411 : ADFULD1 port map( A => mult_21_C247_n526, B => 
                           mult_21_C247_n505, CI => mult_21_C247_n520, CO => 
                           mult_21_C247_n494, S => mult_21_C247_n495);
   mult_21_C247_U410 : ADFULD1 port map( A => mult_21_C247_n522, B => 
                           mult_21_C247_n524, CI => mult_21_C247_n499, CO => 
                           mult_21_C247_n492, S => mult_21_C247_n493);
   mult_21_C247_U409 : ADFULD1 port map( A => mult_21_C247_n501, B => 
                           mult_21_C247_n503, CI => mult_21_C247_n497, CO => 
                           mult_21_C247_n490, S => mult_21_C247_n491);
   mult_21_C247_U408 : ADFULD1 port map( A => mult_21_C247_n516, B => 
                           mult_21_C247_n518, CI => mult_21_C247_n495, CO => 
                           mult_21_C247_n488, S => mult_21_C247_n489);
   mult_21_C247_U407 : ADFULD1 port map( A => mult_21_C247_n493, B => 
                           mult_21_C247_n514, CI => mult_21_C247_n491, CO => 
                           mult_21_C247_n486, S => mult_21_C247_n487);
   mult_21_C247_U406 : ADFULD1 port map( A => mult_21_C247_n510, B => 
                           mult_21_C247_n512, CI => mult_21_C247_n489, CO => 
                           mult_21_C247_n484, S => mult_21_C247_n485);
   mult_21_C247_U405 : ADFULD1 port map( A => mult_21_C247_n508, B => 
                           mult_21_C247_n487, CI => mult_21_C247_n485, CO => 
                           mult_21_C247_n482, S => mult_21_C247_n483);
   mult_21_C247_U403 : ADFULD1 port map( A => mult_21_C247_n1114, B => 
                           mult_21_C247_n1342, CI => mult_21_C247_n1312, CO => 
                           mult_21_C247_n478, S => mult_21_C247_n479);
   mult_21_C247_U402 : ADFULD1 port map( A => mult_21_C247_n1284, B => 
                           mult_21_C247_n1174, CI => mult_21_C247_n1212, CO => 
                           mult_21_C247_n476, S => mult_21_C247_n477);
   mult_21_C247_U401 : ADFULD1 port map( A => mult_21_C247_n1258, B => 
                           mult_21_C247_n1132, CI => mult_21_C247_n1122, CO => 
                           mult_21_C247_n474, S => mult_21_C247_n475);
   mult_21_C247_U400 : ADFULD1 port map( A => mult_21_C247_n1144, B => 
                           mult_21_C247_n1234, CI => mult_21_C247_n1158, CO => 
                           mult_21_C247_n472, S => mult_21_C247_n473);
   mult_21_C247_U399 : ADFULD1 port map( A => mult_21_C247_n504, B => 
                           mult_21_C247_n1192, CI => mult_21_C247_n481, CO => 
                           mult_21_C247_n470, S => mult_21_C247_n471);
   mult_21_C247_U398 : ADFULD1 port map( A => mult_21_C247_n498, B => 
                           mult_21_C247_n502, CI => mult_21_C247_n496, CO => 
                           mult_21_C247_n468, S => mult_21_C247_n469);
   mult_21_C247_U397 : ADFULD1 port map( A => mult_21_C247_n479, B => 
                           mult_21_C247_n500, CI => mult_21_C247_n473, CO => 
                           mult_21_C247_n466, S => mult_21_C247_n467);
   mult_21_C247_U396 : ADFULD1 port map( A => mult_21_C247_n475, B => 
                           mult_21_C247_n477, CI => mult_21_C247_n471, CO => 
                           mult_21_C247_n464, S => mult_21_C247_n465);
   mult_21_C247_U395 : ADFULD1 port map( A => mult_21_C247_n492, B => 
                           mult_21_C247_n494, CI => mult_21_C247_n490, CO => 
                           mult_21_C247_n462, S => mult_21_C247_n463);
   mult_21_C247_U394 : ADFULD1 port map( A => mult_21_C247_n467, B => 
                           mult_21_C247_n469, CI => mult_21_C247_n465, CO => 
                           mult_21_C247_n460, S => mult_21_C247_n461);
   mult_21_C247_U393 : ADFULD1 port map( A => mult_21_C247_n486, B => 
                           mult_21_C247_n488, CI => mult_21_C247_n463, CO => 
                           mult_21_C247_n458, S => mult_21_C247_n459);
   mult_21_C247_U392 : ADFULD1 port map( A => mult_21_C247_n484, B => 
                           mult_21_C247_n461, CI => mult_21_C247_n459, CO => 
                           mult_21_C247_n456, S => mult_21_C247_n457);
   mult_21_C247_U390 : ADFULD1 port map( A => mult_21_C247_n1107, B => 
                           mult_21_C247_n1157, CI => mult_21_C247_n1211, CO => 
                           mult_21_C247_n452, S => mult_21_C247_n453);
   mult_21_C247_U389 : ADFULD1 port map( A => mult_21_C247_n1283, B => 
                           mult_21_C247_n1143, CI => mult_21_C247_n1257, CO => 
                           mult_21_C247_n450, S => mult_21_C247_n451);
   mult_21_C247_U388 : ADFULD1 port map( A => mult_21_C247_n1113, B => 
                           mult_21_C247_n1233, CI => mult_21_C247_n1121, CO => 
                           mult_21_C247_n448, S => mult_21_C247_n449);
   mult_21_C247_U387 : ADFULD1 port map( A => mult_21_C247_n1131, B => 
                           mult_21_C247_n1191, CI => mult_21_C247_n1173, CO => 
                           mult_21_C247_n446, S => mult_21_C247_n447);
   mult_21_C247_U386 : ADFULD1 port map( A => mult_21_C247_n455, B => 
                           mult_21_C247_n480, CI => mult_21_C247_n478, CO => 
                           mult_21_C247_n444, S => mult_21_C247_n445);
   mult_21_C247_U385 : ADFULD1 port map( A => mult_21_C247_n474, B => 
                           mult_21_C247_n472, CI => mult_21_C247_n476, CO => 
                           mult_21_C247_n442, S => mult_21_C247_n443);
   mult_21_C247_U384 : ADFULD1 port map( A => mult_21_C247_n453, B => 
                           mult_21_C247_n447, CI => mult_21_C247_n470, CO => 
                           mult_21_C247_n440, S => mult_21_C247_n441);
   mult_21_C247_U383 : ADFULD1 port map( A => mult_21_C247_n449, B => 
                           mult_21_C247_n451, CI => mult_21_C247_n468, CO => 
                           mult_21_C247_n438, S => mult_21_C247_n439);
   mult_21_C247_U382 : ADFULD1 port map( A => mult_21_C247_n466, B => 
                           mult_21_C247_n445, CI => mult_21_C247_n443, CO => 
                           mult_21_C247_n436, S => mult_21_C247_n437);
   mult_21_C247_U381 : ADFULD1 port map( A => mult_21_C247_n441, B => 
                           mult_21_C247_n464, CI => mult_21_C247_n462, CO => 
                           mult_21_C247_n434, S => mult_21_C247_n435);
   mult_21_C247_U380 : ADFULD1 port map( A => mult_21_C247_n437, B => 
                           mult_21_C247_n439, CI => mult_21_C247_n460, CO => 
                           mult_21_C247_n432, S => mult_21_C247_n433);
   mult_21_C247_U379 : ADFULD1 port map( A => mult_21_C247_n458, B => 
                           mult_21_C247_n435, CI => mult_21_C247_n433, CO => 
                           mult_21_C247_n430, S => mult_21_C247_n431);
   mult_21_C247_U377 : ADFULD1 port map( A => mult_21_C247_n1106, B => 
                           mult_21_C247_n1340, CI => mult_21_C247_n1310, CO => 
                           mult_21_C247_n426, S => mult_21_C247_n427);
   mult_21_C247_U376 : ADFULD1 port map( A => mult_21_C247_n1282, B => 
                           mult_21_C247_n1156, CI => mult_21_C247_n1210, CO => 
                           mult_21_C247_n424, S => mult_21_C247_n425);
   mult_21_C247_U375 : ADFULD1 port map( A => mult_21_C247_n1112, B => 
                           mult_21_C247_n1130, CI => mult_21_C247_n1120, CO => 
                           mult_21_C247_n422, S => mult_21_C247_n423);
   mult_21_C247_U374 : ADFULD1 port map( A => mult_21_C247_n1142, B => 
                           mult_21_C247_n1256, CI => mult_21_C247_n1172, CO => 
                           mult_21_C247_n420, S => mult_21_C247_n421);
   mult_21_C247_U373 : ADFULD1 port map( A => mult_21_C247_n1232, B => 
                           mult_21_C247_n1190, CI => mult_21_C247_n454, CO => 
                           mult_21_C247_n418, S => mult_21_C247_n419);
   mult_21_C247_U372 : ADFULD1 port map( A => mult_21_C247_n452, B => 
                           mult_21_C247_n429, CI => mult_21_C247_n450, CO => 
                           mult_21_C247_n416, S => mult_21_C247_n417);
   mult_21_C247_U371 : ADFULD1 port map( A => mult_21_C247_n448, B => 
                           mult_21_C247_n446, CI => mult_21_C247_n427, CO => 
                           mult_21_C247_n414, S => mult_21_C247_n415);
   mult_21_C247_U370 : ADFULD1 port map( A => mult_21_C247_n421, B => 
                           mult_21_C247_n423, CI => mult_21_C247_n425, CO => 
                           mult_21_C247_n412, S => mult_21_C247_n413);
   mult_21_C247_U369 : ADFULD1 port map( A => mult_21_C247_n444, B => 
                           mult_21_C247_n419, CI => mult_21_C247_n442, CO => 
                           mult_21_C247_n410, S => mult_21_C247_n411);
   mult_21_C247_U368 : ADFULD1 port map( A => mult_21_C247_n440, B => 
                           mult_21_C247_n417, CI => mult_21_C247_n415, CO => 
                           mult_21_C247_n408, S => mult_21_C247_n409);
   mult_21_C247_U367 : ADFULD1 port map( A => mult_21_C247_n438, B => 
                           mult_21_C247_n413, CI => mult_21_C247_n411, CO => 
                           mult_21_C247_n406, S => mult_21_C247_n407);
   mult_21_C247_U366 : ADFULD1 port map( A => mult_21_C247_n409, B => 
                           mult_21_C247_n436, CI => mult_21_C247_n434, CO => 
                           mult_21_C247_n404, S => mult_21_C247_n405);
   mult_21_C247_U365 : ADFULD1 port map( A => mult_21_C247_n432, B => 
                           mult_21_C247_n407, CI => mult_21_C247_n405, CO => 
                           mult_21_C247_n402, S => mult_21_C247_n403);
   mult_21_C247_U363 : ADFULD1 port map( A => mult_21_C247_n1101, B => 
                           mult_21_C247_n1155, CI => mult_21_C247_n1209, CO => 
                           mult_21_C247_n398, S => mult_21_C247_n399);
   mult_21_C247_U362 : ADFULD1 port map( A => mult_21_C247_n1281, B => 
                           mult_21_C247_n1129, CI => mult_21_C247_n1105, CO => 
                           mult_21_C247_n396, S => mult_21_C247_n397);
   mult_21_C247_U361 : ADFULD1 port map( A => mult_21_C247_n1255, B => 
                           mult_21_C247_n1119, CI => mult_21_C247_n1111, CO => 
                           mult_21_C247_n394, S => mult_21_C247_n395);
   mult_21_C247_U360 : ADFULD1 port map( A => mult_21_C247_n1141, B => 
                           mult_21_C247_n1231, CI => mult_21_C247_n1171, CO => 
                           mult_21_C247_n392, S => mult_21_C247_n393);
   mult_21_C247_U359 : ADFULD1 port map( A => mult_21_C247_n428, B => 
                           mult_21_C247_n1189, CI => mult_21_C247_n401, CO => 
                           mult_21_C247_n390, S => mult_21_C247_n391);
   mult_21_C247_U358 : ADFULD1 port map( A => mult_21_C247_n424, B => 
                           mult_21_C247_n426, CI => mult_21_C247_n420, CO => 
                           mult_21_C247_n388, S => mult_21_C247_n389);
   mult_21_C247_U357 : ADFULD1 port map( A => mult_21_C247_n418, B => 
                           mult_21_C247_n422, CI => mult_21_C247_n393, CO => 
                           mult_21_C247_n386, S => mult_21_C247_n387);
   mult_21_C247_U356 : ADFULD1 port map( A => mult_21_C247_n395, B => 
                           mult_21_C247_n397, CI => mult_21_C247_n399, CO => 
                           mult_21_C247_n384, S => mult_21_C247_n385);
   mult_21_C247_U355 : ADFULD1 port map( A => mult_21_C247_n391, B => 
                           mult_21_C247_n416, CI => mult_21_C247_n414, CO => 
                           mult_21_C247_n382, S => mult_21_C247_n383);
   mult_21_C247_U354 : ADFULD1 port map( A => mult_21_C247_n412, B => 
                           mult_21_C247_n389, CI => mult_21_C247_n387, CO => 
                           mult_21_C247_n380, S => mult_21_C247_n381);
   mult_21_C247_U353 : ADFULD1 port map( A => mult_21_C247_n410, B => 
                           mult_21_C247_n385, CI => mult_21_C247_n383, CO => 
                           mult_21_C247_n378, S => mult_21_C247_n379);
   mult_21_C247_U352 : ADFULD1 port map( A => mult_21_C247_n381, B => 
                           mult_21_C247_n408, CI => mult_21_C247_n406, CO => 
                           mult_21_C247_n376, S => mult_21_C247_n377);
   mult_21_C247_U351 : ADFULD1 port map( A => mult_21_C247_n404, B => 
                           mult_21_C247_n379, CI => mult_21_C247_n377, CO => 
                           mult_21_C247_n374, S => mult_21_C247_n375);
   mult_21_C247_U349 : ADFULD1 port map( A => mult_21_C247_n1100, B => 
                           mult_21_C247_n1338, CI => mult_21_C247_n1308, CO => 
                           mult_21_C247_n370, S => mult_21_C247_n371);
   mult_21_C247_U348 : ADFULD1 port map( A => mult_21_C247_n1280, B => 
                           mult_21_C247_n1154, CI => mult_21_C247_n1208, CO => 
                           mult_21_C247_n368, S => mult_21_C247_n369);
   mult_21_C247_U347 : ADFULD1 port map( A => mult_21_C247_n1254, B => 
                           mult_21_C247_n1128, CI => mult_21_C247_n1230, CO => 
                           mult_21_C247_n366, S => mult_21_C247_n367);
   mult_21_C247_U346 : ADFULD1 port map( A => mult_21_C247_n1104, B => 
                           mult_21_C247_n1188, CI => mult_21_C247_n1110, CO => 
                           mult_21_C247_n364, S => mult_21_C247_n365);
   mult_21_C247_U345 : ADFULD1 port map( A => mult_21_C247_n1170, B => 
                           mult_21_C247_n1118, CI => mult_21_C247_n1140, CO => 
                           mult_21_C247_n362, S => mult_21_C247_n363);
   mult_21_C247_U344 : ADFULD1 port map( A => mult_21_C247_n373, B => 
                           mult_21_C247_n400, CI => mult_21_C247_n392, CO => 
                           mult_21_C247_n360, S => mult_21_C247_n361);
   mult_21_C247_U343 : ADFULD1 port map( A => mult_21_C247_n398, B => 
                           mult_21_C247_n394, CI => mult_21_C247_n396, CO => 
                           mult_21_C247_n358, S => mult_21_C247_n359);
   mult_21_C247_U342 : ADFULD1 port map( A => mult_21_C247_n369, B => 
                           mult_21_C247_n371, CI => mult_21_C247_n367, CO => 
                           mult_21_C247_n356, S => mult_21_C247_n357);
   mult_21_C247_U341 : ADFULD1 port map( A => mult_21_C247_n365, B => 
                           mult_21_C247_n363, CI => mult_21_C247_n390, CO => 
                           mult_21_C247_n354, S => mult_21_C247_n355);
   mult_21_C247_U340 : ADFULD1 port map( A => mult_21_C247_n361, B => 
                           mult_21_C247_n388, CI => mult_21_C247_n386, CO => 
                           mult_21_C247_n352, S => mult_21_C247_n353);
   mult_21_C247_U339 : ADFULD1 port map( A => mult_21_C247_n359, B => 
                           mult_21_C247_n384, CI => mult_21_C247_n357, CO => 
                           mult_21_C247_n350, S => mult_21_C247_n351);
   mult_21_C247_U338 : ADFULD1 port map( A => mult_21_C247_n382, B => 
                           mult_21_C247_n355, CI => mult_21_C247_n380, CO => 
                           mult_21_C247_n348, S => mult_21_C247_n349);
   mult_21_C247_U337 : ADFULD1 port map( A => mult_21_C247_n351, B => 
                           mult_21_C247_n353, CI => mult_21_C247_n378, CO => 
                           mult_21_C247_n346, S => mult_21_C247_n347);
   mult_21_C247_U336 : ADFULD1 port map( A => mult_21_C247_n376, B => 
                           mult_21_C247_n349, CI => mult_21_C247_n347, CO => 
                           mult_21_C247_n344, S => mult_21_C247_n345);
   mult_21_C247_U334 : EXOR3D1 port map( A1 => mult_21_C247_n1097, A2 => 
                           mult_21_C247_n1279, A3 => mult_21_C247_n1207, Z => 
                           mult_21_C247_n342);
   mult_21_C247_U333 : EXOR3D1 port map( A1 => mult_21_C247_n1253, A2 => 
                           mult_21_C247_n1127, A3 => mult_21_C247_n1099, Z => 
                           mult_21_C247_n341);
   mult_21_C247_U332 : EXOR3D1 port map( A1 => mult_21_C247_n1103, A2 => 
                           mult_21_C247_n1117, A3 => mult_21_C247_n1109, Z => 
                           mult_21_C247_n340);
   mult_21_C247_U331 : EXOR3D1 port map( A1 => mult_21_C247_n1139, A2 => 
                           mult_21_C247_n1229, A3 => mult_21_C247_n1153, Z => 
                           mult_21_C247_n339);
   mult_21_C247_U330 : EXOR3D1 port map( A1 => mult_21_C247_n1187, A2 => 
                           mult_21_C247_n1169, A3 => mult_21_C247_n372, Z => 
                           mult_21_C247_n338);
   mult_21_C247_U329 : EXOR3D1 port map( A1 => mult_21_C247_n368, A2 => 
                           mult_21_C247_n370, A3 => mult_21_C247_n364, Z => 
                           mult_21_C247_n337);
   mult_21_C247_U328 : EXOR3D1 port map( A1 => mult_21_C247_n366, A2 => 
                           mult_21_C247_n343, A3 => mult_21_C247_n362, Z => 
                           mult_21_C247_n336);
   mult_21_C247_U327 : EXOR3D1 port map( A1 => mult_21_C247_n342, A2 => 
                           mult_21_C247_n338, A3 => mult_21_C247_n341, Z => 
                           mult_21_C247_n335);
   mult_21_C247_U326 : EXOR3D1 port map( A1 => mult_21_C247_n339, A2 => 
                           mult_21_C247_n340, A3 => mult_21_C247_n360, Z => 
                           mult_21_C247_n334);
   mult_21_C247_U325 : EXOR3D1 port map( A1 => mult_21_C247_n337, A2 => 
                           mult_21_C247_n358, A3 => mult_21_C247_n336, Z => 
                           mult_21_C247_n333);
   mult_21_C247_U324 : EXOR3D1 port map( A1 => mult_21_C247_n354, A2 => 
                           mult_21_C247_n356, A3 => mult_21_C247_n335, Z => 
                           mult_21_C247_n332);
   mult_21_C247_U323 : EXOR3D1 port map( A1 => mult_21_C247_n352, A2 => 
                           mult_21_C247_n334, A3 => mult_21_C247_n333, Z => 
                           mult_21_C247_n331);
   mult_21_C247_U322 : EXOR3D1 port map( A1 => mult_21_C247_n332, A2 => 
                           mult_21_C247_n350, A3 => mult_21_C247_n348, Z => 
                           mult_21_C247_n330);
   mult_21_C247_U321 : EXOR3D1 port map( A1 => mult_21_C247_n346, A2 => 
                           mult_21_C247_n331, A3 => mult_21_C247_n330, Z => 
                           mult_21_C247_n329);
   mult_21_C247_U313 : EXOR2D1 port map( A1 => mult_21_C247_n303, A2 => 
                           mult_21_C247_n305, Z => N3330);
   mult_21_C247_U305 : EXNOR2D1 port map( A1 => mult_21_C247_n176, A2 => 
                           mult_21_C247_n302, Z => N3331);
   mult_21_C247_U300 : OAI21D1 port map( A1 => mult_21_C247_n297, A2 => 
                           mult_21_C247_n295, B => mult_21_C247_n296, Z => 
                           mult_21_C247_n294);
   mult_21_C247_U299 : EXOR2D1 port map( A1 => mult_21_C247_n297, A2 => 
                           mult_21_C247_n175, Z => N3332);
   mult_21_C247_U291 : EXNOR2D1 port map( A1 => mult_21_C247_n174, A2 => 
                           mult_21_C247_n294, Z => N3333);
   mult_21_C247_U286 : OAI21D1 port map( A1 => mult_21_C247_n289, A2 => 
                           mult_21_C247_n287, B => mult_21_C247_n288, Z => 
                           mult_21_C247_n286);
   mult_21_C247_U284 : EXOR2D1 port map( A1 => mult_21_C247_n173, A2 => 
                           mult_21_C247_n289, Z => N3334);
   mult_21_C247_U279 : OAI21D1 port map( A1 => mult_21_C247_n285, A2 => 
                           mult_21_C247_n283, B => mult_21_C247_n284, Z => 
                           mult_21_C247_n282);
   mult_21_C247_U278 : EXOR2D1 port map( A1 => mult_21_C247_n172, A2 => 
                           mult_21_C247_n285, Z => N3335);
   mult_21_C247_U273 : OAI21D1 port map( A1 => mult_21_C247_n280, A2 => 
                           mult_21_C247_n284, B => mult_21_C247_n281, Z => 
                           mult_21_C247_n279);
   mult_21_C247_U271 : AOI21D1 port map( A1 => mult_21_C247_n278, A2 => 
                           mult_21_C247_n286, B => mult_21_C247_n279, Z => 
                           mult_21_C247_n277);
   mult_21_C247_U269 : EXNOR2D1 port map( A1 => mult_21_C247_n282, A2 => 
                           mult_21_C247_n171, Z => N3336);
   mult_21_C247_U262 : AOI21D1 port map( A1 => mult_21_C247_n276, A2 => 
                           mult_21_C247_n1527, B => mult_21_C247_n273, Z => 
                           mult_21_C247_n271);
   mult_21_C247_U261 : EXNOR2D1 port map( A1 => mult_21_C247_n276, A2 => 
                           mult_21_C247_n170, Z => N3337);
   mult_21_C247_U254 : AOI21D1 port map( A1 => mult_21_C247_n1524, A2 => 
                           mult_21_C247_n273, B => mult_21_C247_n268, Z => 
                           mult_21_C247_n266);
   mult_21_C247_U252 : OAI21D1 port map( A1 => mult_21_C247_n265, A2 => 
                           mult_21_C247_n277, B => mult_21_C247_n266, Z => 
                           mult_21_C247_n264);
   mult_21_C247_U250 : EXOR2D1 port map( A1 => mult_21_C247_n271, A2 => 
                           mult_21_C247_n169, Z => N3338);
   mult_21_C247_U245 : OAI21D1 port map( A1 => mult_21_C247_n263, A2 => 
                           mult_21_C247_n261, B => mult_21_C247_n262, Z => 
                           mult_21_C247_n260);
   mult_21_C247_U244 : EXOR2D1 port map( A1 => mult_21_C247_n263, A2 => 
                           mult_21_C247_n168, Z => N3339);
   mult_21_C247_U239 : OAI21D1 port map( A1 => mult_21_C247_n258, A2 => 
                           mult_21_C247_n262, B => mult_21_C247_n259, Z => 
                           mult_21_C247_n257);
   mult_21_C247_U237 : AOI21D1 port map( A1 => mult_21_C247_n256, A2 => 
                           mult_21_C247_n264, B => mult_21_C247_n257, Z => 
                           mult_21_C247_n255);
   mult_21_C247_U235 : EXNOR2D1 port map( A1 => mult_21_C247_n260, A2 => 
                           mult_21_C247_n167, Z => N3340);
   mult_21_C247_U228 : AOI21D1 port map( A1 => mult_21_C247_n254, A2 => 
                           mult_21_C247_n1529, B => mult_21_C247_n251, Z => 
                           mult_21_C247_n249);
   mult_21_C247_U227 : EXNOR2D1 port map( A1 => mult_21_C247_n254, A2 => 
                           mult_21_C247_n166, Z => N3341);
   mult_21_C247_U220 : AOI21D1 port map( A1 => mult_21_C247_n1530, A2 => 
                           mult_21_C247_n251, B => mult_21_C247_n246, Z => 
                           mult_21_C247_n244);
   mult_21_C247_U218 : OAI21D1 port map( A1 => mult_21_C247_n255, A2 => 
                           mult_21_C247_n243, B => mult_21_C247_n244, Z => 
                           mult_21_C247_n242);
   mult_21_C247_U216 : EXOR2D1 port map( A1 => mult_21_C247_n249, A2 => 
                           mult_21_C247_n165, Z => N3342);
   mult_21_C247_U211 : OAI21D1 port map( A1 => mult_21_C247_n241, A2 => 
                           mult_21_C247_n239, B => mult_21_C247_n240, Z => 
                           mult_21_C247_n238);
   mult_21_C247_U210 : EXOR2D1 port map( A1 => mult_21_C247_n241, A2 => 
                           mult_21_C247_n164, Z => N3343);
   mult_21_C247_U205 : OAI21D1 port map( A1 => mult_21_C247_n236, A2 => 
                           mult_21_C247_n240, B => mult_21_C247_n237, Z => 
                           mult_21_C247_n235);
   mult_21_C247_U203 : AOI21D1 port map( A1 => mult_21_C247_n242, A2 => 
                           mult_21_C247_n234, B => mult_21_C247_n235, Z => 
                           mult_21_C247_n233);
   mult_21_C247_U201 : EXNOR2D1 port map( A1 => mult_21_C247_n238, A2 => 
                           mult_21_C247_n163, Z => N3344);
   mult_21_C247_U194 : AOI21D1 port map( A1 => mult_21_C247_n232, A2 => 
                           mult_21_C247_n313, B => mult_21_C247_n229, Z => 
                           mult_21_C247_n227);
   mult_21_C247_U193 : EXNOR2D1 port map( A1 => mult_21_C247_n232, A2 => 
                           mult_21_C247_n162, Z => N3345);
   mult_21_C247_U188 : OAI21D1 port map( A1 => mult_21_C247_n225, A2 => 
                           mult_21_C247_n231, B => mult_21_C247_n226, Z => 
                           mult_21_C247_n224);
   mult_21_C247_U186 : AOI21D1 port map( A1 => mult_21_C247_n232, A2 => 
                           mult_21_C247_n223, B => mult_21_C247_n224, Z => 
                           mult_21_C247_n222);
   mult_21_C247_U185 : EXOR2D1 port map( A1 => mult_21_C247_n227, A2 => 
                           mult_21_C247_n161, Z => N3346);
   mult_21_C247_U178 : AOI21D1 port map( A1 => mult_21_C247_n224, A2 => 
                           mult_21_C247_n1528, B => mult_21_C247_n219, Z => 
                           mult_21_C247_n217);
   mult_21_C247_U176 : OAI21D1 port map( A1 => mult_21_C247_n233, A2 => 
                           mult_21_C247_n216, B => mult_21_C247_n217, Z => 
                           mult_21_C247_n215);
   mult_21_C247_U174 : EXOR2D1 port map( A1 => mult_21_C247_n222, A2 => 
                           mult_21_C247_n160, Z => N3347);
   mult_21_C247_U165 : OAI21D1 port map( A1 => mult_21_C247_n214, A2 => 
                           mult_21_C247_n208, B => mult_21_C247_n209, Z => 
                           mult_21_C247_n207);
   mult_21_C247_U164 : EXOR2D1 port map( A1 => mult_21_C247_n214, A2 => 
                           mult_21_C247_n159, Z => N3348);
   mult_21_C247_U157 : AOI21D1 port map( A1 => mult_21_C247_n1525, A2 => 
                           mult_21_C247_n211, B => mult_21_C247_n204, Z => 
                           mult_21_C247_n202);
   mult_21_C247_U155 : OAI21D1 port map( A1 => mult_21_C247_n214, A2 => 
                           mult_21_C247_n201, B => mult_21_C247_n202, Z => 
                           mult_21_C247_n200);
   mult_21_C247_U154 : EXNOR2D1 port map( A1 => mult_21_C247_n207, A2 => 
                           mult_21_C247_n158, Z => N3349);
   mult_21_C247_U147 : AOI21D1 port map( A1 => mult_21_C247_n200, A2 => 
                           mult_21_C247_n1526, B => mult_21_C247_n197, Z => 
                           mult_21_C247_n195);
   mult_21_C247_U146 : EXNOR2D1 port map( A1 => mult_21_C247_n200, A2 => 
                           mult_21_C247_n157, Z => N3350);
   mult_21_C247_U137 : OAI21D1 port map( A1 => mult_21_C247_n202, A2 => 
                           mult_21_C247_n189, B => mult_21_C247_n190, Z => 
                           mult_21_C247_n188);
   mult_21_C247_U134 : EXOR2D1 port map( A1 => mult_21_C247_n195, A2 => 
                           mult_21_C247_n156, Z => N3351);
   mult_21_C247_U132 : ADFULD1 port map( A => mult_21_C247_n531, B => 
                           mult_21_C247_n552, CI => mult_21_C247_n1521, CO => 
                           mult_21_C247_n185, S => N3352);
   mult_21_C247_U131 : ADFULD1 port map( A => mult_21_C247_n507, B => 
                           mult_21_C247_n530, CI => mult_21_C247_n185, CO => 
                           mult_21_C247_n184, S => N3353);
   mult_21_C247_U130 : ADFULD1 port map( A => mult_21_C247_n483, B => 
                           mult_21_C247_n506, CI => mult_21_C247_n184, CO => 
                           mult_21_C247_n183, S => N3354);
   mult_21_C247_U129 : ADFULD1 port map( A => mult_21_C247_n457, B => 
                           mult_21_C247_n482, CI => mult_21_C247_n183, CO => 
                           mult_21_C247_n182, S => N3355);
   mult_21_C247_U128 : ADFULD1 port map( A => mult_21_C247_n431, B => 
                           mult_21_C247_n456, CI => mult_21_C247_n182, CO => 
                           mult_21_C247_n181, S => N3356);
   mult_21_C247_U127 : ADFULD1 port map( A => mult_21_C247_n403, B => 
                           mult_21_C247_n430, CI => mult_21_C247_n181, CO => 
                           mult_21_C247_n180, S => N3357);
   mult_21_C247_U126 : ADFULD1 port map( A => mult_21_C247_n375, B => 
                           mult_21_C247_n402, CI => mult_21_C247_n180, CO => 
                           mult_21_C247_n179, S => N3358);
   mult_21_C247_U125 : ADFULD1 port map( A => mult_21_C247_n345, B => 
                           mult_21_C247_n374, CI => mult_21_C247_n179, CO => 
                           mult_21_C247_n178, S => N3359);
   mult_21_C249_U1403 : INVD1 port map( A => N3072, Z => mult_21_C249_n1066);
   mult_21_C249_U1402 : AO21D1 port map( A1 => N3070, A2 => N3071, B => 
                           mult_21_C249_n1066, Z => mult_21_C249_n105);
   mult_21_C249_U1401 : INVD1 port map( A => N3070, Z => mult_21_C249_n1067);
   mult_21_C249_U1400 : AO21D1 port map( A1 => N3068, A2 => N3069, B => 
                           mult_21_C249_n1067, Z => mult_21_C249_n101);
   mult_21_C249_U1399 : INVD1 port map( A => N3068, Z => mult_21_C249_n1068);
   mult_21_C249_U1398 : AO21D1 port map( A1 => N3066, A2 => N3067, B => 
                           mult_21_C249_n1068, Z => mult_21_C249_n96);
   mult_21_C249_U1397 : ADHALFDL port map( A => mult_21_C249_n1309, B => 
                           mult_21_C249_n1339, CO => mult_21_C249_n400, S => 
                           mult_21_C249_n401);
   mult_21_C249_U1396 : AO21D1 port map( A1 => N3064, A2 => N3065, B => 
                           mult_21_C249_n1069, Z => mult_21_C249_n91);
   mult_21_C249_U1395 : INVD1 port map( A => N3066, Z => mult_21_C249_n1069);
   mult_21_C249_U1394 : ADHALFDL port map( A => mult_21_C249_n1311, B => 
                           mult_21_C249_n1341, CO => mult_21_C249_n454, S => 
                           mult_21_C249_n455);
   mult_21_C249_U1393 : OAI21D1 port map( A1 => N3064, A2 => N3065, B => 
                           mult_21_C249_n1069, Z => mult_21_C249_n89);
   mult_21_C249_U1392 : ADHALFDL port map( A => mult_21_C249_n1313, B => 
                           mult_21_C249_n1343, CO => mult_21_C249_n504, S => 
                           mult_21_C249_n505);
   mult_21_C249_U1391 : AO21D1 port map( A1 => N3062, A2 => N3063, B => 
                           mult_21_C249_n1070, Z => mult_21_C249_n86);
   mult_21_C249_U1390 : INVD1 port map( A => N3064, Z => mult_21_C249_n1070);
   mult_21_C249_U1389 : OAI21D1 port map( A1 => N3062, A2 => N3063, B => 
                           mult_21_C249_n1070, Z => mult_21_C249_n84);
   mult_21_C249_U1388 : AO21D1 port map( A1 => N3060, A2 => N3061, B => 
                           mult_21_C249_n1071, Z => mult_21_C249_n81);
   mult_21_C249_U1387 : INVD1 port map( A => N3062, Z => mult_21_C249_n1071);
   mult_21_C249_U1386 : OAI21D1 port map( A1 => N3060, A2 => N3061, B => 
                           mult_21_C249_n1071, Z => mult_21_C249_n79);
   mult_21_C249_U1385 : EXNOR2D1 port map( A1 => N3062, A2 => N3063, Z => 
                           mult_21_C249_n88);
   mult_21_C249_U1384 : AO21D1 port map( A1 => N3058, A2 => N3059, B => 
                           mult_21_C249_n1072, Z => mult_21_C249_n76);
   mult_21_C249_U1383 : OAI21D1 port map( A1 => N3050, A2 => N3051, B => 
                           mult_21_C249_n1076, Z => mult_21_C249_n42);
   mult_21_C249_U1382 : INVD1 port map( A => N3060, Z => mult_21_C249_n1072);
   mult_21_C249_U1381 : OAI21D1 port map( A1 => N3058, A2 => N3059, B => 
                           mult_21_C249_n1072, Z => mult_21_C249_n73);
   mult_21_C249_U1380 : INVD1 port map( A => N3052, Z => mult_21_C249_n1076);
   mult_21_C249_U1379 : AO21D1 port map( A1 => N3050, A2 => N3051, B => 
                           mult_21_C249_n1076, Z => mult_21_C249_n45);
   mult_21_C249_U1378 : OAI21D1 port map( A1 => N3056, A2 => N3057, B => 
                           mult_21_C249_n1073, Z => mult_21_C249_n66);
   mult_21_C249_U1377 : INVD1 port map( A => N3058, Z => mult_21_C249_n1073);
   mult_21_C249_U1376 : OAI21D1 port map( A1 => N3054, A2 => N3055, B => 
                           mult_21_C249_n1074, Z => mult_21_C249_n58);
   mult_21_C249_U1375 : INVD1 port map( A => N3056, Z => mult_21_C249_n1074);
   mult_21_C249_U1374 : AO21D1 port map( A1 => N3056, A2 => N3057, B => 
                           mult_21_C249_n1073, Z => mult_21_C249_n69);
   mult_21_C249_U1373 : AO21D1 port map( A1 => N3054, A2 => N3055, B => 
                           mult_21_C249_n1074, Z => mult_21_C249_n61);
   mult_21_C249_U1372 : OAI21D1 port map( A1 => N3052, A2 => N3053, B => 
                           mult_21_C249_n1075, Z => mult_21_C249_n50);
   mult_21_C249_U1371 : AO21D1 port map( A1 => N3048, A2 => N3049, B => 
                           mult_21_C249_n1077, Z => mult_21_C249_n38);
   mult_21_C249_U1370 : AO21D1 port map( A1 => N3044, A2 => N3045, B => 
                           mult_21_C249_n1079, Z => mult_21_C249_n22);
   mult_21_C249_U1369 : ADHALFDL port map( A => mult_21_C249_n1315, B => 
                           mult_21_C249_n1345, CO => mult_21_C249_n550, S => 
                           mult_21_C249_n551);
   mult_21_C249_U1368 : INVD1 port map( A => N3054, Z => mult_21_C249_n1075);
   mult_21_C249_U1367 : AO21D1 port map( A1 => N3052, A2 => N3053, B => 
                           mult_21_C249_n1075, Z => mult_21_C249_n53);
   mult_21_C249_U1366 : INVD1 port map( A => N3041, Z => mult_21_C249_n8);
   mult_21_C249_U1365 : EXNOR2D1 port map( A1 => N3060, A2 => N3061, Z => 
                           mult_21_C249_n83);
   mult_21_C249_U1364 : AO21D1 port map( A1 => N3046, A2 => N3047, B => 
                           mult_21_C249_n1078, Z => mult_21_C249_n30);
   mult_21_C249_U1363 : AO21D1 port map( A1 => N3042, A2 => N3043, B => 
                           mult_21_C249_n1080, Z => mult_21_C249_n14);
   mult_21_C249_U1362 : EXNOR2D1 port map( A1 => N3058, A2 => N3059, Z => 
                           mult_21_C249_n78);
   mult_21_C249_U1361 : EXNOR2D1 port map( A1 => N3050, A2 => N3051, Z => 
                           mult_21_C249_n48);
   mult_21_C249_U1360 : INVD1 port map( A => N3046, Z => mult_21_C249_n1079);
   mult_21_C249_U1359 : INVD1 port map( A => n288, Z => mult_21_C249_n1557);
   mult_21_C249_U1358 : EXNOR2D1 port map( A1 => N3056, A2 => N3057, Z => 
                           mult_21_C249_n71);
   mult_21_C249_U1357 : EXNOR2D1 port map( A1 => N3054, A2 => N3055, Z => 
                           mult_21_C249_n63);
   mult_21_C249_U1356 : INVD1 port map( A => n287, Z => mult_21_C249_n1550);
   mult_21_C249_U1355 : INVD1 port map( A => n286, Z => mult_21_C249_n1552);
   mult_21_C249_U1354 : INVD1 port map( A => N3050, Z => mult_21_C249_n1077);
   mult_21_C249_U1353 : INVD1 port map( A => N3042, Z => mult_21_C249_n6);
   mult_21_C249_U1352 : NAN2D1 port map( A1 => N3041, A2 => mult_21_C249_n6, Z 
                           => mult_21_C249_n3);
   mult_21_C249_U1351 : INVD1 port map( A => n283, Z => mult_21_C249_n1555);
   mult_21_C249_U1350 : INVD1 port map( A => n282, Z => mult_21_C249_n1548);
   mult_21_C249_U1349 : INVD1 port map( A => N3048, Z => mult_21_C249_n1078);
   mult_21_C249_U1348 : INVD1 port map( A => n281, Z => mult_21_C249_n1542);
   mult_21_C249_U1347 : EXNOR2D1 port map( A1 => N3052, A2 => N3053, Z => 
                           mult_21_C249_n56);
   mult_21_C249_U1346 : INVD1 port map( A => N3044, Z => mult_21_C249_n1080);
   mult_21_C249_U1345 : INVD1 port map( A => n279, Z => mult_21_C249_n1544);
   mult_21_C249_U1344 : INVD1 port map( A => n278, Z => mult_21_C249_n1546);
   mult_21_C249_U1343 : OA21D1 port map( A1 => N3046, A2 => N3047, B => 
                           mult_21_C249_n1078, Z => mult_21_C249_n1537);
   mult_21_C249_U1342 : ADHALFDL port map( A => mult_21_C249_n1325, B => 
                           mult_21_C249_n1355, CO => mult_21_C249_n720, S => 
                           mult_21_C249_n721);
   mult_21_C249_U1341 : ADHALFDL port map( A => mult_21_C249_n1321, B => 
                           mult_21_C249_n1351, CO => mult_21_C249_n664, S => 
                           mult_21_C249_n665);
   mult_21_C249_U1340 : ADHALFDL port map( A => mult_21_C249_n1319, B => 
                           mult_21_C249_n1349, CO => mult_21_C249_n630, S => 
                           mult_21_C249_n631);
   mult_21_C249_U1339 : ADHALFDL port map( A => mult_21_C249_n1327, B => 
                           mult_21_C249_n1357, CO => mult_21_C249_n742, S => 
                           mult_21_C249_n743);
   mult_21_C249_U1338 : ADHALFDL port map( A => mult_21_C249_n1317, B => 
                           mult_21_C249_n1347, CO => mult_21_C249_n592, S => 
                           mult_21_C249_n593);
   mult_21_C249_U1337 : EXOR2D1 port map( A1 => N3044, A2 => N3045, Z => 
                           mult_21_C249_n1536);
   mult_21_C249_U1336 : ADHALFDL port map( A => mult_21_C249_n1323, B => 
                           mult_21_C249_n1353, CO => mult_21_C249_n694, S => 
                           mult_21_C249_n695);
   mult_21_C249_U1335 : EXOR2D1 port map( A1 => N3042, A2 => N3043, Z => 
                           mult_21_C249_n1535);
   mult_21_C249_U1334 : ADHALFDL port map( A => mult_21_C249_n1098, B => 
                           mult_21_C249_n1081, CO => mult_21_C249_n372, S => 
                           mult_21_C249_n373);
   mult_21_C249_U1333 : EXOR2D1 port map( A1 => mult_21_C249_n1307, A2 => 
                           mult_21_C249_n1337, Z => mult_21_C249_n343);
   mult_21_C249_U1332 : ADHALFDL port map( A => mult_21_C249_n1102, B => 
                           mult_21_C249_n1082, CO => mult_21_C249_n428, S => 
                           mult_21_C249_n429);
   mult_21_C249_U1331 : ADHALFDL port map( A => mult_21_C249_n1108, B => 
                           mult_21_C249_n1083, CO => mult_21_C249_n480, S => 
                           mult_21_C249_n481);
   mult_21_C249_U1330 : ADHALFDL port map( A => mult_21_C249_n1116, B => 
                           mult_21_C249_n1084, CO => mult_21_C249_n528, S => 
                           mult_21_C249_n529);
   mult_21_C249_U1329 : ADHALFDL port map( A => mult_21_C249_n1126, B => 
                           mult_21_C249_n1085, CO => mult_21_C249_n572, S => 
                           mult_21_C249_n573);
   mult_21_C249_U1328 : INVD1 port map( A => mult_21_C249_n1367, Z => 
                           mult_21_C249_n303);
   mult_21_C249_U1327 : ADHALFDL port map( A => mult_21_C249_n1138, B => 
                           mult_21_C249_n1086, CO => mult_21_C249_n612, S => 
                           mult_21_C249_n613);
   mult_21_C249_U1326 : ADHALFDL port map( A => mult_21_C249_n1186, B => 
                           mult_21_C249_n1089, CO => mult_21_C249_n708, S => 
                           mult_21_C249_n709);
   mult_21_C249_U1325 : ADHALFDL port map( A => mult_21_C249_n1228, B => 
                           mult_21_C249_n1091, CO => mult_21_C249_n752, S => 
                           mult_21_C249_n753);
   mult_21_C249_U1324 : ADHALFDL port map( A => mult_21_C249_n1152, B => 
                           mult_21_C249_n1087, CO => mult_21_C249_n648, S => 
                           mult_21_C249_n649);
   mult_21_C249_U1323 : ADHALFDL port map( A => mult_21_C249_n1168, B => 
                           mult_21_C249_n1088, CO => mult_21_C249_n680, S => 
                           mult_21_C249_n681);
   mult_21_C249_U1322 : ADHALFDL port map( A => mult_21_C249_n1206, B => 
                           mult_21_C249_n1090, CO => mult_21_C249_n732, S => 
                           mult_21_C249_n733);
   mult_21_C249_U1321 : INVD1 port map( A => mult_21_C249_n1557, Z => 
                           mult_21_C249_n1556);
   mult_21_C249_U1320 : INVD1 port map( A => mult_21_C249_n1555, Z => 
                           mult_21_C249_n1553);
   mult_21_C249_U1319 : INVD1 port map( A => mult_21_C249_n1550, Z => 
                           mult_21_C249_n1549);
   mult_21_C249_U1318 : INVD1 port map( A => mult_21_C249_n1552, Z => 
                           mult_21_C249_n1551);
   mult_21_C249_U1317 : INVD1 port map( A => mult_21_C249_n1544, Z => 
                           mult_21_C249_n1543);
   mult_21_C249_U1316 : INVD1 port map( A => mult_21_C249_n1555, Z => 
                           mult_21_C249_n1554);
   mult_21_C249_U1315 : INVD1 port map( A => mult_21_C249_n1548, Z => 
                           mult_21_C249_n1547);
   mult_21_C249_U1314 : INVD1 port map( A => mult_21_C249_n1542, Z => 
                           mult_21_C249_n1541);
   mult_21_C249_U1313 : INVD1 port map( A => mult_21_C249_n1546, Z => 
                           mult_21_C249_n1545);
   mult_21_C249_U1312 : INVD1 port map( A => mult_21_C249_n1537, Z => 
                           mult_21_C249_n1538);
   mult_21_C249_U1311 : ADHALFDL port map( A => mult_21_C249_n1306, B => 
                           mult_21_C249_n1094, CO => mult_21_C249_n788, S => 
                           mult_21_C249_n789);
   mult_21_C249_U1310 : ADHALFDL port map( A => mult_21_C249_n1333, B => 
                           mult_21_C249_n1363, CO => mult_21_C249_n784, S => 
                           mult_21_C249_n785);
   mult_21_C249_U1309 : ADHALFDL port map( A => mult_21_C249_n1252, B => 
                           mult_21_C249_n1092, CO => mult_21_C249_n768, S => 
                           mult_21_C249_n769);
   mult_21_C249_U1308 : ADHALFDL port map( A => mult_21_C249_n1331, B => 
                           mult_21_C249_n1361, CO => mult_21_C249_n774, S => 
                           mult_21_C249_n775);
   mult_21_C249_U1307 : INVD1 port map( A => mult_21_C249_n1536, Z => 
                           mult_21_C249_n1539);
   mult_21_C249_U1306 : NOR2D1 port map( A1 => mult_21_C249_n1537, A2 => 
                           mult_21_C249_n30, Z => mult_21_C249_n1093);
   mult_21_C249_U1305 : ADHALFDL port map( A => mult_21_C249_n1336, B => 
                           mult_21_C249_n1095, CO => mult_21_C249_n792, S => 
                           mult_21_C249_n793);
   mult_21_C249_U1304 : ADHALFDL port map( A => mult_21_C249_n1335, B => 
                           mult_21_C249_n1365, CO => mult_21_C249_n790, S => 
                           mult_21_C249_n791);
   mult_21_C249_U1303 : INVD1 port map( A => mult_21_C249_n1535, Z => 
                           mult_21_C249_n1540);
   mult_21_C249_U1302 : ADHALFDL port map( A => mult_21_C249_n1329, B => 
                           mult_21_C249_n1359, CO => mult_21_C249_n760, S => 
                           mult_21_C249_n761);
   mult_21_C249_U1301 : NOR2D1 port map( A1 => mult_21_C249_n303, A2 => 
                           mult_21_C249_n305, Z => mult_21_C249_n302);
   mult_21_C249_U1300 : NAN2D1 port map( A1 => mult_21_C249_n1368, A2 => 
                           mult_21_C249_n1096, Z => mult_21_C249_n305);
   mult_21_C249_U1299 : NAN2D1 port map( A1 => mult_21_C249_n791, A2 => 
                           mult_21_C249_n792, Z => mult_21_C249_n296);
   mult_21_C249_U1298 : NAN2D1 port map( A1 => mult_21_C249_n783, A2 => 
                           mult_21_C249_n786, Z => mult_21_C249_n288);
   mult_21_C249_U1297 : NOR2D1 port map( A1 => mult_21_C249_n791, A2 => 
                           mult_21_C249_n792, Z => mult_21_C249_n295);
   mult_21_C249_U1296 : NOR2D1 port map( A1 => mult_21_C249_n783, A2 => 
                           mult_21_C249_n786, Z => mult_21_C249_n287);
   mult_21_C249_U1295 : NAN2D1 port map( A1 => mult_21_C249_n777, A2 => 
                           mult_21_C249_n782, Z => mult_21_C249_n284);
   mult_21_C249_U1294 : NAN2D1 port map( A1 => mult_21_C249_n793, A2 => 
                           mult_21_C249_n1366, Z => mult_21_C249_n301);
   mult_21_C249_U1293 : NAN2D1 port map( A1 => mult_21_C249_n787, A2 => 
                           mult_21_C249_n789, Z => mult_21_C249_n293);
   mult_21_C249_U1292 : NOR2D1 port map( A1 => mult_21_C249_n777, A2 => 
                           mult_21_C249_n782, Z => mult_21_C249_n283);
   mult_21_C249_U1291 : OR2D1 port map( A1 => mult_21_C249_n793, A2 => 
                           mult_21_C249_n1366, Z => mult_21_C249_n1534);
   mult_21_C249_U1290 : OR2D1 port map( A1 => mult_21_C249_n787, A2 => 
                           mult_21_C249_n789, Z => mult_21_C249_n1533);
   mult_21_C249_U1289 : EXOR2D1 port map( A1 => mult_21_C249_n329, A2 => 
                           mult_21_C249_n344, Z => mult_21_C249_n155);
   mult_21_C249_U1288 : EXOR2D1 port map( A1 => mult_21_C249_n178, A2 => 
                           mult_21_C249_n155, Z => N3392);
   mult_21_C249_U1287 : NAN2D1 port map( A1 => mult_21_C249_n1534, A2 => 
                           mult_21_C249_n301, Z => mult_21_C249_n176);
   mult_21_C249_U1286 : INVD1 port map( A => mult_21_C249_n295, Z => 
                           mult_21_C249_n326);
   mult_21_C249_U1285 : NAN2D1 port map( A1 => mult_21_C249_n326, A2 => 
                           mult_21_C249_n296, Z => mult_21_C249_n175);
   mult_21_C249_U1284 : NAN2D1 port map( A1 => mult_21_C249_n1533, A2 => 
                           mult_21_C249_n293, Z => mult_21_C249_n174);
   mult_21_C249_U1283 : INVD1 port map( A => mult_21_C249_n287, Z => 
                           mult_21_C249_n324);
   mult_21_C249_U1282 : NAN2D1 port map( A1 => mult_21_C249_n324, A2 => 
                           mult_21_C249_n288, Z => mult_21_C249_n173);
   mult_21_C249_U1281 : INVD1 port map( A => mult_21_C249_n283, Z => 
                           mult_21_C249_n323);
   mult_21_C249_U1280 : NAN2D1 port map( A1 => mult_21_C249_n323, A2 => 
                           mult_21_C249_n284, Z => mult_21_C249_n172);
   mult_21_C249_U1279 : INVD1 port map( A => mult_21_C249_n280, Z => 
                           mult_21_C249_n322);
   mult_21_C249_U1278 : NAN2D1 port map( A1 => mult_21_C249_n322, A2 => 
                           mult_21_C249_n281, Z => mult_21_C249_n171);
   mult_21_C249_U1277 : NAN2D1 port map( A1 => mult_21_C249_n697, A2 => 
                           mult_21_C249_n710, Z => mult_21_C249_n240);
   mult_21_C249_U1276 : NAN2D1 port map( A1 => mult_21_C249_n711, A2 => 
                           mult_21_C249_n722, Z => mult_21_C249_n248);
   mult_21_C249_U1275 : NAN2D1 port map( A1 => mult_21_C249_n633, A2 => 
                           mult_21_C249_n650, Z => mult_21_C249_n221);
   mult_21_C249_U1274 : NOR2D1 port map( A1 => mult_21_C249_n615, A2 => 
                           mult_21_C249_n632, Z => mult_21_C249_n208);
   mult_21_C249_U1273 : NOR2D1 port map( A1 => mult_21_C249_n697, A2 => 
                           mult_21_C249_n710, Z => mult_21_C249_n239);
   mult_21_C249_U1272 : NAN2D1 port map( A1 => mult_21_C249_n735, A2 => 
                           mult_21_C249_n744, Z => mult_21_C249_n259);
   mult_21_C249_U1271 : NAN2D1 port map( A1 => mult_21_C249_n615, A2 => 
                           mult_21_C249_n632, Z => mult_21_C249_n209);
   mult_21_C249_U1270 : NAN2D1 port map( A1 => mult_21_C249_n771, A2 => 
                           mult_21_C249_n776, Z => mult_21_C249_n281);
   mult_21_C249_U1269 : OR2D1 port map( A1 => mult_21_C249_n711, A2 => 
                           mult_21_C249_n722, Z => mult_21_C249_n1532);
   mult_21_C249_U1268 : OR2D1 port map( A1 => mult_21_C249_n723, A2 => 
                           mult_21_C249_n734, Z => mult_21_C249_n1531);
   mult_21_C249_U1267 : NAN2D1 port map( A1 => mult_21_C249_n745, A2 => 
                           mult_21_C249_n754, Z => mult_21_C249_n262);
   mult_21_C249_U1266 : OR2D1 port map( A1 => mult_21_C249_n633, A2 => 
                           mult_21_C249_n650, Z => mult_21_C249_n1530);
   mult_21_C249_U1265 : NAN2D1 port map( A1 => mult_21_C249_n595, A2 => 
                           mult_21_C249_n614, Z => mult_21_C249_n206);
   mult_21_C249_U1264 : OR2D1 port map( A1 => mult_21_C249_n763, A2 => 
                           mult_21_C249_n770, Z => mult_21_C249_n1529);
   mult_21_C249_U1263 : NAN2D1 port map( A1 => mult_21_C249_n651, A2 => 
                           mult_21_C249_n666, Z => mult_21_C249_n226);
   mult_21_C249_U1262 : NAN2D1 port map( A1 => mult_21_C249_n723, A2 => 
                           mult_21_C249_n734, Z => mult_21_C249_n253);
   mult_21_C249_U1261 : NAN2D1 port map( A1 => mult_21_C249_n575, A2 => 
                           mult_21_C249_n594, Z => mult_21_C249_n199);
   mult_21_C249_U1260 : OR2D1 port map( A1 => mult_21_C249_n575, A2 => 
                           mult_21_C249_n594, Z => mult_21_C249_n1528);
   mult_21_C249_U1259 : NAN2D1 port map( A1 => mult_21_C249_n763, A2 => 
                           mult_21_C249_n770, Z => mult_21_C249_n275);
   mult_21_C249_U1258 : NOR2D1 port map( A1 => mult_21_C249_n735, A2 => 
                           mult_21_C249_n744, Z => mult_21_C249_n258);
   mult_21_C249_U1257 : NOR2D1 port map( A1 => mult_21_C249_n745, A2 => 
                           mult_21_C249_n754, Z => mult_21_C249_n261);
   mult_21_C249_U1256 : NOR2D1 port map( A1 => mult_21_C249_n771, A2 => 
                           mult_21_C249_n776, Z => mult_21_C249_n280);
   mult_21_C249_U1255 : OR2D1 port map( A1 => mult_21_C249_n595, A2 => 
                           mult_21_C249_n614, Z => mult_21_C249_n1527);
   mult_21_C249_U1254 : OA21M20D1 port map( A1 => mult_21_C249_n1534, A2 => 
                           mult_21_C249_n302, B => mult_21_C249_n301, Z => 
                           mult_21_C249_n297);
   mult_21_C249_U1253 : NOR2D1 port map( A1 => mult_21_C249_n651, A2 => 
                           mult_21_C249_n666, Z => mult_21_C249_n225);
   mult_21_C249_U1252 : OA21M20D1 port map( A1 => mult_21_C249_n1533, A2 => 
                           mult_21_C249_n294, B => mult_21_C249_n293, Z => 
                           mult_21_C249_n289);
   mult_21_C249_U1251 : NOR2D1 port map( A1 => mult_21_C249_n280, A2 => 
                           mult_21_C249_n283, Z => mult_21_C249_n278);
   mult_21_C249_U1250 : NAN2D1 port map( A1 => mult_21_C249_n755, A2 => 
                           mult_21_C249_n762, Z => mult_21_C249_n270);
   mult_21_C249_U1249 : OR2D1 port map( A1 => mult_21_C249_n755, A2 => 
                           mult_21_C249_n762, Z => mult_21_C249_n1526);
   mult_21_C249_U1248 : INVD1 port map( A => mult_21_C249_n286, Z => 
                           mult_21_C249_n285);
   mult_21_C249_U1247 : NAN2D1 port map( A1 => mult_21_C249_n1529, A2 => 
                           mult_21_C249_n275, Z => mult_21_C249_n170);
   mult_21_C249_U1246 : NAN2D1 port map( A1 => mult_21_C249_n1526, A2 => 
                           mult_21_C249_n270, Z => mult_21_C249_n169);
   mult_21_C249_U1245 : INVD1 port map( A => mult_21_C249_n277, Z => 
                           mult_21_C249_n276);
   mult_21_C249_U1244 : INVD1 port map( A => mult_21_C249_n261, Z => 
                           mult_21_C249_n319);
   mult_21_C249_U1243 : NAN2D1 port map( A1 => mult_21_C249_n319, A2 => 
                           mult_21_C249_n262, Z => mult_21_C249_n168);
   mult_21_C249_U1242 : INVD1 port map( A => mult_21_C249_n258, Z => 
                           mult_21_C249_n318);
   mult_21_C249_U1241 : NAN2D1 port map( A1 => mult_21_C249_n318, A2 => 
                           mult_21_C249_n259, Z => mult_21_C249_n167);
   mult_21_C249_U1240 : NAN2D1 port map( A1 => mult_21_C249_n1531, A2 => 
                           mult_21_C249_n253, Z => mult_21_C249_n166);
   mult_21_C249_U1239 : INVD1 port map( A => mult_21_C249_n239, Z => 
                           mult_21_C249_n315);
   mult_21_C249_U1238 : NAN2D1 port map( A1 => mult_21_C249_n315, A2 => 
                           mult_21_C249_n240, Z => mult_21_C249_n164);
   mult_21_C249_U1237 : NAN2D1 port map( A1 => mult_21_C249_n1532, A2 => 
                           mult_21_C249_n248, Z => mult_21_C249_n165);
   mult_21_C249_U1236 : INVD1 port map( A => mult_21_C249_n236, Z => 
                           mult_21_C249_n314);
   mult_21_C249_U1235 : NAN2D1 port map( A1 => mult_21_C249_n314, A2 => 
                           mult_21_C249_n237, Z => mult_21_C249_n163);
   mult_21_C249_U1234 : NAN2D1 port map( A1 => mult_21_C249_n1530, A2 => 
                           mult_21_C249_n221, Z => mult_21_C249_n160);
   mult_21_C249_U1233 : INVD1 port map( A => mult_21_C249_n225, Z => 
                           mult_21_C249_n312);
   mult_21_C249_U1232 : NAN2D1 port map( A1 => mult_21_C249_n312, A2 => 
                           mult_21_C249_n226, Z => mult_21_C249_n161);
   mult_21_C249_U1231 : NAN2D1 port map( A1 => mult_21_C249_n310, A2 => 
                           mult_21_C249_n209, Z => mult_21_C249_n159);
   mult_21_C249_U1230 : NAN2D1 port map( A1 => mult_21_C249_n1527, A2 => 
                           mult_21_C249_n206, Z => mult_21_C249_n158);
   mult_21_C249_U1229 : NAN2D1 port map( A1 => mult_21_C249_n1528, A2 => 
                           mult_21_C249_n199, Z => mult_21_C249_n157);
   mult_21_C249_U1228 : NAN2D1 port map( A1 => mult_21_C249_n1525, A2 => 
                           mult_21_C249_n194, Z => mult_21_C249_n156);
   mult_21_C249_U1227 : NAN2D1 port map( A1 => mult_21_C249_n683, A2 => 
                           mult_21_C249_n696, Z => mult_21_C249_n237);
   mult_21_C249_U1226 : INVD1 port map( A => mult_21_C249_n208, Z => 
                           mult_21_C249_n310);
   mult_21_C249_U1225 : NOR2D1 port map( A1 => mult_21_C249_n667, A2 => 
                           mult_21_C249_n682, Z => mult_21_C249_n230);
   mult_21_C249_U1224 : NAN2D1 port map( A1 => mult_21_C249_n553, A2 => 
                           mult_21_C249_n574, Z => mult_21_C249_n194);
   mult_21_C249_U1223 : NOR2D1 port map( A1 => mult_21_C249_n683, A2 => 
                           mult_21_C249_n696, Z => mult_21_C249_n236);
   mult_21_C249_U1222 : NAN2D1 port map( A1 => mult_21_C249_n1527, A2 => 
                           mult_21_C249_n310, Z => mult_21_C249_n201);
   mult_21_C249_U1221 : NOR2D1 port map( A1 => mult_21_C249_n225, A2 => 
                           mult_21_C249_n230, Z => mult_21_C249_n223);
   mult_21_C249_U1220 : INVD1 port map( A => mult_21_C249_n253, Z => 
                           mult_21_C249_n251);
   mult_21_C249_U1219 : NAN2D1 port map( A1 => mult_21_C249_n667, A2 => 
                           mult_21_C249_n682, Z => mult_21_C249_n231);
   mult_21_C249_U1218 : INVD1 port map( A => mult_21_C249_n199, Z => 
                           mult_21_C249_n197);
   mult_21_C249_U1217 : NAN2D1 port map( A1 => mult_21_C249_n1525, A2 => 
                           mult_21_C249_n1528, Z => mult_21_C249_n189);
   mult_21_C249_U1216 : OR2D1 port map( A1 => mult_21_C249_n553, A2 => 
                           mult_21_C249_n574, Z => mult_21_C249_n1525);
   mult_21_C249_U1215 : INVD1 port map( A => mult_21_C249_n275, Z => 
                           mult_21_C249_n273);
   mult_21_C249_U1214 : INVD1 port map( A => mult_21_C249_n206, Z => 
                           mult_21_C249_n204);
   mult_21_C249_U1213 : INVD1 port map( A => mult_21_C249_n209, Z => 
                           mult_21_C249_n211);
   mult_21_C249_U1212 : NOR2D1 port map( A1 => mult_21_C249_n189, A2 => 
                           mult_21_C249_n201, Z => mult_21_C249_n187);
   mult_21_C249_U1211 : NOR2D1 port map( A1 => mult_21_C249_n236, A2 => 
                           mult_21_C249_n239, Z => mult_21_C249_n234);
   mult_21_C249_U1210 : NOR2D1 port map( A1 => mult_21_C249_n258, A2 => 
                           mult_21_C249_n261, Z => mult_21_C249_n256);
   mult_21_C249_U1209 : INVD1 port map( A => mult_21_C249_n270, Z => 
                           mult_21_C249_n268);
   mult_21_C249_U1208 : NAN2D1 port map( A1 => mult_21_C249_n1526, A2 => 
                           mult_21_C249_n1529, Z => mult_21_C249_n265);
   mult_21_C249_U1207 : INVD1 port map( A => mult_21_C249_n248, Z => 
                           mult_21_C249_n246);
   mult_21_C249_U1206 : NAN2D1 port map( A1 => mult_21_C249_n1532, A2 => 
                           mult_21_C249_n1531, Z => mult_21_C249_n243);
   mult_21_C249_U1205 : INVD1 port map( A => mult_21_C249_n221, Z => 
                           mult_21_C249_n219);
   mult_21_C249_U1204 : NAN2D1 port map( A1 => mult_21_C249_n223, A2 => 
                           mult_21_C249_n1530, Z => mult_21_C249_n216);
   mult_21_C249_U1203 : INVD1 port map( A => mult_21_C249_n264, Z => 
                           mult_21_C249_n263);
   mult_21_C249_U1202 : INVD1 port map( A => mult_21_C249_n231, Z => 
                           mult_21_C249_n229);
   mult_21_C249_U1201 : INVD1 port map( A => mult_21_C249_n230, Z => 
                           mult_21_C249_n313);
   mult_21_C249_U1200 : INVD1 port map( A => mult_21_C249_n255, Z => 
                           mult_21_C249_n254);
   mult_21_C249_U1199 : INVD1 port map( A => mult_21_C249_n242, Z => 
                           mult_21_C249_n241);
   mult_21_C249_U1198 : NAN2D1 port map( A1 => mult_21_C249_n313, A2 => 
                           mult_21_C249_n231, Z => mult_21_C249_n162);
   mult_21_C249_U1197 : INVD1 port map( A => mult_21_C249_n233, Z => 
                           mult_21_C249_n232);
   mult_21_C249_U1196 : INVD1 port map( A => mult_21_C249_n215, Z => 
                           mult_21_C249_n214);
   mult_21_C249_U1195 : OA21M20D1 port map( A1 => mult_21_C249_n1525, A2 => 
                           mult_21_C249_n197, B => mult_21_C249_n194, Z => 
                           mult_21_C249_n190);
   mult_21_C249_U1194 : OR2D1 port map( A1 => mult_21_C249_n1368, A2 => 
                           mult_21_C249_n1096, Z => mult_21_C249_n1524);
   mult_21_C249_U1193 : AO21D1 port map( A1 => mult_21_C249_n215, A2 => 
                           mult_21_C249_n187, B => mult_21_C249_n188, Z => 
                           mult_21_C249_n1523);
   mult_21_C249_U1192 : AND2D1 port map( A1 => mult_21_C249_n1524, A2 => 
                           mult_21_C249_n305, Z => N3361);
   mult_21_C249_U1191 : OAI21D1 port map( A1 => N3048, A2 => N3049, B => 
                           mult_21_C249_n1077, Z => mult_21_C249_n1521);
   mult_21_C249_U1190 : OAI21D1 port map( A1 => N3044, A2 => N3045, B => 
                           mult_21_C249_n1079, Z => mult_21_C249_n1520);
   mult_21_C249_U1189 : OAI21D1 port map( A1 => N3042, A2 => N3043, B => 
                           mult_21_C249_n1080, Z => mult_21_C249_n1519);
   mult_21_C249_U1188 : EXNOR2D1 port map( A1 => N3048, A2 => N3049, Z => 
                           mult_21_C249_n1518);
   mult_21_C249_U1187 : EXNOR2D1 port map( A1 => N3046, A2 => N3047, Z => 
                           mult_21_C249_n1517);
   mult_21_C249_U1186 : ADHALFDL port map( A => mult_21_C249_n1278, B => 
                           mult_21_C249_n1093, CO => mult_21_C249_n780, S => 
                           mult_21_C249_n781);
   mult_21_C249_U1135 : EXNOR2D1 port map( A1 => N3064, A2 => N3065, Z => 
                           mult_21_C249_n93);
   mult_21_C249_U1131 : EXNOR2D1 port map( A1 => N3066, A2 => N3067, Z => 
                           mult_21_C249_n98);
   mult_21_C249_U1129 : OAI21D1 port map( A1 => N3066, A2 => N3067, B => 
                           mult_21_C249_n1068, Z => mult_21_C249_n94);
   mult_21_C249_U1127 : EXNOR2D1 port map( A1 => N3068, A2 => N3069, Z => 
                           mult_21_C249_n103);
   mult_21_C249_U1125 : OAI21D1 port map( A1 => N3068, A2 => N3069, B => 
                           mult_21_C249_n1067, Z => mult_21_C249_n99);
   mult_21_C249_U1123 : EXNOR2D1 port map( A1 => N3070, A2 => N3071, Z => 
                           mult_21_C249_n106);
   mult_21_C249_U1121 : OAI21D1 port map( A1 => N3070, A2 => N3071, B => 
                           mult_21_C249_n1066, Z => mult_21_C249_n104);
   mult_21_C249_U1120 : NAN2M1D1 port map( A1 => mult_21_C249_n8, A2 => n288, Z
                           => mult_21_C249_n1065);
   mult_21_C249_U1119 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1065, Z => 
                           mult_21_C249_n1368);
   mult_21_C249_U1118 : MUXB2DL port map( A0 => mult_21_C249_n1553, A1 => n288,
                           SL => mult_21_C249_n8, Z => mult_21_C249_n1064);
   mult_21_C249_U1117 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1064, Z => 
                           mult_21_C249_n1367);
   mult_21_C249_U1116 : MUXB2DL port map( A0 => n284, A1 => mult_21_C249_n1554,
                           SL => mult_21_C249_n8, Z => mult_21_C249_n1063);
   mult_21_C249_U1115 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1063, Z => 
                           mult_21_C249_n1366);
   mult_21_C249_U1114 : MUXB2DL port map( A0 => mult_21_C249_n1551, A1 => n284,
                           SL => mult_21_C249_n8, Z => mult_21_C249_n1062);
   mult_21_C249_U1113 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1062, Z => 
                           mult_21_C249_n1365);
   mult_21_C249_U1112 : MUXB2DL port map( A0 => n287, A1 => n286, SL => 
                           mult_21_C249_n8, Z => mult_21_C249_n1061);
   mult_21_C249_U1111 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1061, Z => 
                           mult_21_C249_n1364);
   mult_21_C249_U1110 : MUXB2DL port map( A0 => n282, A1 => mult_21_C249_n1549,
                           SL => mult_21_C249_n8, Z => mult_21_C249_n1060);
   mult_21_C249_U1109 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1060, Z => 
                           mult_21_C249_n1363);
   mult_21_C249_U1108 : MUXB2DL port map( A0 => n278, A1 => mult_21_C249_n1547,
                           SL => mult_21_C249_n8, Z => mult_21_C249_n1059);
   mult_21_C249_U1107 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1059, Z => 
                           mult_21_C249_n1362);
   mult_21_C249_U1106 : MUXB2DL port map( A0 => n279, A1 => mult_21_C249_n1545,
                           SL => mult_21_C249_n8, Z => mult_21_C249_n1058);
   mult_21_C249_U1105 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1058, Z => 
                           mult_21_C249_n1361);
   mult_21_C249_U1104 : MUXB2DL port map( A0 => n280, A1 => mult_21_C249_n1543,
                           SL => mult_21_C249_n8, Z => mult_21_C249_n1057);
   mult_21_C249_U1103 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1057, Z => 
                           mult_21_C249_n1360);
   mult_21_C249_U1102 : MUXB2DL port map( A0 => mult_21_C249_n1541, A1 => n280,
                           SL => mult_21_C249_n8, Z => mult_21_C249_n1056);
   mult_21_C249_U1101 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1056, Z => 
                           mult_21_C249_n1359);
   mult_21_C249_U1100 : MUXB2DL port map( A0 => n285, A1 => n281, SL => 
                           mult_21_C249_n8, Z => mult_21_C249_n1055);
   mult_21_C249_U1099 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1055, Z => 
                           mult_21_C249_n1358);
   mult_21_C249_U1098 : MUXB2DL port map( A0 => n274, A1 => n285, SL => 
                           mult_21_C249_n8, Z => mult_21_C249_n1054);
   mult_21_C249_U1097 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1054, Z => 
                           mult_21_C249_n1357);
   mult_21_C249_U1096 : MUXB2DL port map( A0 => n271, A1 => n274, SL => 
                           mult_21_C249_n8, Z => mult_21_C249_n1053);
   mult_21_C249_U1095 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1053, Z => 
                           mult_21_C249_n1356);
   mult_21_C249_U1094 : MUXB2DL port map( A0 => n272, A1 => n271, SL => 
                           mult_21_C249_n8, Z => mult_21_C249_n1052);
   mult_21_C249_U1093 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1052, Z => 
                           mult_21_C249_n1355);
   mult_21_C249_U1092 : MUXB2DL port map( A0 => n273, A1 => n272, SL => 
                           mult_21_C249_n8, Z => mult_21_C249_n1051);
   mult_21_C249_U1091 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1051, Z => 
                           mult_21_C249_n1354);
   mult_21_C249_U1090 : MUXB2DL port map( A0 => n291, A1 => n273, SL => 
                           mult_21_C249_n8, Z => mult_21_C249_n1050);
   mult_21_C249_U1089 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1050, Z => 
                           mult_21_C249_n1353);
   mult_21_C249_U1088 : MUXB2DL port map( A0 => n292, A1 => n291, SL => 
                           mult_21_C249_n8, Z => mult_21_C249_n1049);
   mult_21_C249_U1087 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1049, Z => 
                           mult_21_C249_n1352);
   mult_21_C249_U1086 : MUXB2DL port map( A0 => n289, A1 => n292, SL => 
                           mult_21_C249_n8, Z => mult_21_C249_n1048);
   mult_21_C249_U1085 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1048, Z => 
                           mult_21_C249_n1351);
   mult_21_C249_U1084 : MUXB2DL port map( A0 => n290, A1 => n289, SL => 
                           mult_21_C249_n8, Z => mult_21_C249_n1047);
   mult_21_C249_U1083 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1047, Z => 
                           mult_21_C249_n1350);
   mult_21_C249_U1082 : MUXB2DL port map( A0 => n293, A1 => n290, SL => 
                           mult_21_C249_n8, Z => mult_21_C249_n1046);
   mult_21_C249_U1081 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1046, Z => 
                           mult_21_C249_n1349);
   mult_21_C249_U1080 : MUXB2DL port map( A0 => n294, A1 => n293, SL => 
                           mult_21_C249_n8, Z => mult_21_C249_n1045);
   mult_21_C249_U1079 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1045, Z => 
                           mult_21_C249_n1348);
   mult_21_C249_U1078 : MUXB2DL port map( A0 => n295, A1 => n294, SL => 
                           mult_21_C249_n8, Z => mult_21_C249_n1044);
   mult_21_C249_U1077 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1044, Z => 
                           mult_21_C249_n1347);
   mult_21_C249_U1076 : MUXB2DL port map( A0 => n296, A1 => n295, SL => 
                           mult_21_C249_n8, Z => mult_21_C249_n1043);
   mult_21_C249_U1075 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1043, Z => 
                           mult_21_C249_n1346);
   mult_21_C249_U1074 : MUXB2DL port map( A0 => n297, A1 => n296, SL => 
                           mult_21_C249_n8, Z => mult_21_C249_n1042);
   mult_21_C249_U1073 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1042, Z => 
                           mult_21_C249_n1345);
   mult_21_C249_U1072 : MUXB2DL port map( A0 => n298, A1 => n297, SL => 
                           mult_21_C249_n8, Z => mult_21_C249_n1041);
   mult_21_C249_U1071 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1041, Z => 
                           mult_21_C249_n1344);
   mult_21_C249_U1070 : MUXB2DL port map( A0 => n299, A1 => n298, SL => 
                           mult_21_C249_n8, Z => mult_21_C249_n1040);
   mult_21_C249_U1069 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1040, Z => 
                           mult_21_C249_n1343);
   mult_21_C249_U1068 : MUXB2DL port map( A0 => n302, A1 => n299, SL => 
                           mult_21_C249_n8, Z => mult_21_C249_n1039);
   mult_21_C249_U1067 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1039, Z => 
                           mult_21_C249_n1342);
   mult_21_C249_U1066 : MUXB2DL port map( A0 => n303, A1 => n302, SL => 
                           mult_21_C249_n8, Z => mult_21_C249_n1038);
   mult_21_C249_U1065 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1038, Z => 
                           mult_21_C249_n1341);
   mult_21_C249_U1064 : MUXB2DL port map( A0 => n305, A1 => n303, SL => 
                           mult_21_C249_n8, Z => mult_21_C249_n1037);
   mult_21_C249_U1063 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1037, Z => 
                           mult_21_C249_n1340);
   mult_21_C249_U1062 : MUXB2DL port map( A0 => n310, A1 => n305, SL => 
                           mult_21_C249_n8, Z => mult_21_C249_n1036);
   mult_21_C249_U1061 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1036, Z => 
                           mult_21_C249_n1339);
   mult_21_C249_U1060 : MUXB2DL port map( A0 => n311, A1 => n310, SL => 
                           mult_21_C249_n8, Z => mult_21_C249_n1035);
   mult_21_C249_U1059 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1035, Z => 
                           mult_21_C249_n1338);
   mult_21_C249_U1058 : MUXB2DL port map( A0 => n312, A1 => n311, SL => 
                           mult_21_C249_n8, Z => mult_21_C249_n1034);
   mult_21_C249_U1057 : MUXB2DL port map( A0 => mult_21_C249_n3, A1 => 
                           mult_21_C249_n6, SL => mult_21_C249_n1034, Z => 
                           mult_21_C249_n1337);
   mult_21_C249_U1056 : NOR2M1D1 port map( A1 => mult_21_C249_n3, A2 => 
                           mult_21_C249_n6, Z => mult_21_C249_n1096);
   mult_21_C249_U1055 : NAN2M1D1 port map( A1 => mult_21_C249_n1540, A2 => 
                           mult_21_C249_n1556, Z => mult_21_C249_n1033);
   mult_21_C249_U1054 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1033, Z => 
                           mult_21_C249_n1336);
   mult_21_C249_U1053 : MUXB2DL port map( A0 => mult_21_C249_n1553, A1 => n288,
                           SL => mult_21_C249_n1540, Z => mult_21_C249_n1032);
   mult_21_C249_U1052 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1032, Z => 
                           mult_21_C249_n1335);
   mult_21_C249_U1051 : MUXB2DL port map( A0 => n284, A1 => mult_21_C249_n1554,
                           SL => mult_21_C249_n1540, Z => mult_21_C249_n1031);
   mult_21_C249_U1050 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1031, Z => 
                           mult_21_C249_n1334);
   mult_21_C249_U1049 : MUXB2DL port map( A0 => mult_21_C249_n1551, A1 => n284,
                           SL => mult_21_C249_n1540, Z => mult_21_C249_n1030);
   mult_21_C249_U1048 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1030, Z => 
                           mult_21_C249_n1333);
   mult_21_C249_U1047 : MUXB2DL port map( A0 => n287, A1 => n286, SL => 
                           mult_21_C249_n1540, Z => mult_21_C249_n1029);
   mult_21_C249_U1046 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1029, Z => 
                           mult_21_C249_n1332);
   mult_21_C249_U1045 : MUXB2DL port map( A0 => n282, A1 => mult_21_C249_n1549,
                           SL => mult_21_C249_n1540, Z => mult_21_C249_n1028);
   mult_21_C249_U1044 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1028, Z => 
                           mult_21_C249_n1331);
   mult_21_C249_U1043 : MUXB2DL port map( A0 => n278, A1 => mult_21_C249_n1547,
                           SL => mult_21_C249_n1540, Z => mult_21_C249_n1027);
   mult_21_C249_U1042 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1027, Z => 
                           mult_21_C249_n1330);
   mult_21_C249_U1041 : MUXB2DL port map( A0 => mult_21_C249_n1543, A1 => 
                           mult_21_C249_n1545, SL => mult_21_C249_n1540, Z => 
                           mult_21_C249_n1026);
   mult_21_C249_U1040 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1026, Z => 
                           mult_21_C249_n1329);
   mult_21_C249_U1039 : MUXB2DL port map( A0 => n280, A1 => mult_21_C249_n1543,
                           SL => mult_21_C249_n1540, Z => mult_21_C249_n1025);
   mult_21_C249_U1038 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1025, Z => 
                           mult_21_C249_n1328);
   mult_21_C249_U1037 : MUXB2DL port map( A0 => mult_21_C249_n1541, A1 => n280,
                           SL => mult_21_C249_n1540, Z => mult_21_C249_n1024);
   mult_21_C249_U1036 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1024, Z => 
                           mult_21_C249_n1327);
   mult_21_C249_U1035 : MUXB2DL port map( A0 => n285, A1 => n281, SL => 
                           mult_21_C249_n1540, Z => mult_21_C249_n1023);
   mult_21_C249_U1034 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1023, Z => 
                           mult_21_C249_n1326);
   mult_21_C249_U1033 : MUXB2DL port map( A0 => n274, A1 => n285, SL => 
                           mult_21_C249_n1540, Z => mult_21_C249_n1022);
   mult_21_C249_U1032 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1022, Z => 
                           mult_21_C249_n1325);
   mult_21_C249_U1031 : MUXB2DL port map( A0 => n271, A1 => n274, SL => 
                           mult_21_C249_n1540, Z => mult_21_C249_n1021);
   mult_21_C249_U1030 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1021, Z => 
                           mult_21_C249_n1324);
   mult_21_C249_U1029 : MUXB2DL port map( A0 => n272, A1 => n271, SL => 
                           mult_21_C249_n1540, Z => mult_21_C249_n1020);
   mult_21_C249_U1028 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1020, Z => 
                           mult_21_C249_n1323);
   mult_21_C249_U1027 : MUXB2DL port map( A0 => n273, A1 => n272, SL => 
                           mult_21_C249_n1540, Z => mult_21_C249_n1019);
   mult_21_C249_U1026 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1019, Z => 
                           mult_21_C249_n1322);
   mult_21_C249_U1025 : MUXB2DL port map( A0 => n291, A1 => n273, SL => 
                           mult_21_C249_n1540, Z => mult_21_C249_n1018);
   mult_21_C249_U1024 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1018, Z => 
                           mult_21_C249_n1321);
   mult_21_C249_U1023 : MUXB2DL port map( A0 => n292, A1 => n291, SL => 
                           mult_21_C249_n1540, Z => mult_21_C249_n1017);
   mult_21_C249_U1022 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1017, Z => 
                           mult_21_C249_n1320);
   mult_21_C249_U1021 : MUXB2DL port map( A0 => n289, A1 => n292, SL => 
                           mult_21_C249_n1540, Z => mult_21_C249_n1016);
   mult_21_C249_U1020 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1016, Z => 
                           mult_21_C249_n1319);
   mult_21_C249_U1019 : MUXB2DL port map( A0 => n290, A1 => n289, SL => 
                           mult_21_C249_n1540, Z => mult_21_C249_n1015);
   mult_21_C249_U1018 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1015, Z => 
                           mult_21_C249_n1318);
   mult_21_C249_U1017 : MUXB2DL port map( A0 => n293, A1 => n290, SL => 
                           mult_21_C249_n1540, Z => mult_21_C249_n1014);
   mult_21_C249_U1016 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1014, Z => 
                           mult_21_C249_n1317);
   mult_21_C249_U1015 : MUXB2DL port map( A0 => n294, A1 => n293, SL => 
                           mult_21_C249_n1540, Z => mult_21_C249_n1013);
   mult_21_C249_U1014 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1013, Z => 
                           mult_21_C249_n1316);
   mult_21_C249_U1013 : MUXB2DL port map( A0 => n295, A1 => n294, SL => 
                           mult_21_C249_n1540, Z => mult_21_C249_n1012);
   mult_21_C249_U1012 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1012, Z => 
                           mult_21_C249_n1315);
   mult_21_C249_U1011 : MUXB2DL port map( A0 => n296, A1 => n295, SL => 
                           mult_21_C249_n1540, Z => mult_21_C249_n1011);
   mult_21_C249_U1010 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1011, Z => 
                           mult_21_C249_n1314);
   mult_21_C249_U1009 : MUXB2DL port map( A0 => n297, A1 => n296, SL => 
                           mult_21_C249_n1540, Z => mult_21_C249_n1010);
   mult_21_C249_U1008 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1010, Z => 
                           mult_21_C249_n1313);
   mult_21_C249_U1007 : MUXB2DL port map( A0 => n298, A1 => n297, SL => 
                           mult_21_C249_n1540, Z => mult_21_C249_n1009);
   mult_21_C249_U1006 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1009, Z => 
                           mult_21_C249_n1312);
   mult_21_C249_U1005 : MUXB2DL port map( A0 => n299, A1 => n298, SL => 
                           mult_21_C249_n1540, Z => mult_21_C249_n1008);
   mult_21_C249_U1004 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1008, Z => 
                           mult_21_C249_n1311);
   mult_21_C249_U1003 : MUXB2DL port map( A0 => n302, A1 => n299, SL => 
                           mult_21_C249_n1540, Z => mult_21_C249_n1007);
   mult_21_C249_U1002 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1007, Z => 
                           mult_21_C249_n1310);
   mult_21_C249_U1001 : MUXB2DL port map( A0 => n303, A1 => n302, SL => 
                           mult_21_C249_n1540, Z => mult_21_C249_n1006);
   mult_21_C249_U1000 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1006, Z => 
                           mult_21_C249_n1309);
   mult_21_C249_U999 : MUXB2DL port map( A0 => n305, A1 => n303, SL => 
                           mult_21_C249_n1540, Z => mult_21_C249_n1005);
   mult_21_C249_U998 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1005, Z => 
                           mult_21_C249_n1308);
   mult_21_C249_U997 : MUXB2DL port map( A0 => n310, A1 => n305, SL => 
                           mult_21_C249_n1540, Z => mult_21_C249_n1004);
   mult_21_C249_U996 : MUXB2DL port map( A0 => mult_21_C249_n1519, A1 => 
                           mult_21_C249_n14, SL => mult_21_C249_n1004, Z => 
                           mult_21_C249_n1307);
   mult_21_C249_U995 : NOR2M1D1 port map( A1 => mult_21_C249_n1519, A2 => 
                           mult_21_C249_n14, Z => mult_21_C249_n1095);
   mult_21_C249_U994 : NAN2M1D1 port map( A1 => mult_21_C249_n1539, A2 => 
                           mult_21_C249_n1556, Z => mult_21_C249_n1003);
   mult_21_C249_U993 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n1003, Z => 
                           mult_21_C249_n1306);
   mult_21_C249_U992 : MUXB2DL port map( A0 => mult_21_C249_n1553, A1 => 
                           mult_21_C249_n1556, SL => mult_21_C249_n1539, Z => 
                           mult_21_C249_n1002);
   mult_21_C249_U991 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n1002, Z => 
                           mult_21_C249_n1305);
   mult_21_C249_U990 : MUXB2DL port map( A0 => n284, A1 => mult_21_C249_n1554, 
                           SL => mult_21_C249_n1539, Z => mult_21_C249_n1001);
   mult_21_C249_U989 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n1001, Z => 
                           mult_21_C249_n1304);
   mult_21_C249_U988 : MUXB2DL port map( A0 => mult_21_C249_n1551, A1 => n284, 
                           SL => mult_21_C249_n1539, Z => mult_21_C249_n1000);
   mult_21_C249_U987 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n1000, Z => 
                           mult_21_C249_n1303);
   mult_21_C249_U986 : MUXB2DL port map( A0 => n287, A1 => n286, SL => 
                           mult_21_C249_n1539, Z => mult_21_C249_n999);
   mult_21_C249_U985 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n999, Z => 
                           mult_21_C249_n1302);
   mult_21_C249_U984 : MUXB2DL port map( A0 => n282, A1 => mult_21_C249_n1549, 
                           SL => mult_21_C249_n1539, Z => mult_21_C249_n998);
   mult_21_C249_U983 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n998, Z => 
                           mult_21_C249_n1301);
   mult_21_C249_U982 : MUXB2DL port map( A0 => n278, A1 => mult_21_C249_n1547, 
                           SL => mult_21_C249_n1539, Z => mult_21_C249_n997);
   mult_21_C249_U981 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n997, Z => 
                           mult_21_C249_n1300);
   mult_21_C249_U980 : MUXB2DL port map( A0 => n279, A1 => mult_21_C249_n1545, 
                           SL => mult_21_C249_n1539, Z => mult_21_C249_n996);
   mult_21_C249_U979 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n996, Z => 
                           mult_21_C249_n1299);
   mult_21_C249_U978 : MUXB2DL port map( A0 => n280, A1 => mult_21_C249_n1543, 
                           SL => mult_21_C249_n1539, Z => mult_21_C249_n995);
   mult_21_C249_U977 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n995, Z => 
                           mult_21_C249_n1298);
   mult_21_C249_U976 : MUXB2DL port map( A0 => mult_21_C249_n1541, A1 => n280, 
                           SL => mult_21_C249_n1539, Z => mult_21_C249_n994);
   mult_21_C249_U975 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n994, Z => 
                           mult_21_C249_n1297);
   mult_21_C249_U974 : MUXB2DL port map( A0 => n285, A1 => n281, SL => 
                           mult_21_C249_n1539, Z => mult_21_C249_n993);
   mult_21_C249_U973 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n993, Z => 
                           mult_21_C249_n1296);
   mult_21_C249_U972 : MUXB2DL port map( A0 => n274, A1 => n285, SL => 
                           mult_21_C249_n1539, Z => mult_21_C249_n992);
   mult_21_C249_U971 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n992, Z => 
                           mult_21_C249_n1295);
   mult_21_C249_U970 : MUXB2DL port map( A0 => n271, A1 => n274, SL => 
                           mult_21_C249_n1539, Z => mult_21_C249_n991);
   mult_21_C249_U969 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n991, Z => 
                           mult_21_C249_n1294);
   mult_21_C249_U968 : MUXB2DL port map( A0 => n272, A1 => n271, SL => 
                           mult_21_C249_n1539, Z => mult_21_C249_n990);
   mult_21_C249_U967 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n990, Z => 
                           mult_21_C249_n1293);
   mult_21_C249_U966 : MUXB2DL port map( A0 => n273, A1 => n272, SL => 
                           mult_21_C249_n1539, Z => mult_21_C249_n989);
   mult_21_C249_U965 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n989, Z => 
                           mult_21_C249_n1292);
   mult_21_C249_U964 : MUXB2DL port map( A0 => n291, A1 => n273, SL => 
                           mult_21_C249_n1539, Z => mult_21_C249_n988);
   mult_21_C249_U963 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n988, Z => 
                           mult_21_C249_n1291);
   mult_21_C249_U962 : MUXB2DL port map( A0 => n292, A1 => n291, SL => 
                           mult_21_C249_n1539, Z => mult_21_C249_n987);
   mult_21_C249_U961 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n987, Z => 
                           mult_21_C249_n1290);
   mult_21_C249_U960 : MUXB2DL port map( A0 => n289, A1 => n292, SL => 
                           mult_21_C249_n1539, Z => mult_21_C249_n986);
   mult_21_C249_U959 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n986, Z => 
                           mult_21_C249_n1289);
   mult_21_C249_U958 : MUXB2DL port map( A0 => n290, A1 => n289, SL => 
                           mult_21_C249_n1539, Z => mult_21_C249_n985);
   mult_21_C249_U957 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n985, Z => 
                           mult_21_C249_n1288);
   mult_21_C249_U956 : MUXB2DL port map( A0 => n293, A1 => n290, SL => 
                           mult_21_C249_n1539, Z => mult_21_C249_n984);
   mult_21_C249_U955 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n984, Z => 
                           mult_21_C249_n1287);
   mult_21_C249_U954 : MUXB2DL port map( A0 => n294, A1 => n293, SL => 
                           mult_21_C249_n1539, Z => mult_21_C249_n983);
   mult_21_C249_U953 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n983, Z => 
                           mult_21_C249_n1286);
   mult_21_C249_U952 : MUXB2DL port map( A0 => n295, A1 => n294, SL => 
                           mult_21_C249_n1539, Z => mult_21_C249_n982);
   mult_21_C249_U951 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n982, Z => 
                           mult_21_C249_n1285);
   mult_21_C249_U950 : MUXB2DL port map( A0 => n296, A1 => n295, SL => 
                           mult_21_C249_n1539, Z => mult_21_C249_n981);
   mult_21_C249_U949 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n981, Z => 
                           mult_21_C249_n1284);
   mult_21_C249_U948 : MUXB2DL port map( A0 => n297, A1 => n296, SL => 
                           mult_21_C249_n1539, Z => mult_21_C249_n980);
   mult_21_C249_U947 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n980, Z => 
                           mult_21_C249_n1283);
   mult_21_C249_U946 : MUXB2DL port map( A0 => n298, A1 => n297, SL => 
                           mult_21_C249_n1539, Z => mult_21_C249_n979);
   mult_21_C249_U945 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n979, Z => 
                           mult_21_C249_n1282);
   mult_21_C249_U944 : MUXB2DL port map( A0 => n299, A1 => n298, SL => 
                           mult_21_C249_n1539, Z => mult_21_C249_n978);
   mult_21_C249_U943 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n978, Z => 
                           mult_21_C249_n1281);
   mult_21_C249_U942 : MUXB2DL port map( A0 => n302, A1 => n299, SL => 
                           mult_21_C249_n1539, Z => mult_21_C249_n977);
   mult_21_C249_U941 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n977, Z => 
                           mult_21_C249_n1280);
   mult_21_C249_U940 : MUXB2DL port map( A0 => n303, A1 => n302, SL => 
                           mult_21_C249_n1539, Z => mult_21_C249_n976);
   mult_21_C249_U939 : MUXB2DL port map( A0 => mult_21_C249_n1520, A1 => 
                           mult_21_C249_n22, SL => mult_21_C249_n976, Z => 
                           mult_21_C249_n1279);
   mult_21_C249_U938 : NOR2M1D1 port map( A1 => mult_21_C249_n1520, A2 => 
                           mult_21_C249_n22, Z => mult_21_C249_n1094);
   mult_21_C249_U937 : NAN2M1D1 port map( A1 => mult_21_C249_n1517, A2 => 
                           mult_21_C249_n1556, Z => mult_21_C249_n975);
   mult_21_C249_U936 : MUXB2DL port map( A0 => mult_21_C249_n1538, A1 => 
                           mult_21_C249_n30, SL => mult_21_C249_n975, Z => 
                           mult_21_C249_n1278);
   mult_21_C249_U935 : MUXB2DL port map( A0 => mult_21_C249_n1553, A1 => 
                           mult_21_C249_n1556, SL => mult_21_C249_n1517, Z => 
                           mult_21_C249_n974);
   mult_21_C249_U934 : MUXB2DL port map( A0 => mult_21_C249_n1538, A1 => 
                           mult_21_C249_n30, SL => mult_21_C249_n974, Z => 
                           mult_21_C249_n1277);
   mult_21_C249_U933 : MUXB2DL port map( A0 => n284, A1 => mult_21_C249_n1554, 
                           SL => mult_21_C249_n1517, Z => mult_21_C249_n973);
   mult_21_C249_U932 : MUXB2DL port map( A0 => mult_21_C249_n1538, A1 => 
                           mult_21_C249_n30, SL => mult_21_C249_n973, Z => 
                           mult_21_C249_n1276);
   mult_21_C249_U931 : MUXB2DL port map( A0 => mult_21_C249_n1551, A1 => n284, 
                           SL => mult_21_C249_n1517, Z => mult_21_C249_n972);
   mult_21_C249_U930 : MUXB2DL port map( A0 => mult_21_C249_n1538, A1 => 
                           mult_21_C249_n30, SL => mult_21_C249_n972, Z => 
                           mult_21_C249_n1275);
   mult_21_C249_U929 : MUXB2DL port map( A0 => n287, A1 => mult_21_C249_n1551, 
                           SL => mult_21_C249_n1517, Z => mult_21_C249_n971);
   mult_21_C249_U928 : MUXB2DL port map( A0 => mult_21_C249_n1538, A1 => 
                           mult_21_C249_n30, SL => mult_21_C249_n971, Z => 
                           mult_21_C249_n1274);
   mult_21_C249_U927 : MUXB2DL port map( A0 => n282, A1 => mult_21_C249_n1549, 
                           SL => mult_21_C249_n1517, Z => mult_21_C249_n970);
   mult_21_C249_U926 : MUXB2DL port map( A0 => mult_21_C249_n1538, A1 => 
                           mult_21_C249_n30, SL => mult_21_C249_n970, Z => 
                           mult_21_C249_n1273);
   mult_21_C249_U925 : MUXB2DL port map( A0 => n278, A1 => mult_21_C249_n1547, 
                           SL => mult_21_C249_n1517, Z => mult_21_C249_n969);
   mult_21_C249_U924 : MUXB2DL port map( A0 => mult_21_C249_n1538, A1 => 
                           mult_21_C249_n30, SL => mult_21_C249_n969, Z => 
                           mult_21_C249_n1272);
   mult_21_C249_U923 : MUXB2DL port map( A0 => n279, A1 => mult_21_C249_n1545, 
                           SL => mult_21_C249_n1517, Z => mult_21_C249_n968);
   mult_21_C249_U922 : MUXB2DL port map( A0 => mult_21_C249_n1538, A1 => 
                           mult_21_C249_n30, SL => mult_21_C249_n968, Z => 
                           mult_21_C249_n1271);
   mult_21_C249_U921 : MUXB2DL port map( A0 => n280, A1 => mult_21_C249_n1543, 
                           SL => mult_21_C249_n1517, Z => mult_21_C249_n967);
   mult_21_C249_U920 : MUXB2DL port map( A0 => mult_21_C249_n1538, A1 => 
                           mult_21_C249_n30, SL => mult_21_C249_n967, Z => 
                           mult_21_C249_n1270);
   mult_21_C249_U919 : MUXB2DL port map( A0 => mult_21_C249_n1541, A1 => n280, 
                           SL => mult_21_C249_n1517, Z => mult_21_C249_n966);
   mult_21_C249_U918 : MUXB2DL port map( A0 => mult_21_C249_n1538, A1 => 
                           mult_21_C249_n30, SL => mult_21_C249_n966, Z => 
                           mult_21_C249_n1269);
   mult_21_C249_U917 : MUXB2DL port map( A0 => n285, A1 => mult_21_C249_n1541, 
                           SL => mult_21_C249_n1517, Z => mult_21_C249_n965);
   mult_21_C249_U916 : MUXB2DL port map( A0 => mult_21_C249_n1538, A1 => 
                           mult_21_C249_n30, SL => mult_21_C249_n965, Z => 
                           mult_21_C249_n1268);
   mult_21_C249_U915 : MUXB2DL port map( A0 => n274, A1 => n285, SL => 
                           mult_21_C249_n1517, Z => mult_21_C249_n964);
   mult_21_C249_U914 : MUXB2DL port map( A0 => mult_21_C249_n1538, A1 => 
                           mult_21_C249_n30, SL => mult_21_C249_n964, Z => 
                           mult_21_C249_n1267);
   mult_21_C249_U913 : MUXB2DL port map( A0 => n271, A1 => n274, SL => 
                           mult_21_C249_n1517, Z => mult_21_C249_n963);
   mult_21_C249_U912 : MUXB2DL port map( A0 => mult_21_C249_n1538, A1 => 
                           mult_21_C249_n30, SL => mult_21_C249_n963, Z => 
                           mult_21_C249_n1266);
   mult_21_C249_U911 : MUXB2DL port map( A0 => n272, A1 => n271, SL => 
                           mult_21_C249_n1517, Z => mult_21_C249_n962);
   mult_21_C249_U910 : MUXB2DL port map( A0 => mult_21_C249_n1538, A1 => 
                           mult_21_C249_n30, SL => mult_21_C249_n962, Z => 
                           mult_21_C249_n1265);
   mult_21_C249_U909 : MUXB2DL port map( A0 => n273, A1 => n272, SL => 
                           mult_21_C249_n1517, Z => mult_21_C249_n961);
   mult_21_C249_U908 : MUXB2DL port map( A0 => mult_21_C249_n1538, A1 => 
                           mult_21_C249_n30, SL => mult_21_C249_n961, Z => 
                           mult_21_C249_n1264);
   mult_21_C249_U907 : MUXB2DL port map( A0 => n291, A1 => n273, SL => 
                           mult_21_C249_n1517, Z => mult_21_C249_n960);
   mult_21_C249_U906 : MUXB2DL port map( A0 => mult_21_C249_n1538, A1 => 
                           mult_21_C249_n30, SL => mult_21_C249_n960, Z => 
                           mult_21_C249_n1263);
   mult_21_C249_U905 : MUXB2DL port map( A0 => n292, A1 => n291, SL => 
                           mult_21_C249_n1517, Z => mult_21_C249_n959);
   mult_21_C249_U904 : MUXB2DL port map( A0 => mult_21_C249_n1538, A1 => 
                           mult_21_C249_n30, SL => mult_21_C249_n959, Z => 
                           mult_21_C249_n1262);
   mult_21_C249_U903 : MUXB2DL port map( A0 => n289, A1 => n292, SL => 
                           mult_21_C249_n1517, Z => mult_21_C249_n958);
   mult_21_C249_U902 : MUXB2DL port map( A0 => mult_21_C249_n1538, A1 => 
                           mult_21_C249_n30, SL => mult_21_C249_n958, Z => 
                           mult_21_C249_n1261);
   mult_21_C249_U901 : MUXB2DL port map( A0 => n290, A1 => n289, SL => 
                           mult_21_C249_n1517, Z => mult_21_C249_n957);
   mult_21_C249_U900 : MUXB2DL port map( A0 => mult_21_C249_n1538, A1 => 
                           mult_21_C249_n30, SL => mult_21_C249_n957, Z => 
                           mult_21_C249_n1260);
   mult_21_C249_U899 : MUXB2DL port map( A0 => n293, A1 => n290, SL => 
                           mult_21_C249_n1517, Z => mult_21_C249_n956);
   mult_21_C249_U898 : MUXB2DL port map( A0 => mult_21_C249_n1538, A1 => 
                           mult_21_C249_n30, SL => mult_21_C249_n956, Z => 
                           mult_21_C249_n1259);
   mult_21_C249_U897 : MUXB2DL port map( A0 => n294, A1 => n293, SL => 
                           mult_21_C249_n1517, Z => mult_21_C249_n955);
   mult_21_C249_U896 : MUXB2DL port map( A0 => mult_21_C249_n1538, A1 => 
                           mult_21_C249_n30, SL => mult_21_C249_n955, Z => 
                           mult_21_C249_n1258);
   mult_21_C249_U895 : MUXB2DL port map( A0 => n295, A1 => n294, SL => 
                           mult_21_C249_n1517, Z => mult_21_C249_n954);
   mult_21_C249_U894 : MUXB2DL port map( A0 => mult_21_C249_n1538, A1 => 
                           mult_21_C249_n30, SL => mult_21_C249_n954, Z => 
                           mult_21_C249_n1257);
   mult_21_C249_U893 : MUXB2DL port map( A0 => n296, A1 => n295, SL => 
                           mult_21_C249_n1517, Z => mult_21_C249_n953);
   mult_21_C249_U892 : MUXB2DL port map( A0 => mult_21_C249_n1538, A1 => 
                           mult_21_C249_n30, SL => mult_21_C249_n953, Z => 
                           mult_21_C249_n1256);
   mult_21_C249_U891 : MUXB2DL port map( A0 => n297, A1 => n296, SL => 
                           mult_21_C249_n1517, Z => mult_21_C249_n952);
   mult_21_C249_U890 : MUXB2DL port map( A0 => mult_21_C249_n1538, A1 => 
                           mult_21_C249_n30, SL => mult_21_C249_n952, Z => 
                           mult_21_C249_n1255);
   mult_21_C249_U889 : MUXB2DL port map( A0 => n298, A1 => n297, SL => 
                           mult_21_C249_n1517, Z => mult_21_C249_n951);
   mult_21_C249_U888 : MUXB2DL port map( A0 => mult_21_C249_n1538, A1 => 
                           mult_21_C249_n30, SL => mult_21_C249_n951, Z => 
                           mult_21_C249_n1254);
   mult_21_C249_U887 : MUXB2DL port map( A0 => n299, A1 => n298, SL => 
                           mult_21_C249_n1517, Z => mult_21_C249_n950);
   mult_21_C249_U886 : MUXB2DL port map( A0 => mult_21_C249_n1538, A1 => 
                           mult_21_C249_n30, SL => mult_21_C249_n950, Z => 
                           mult_21_C249_n1253);
   mult_21_C249_U884 : NAN2M1D1 port map( A1 => mult_21_C249_n1518, A2 => 
                           mult_21_C249_n1556, Z => mult_21_C249_n949);
   mult_21_C249_U883 : MUXB2DL port map( A0 => mult_21_C249_n1521, A1 => 
                           mult_21_C249_n38, SL => mult_21_C249_n949, Z => 
                           mult_21_C249_n1252);
   mult_21_C249_U882 : MUXB2DL port map( A0 => mult_21_C249_n1553, A1 => 
                           mult_21_C249_n1556, SL => mult_21_C249_n1518, Z => 
                           mult_21_C249_n948);
   mult_21_C249_U881 : MUXB2DL port map( A0 => mult_21_C249_n1521, A1 => 
                           mult_21_C249_n38, SL => mult_21_C249_n948, Z => 
                           mult_21_C249_n1251);
   mult_21_C249_U880 : MUXB2DL port map( A0 => n284, A1 => mult_21_C249_n1554, 
                           SL => mult_21_C249_n1518, Z => mult_21_C249_n947);
   mult_21_C249_U879 : MUXB2DL port map( A0 => mult_21_C249_n1521, A1 => 
                           mult_21_C249_n38, SL => mult_21_C249_n947, Z => 
                           mult_21_C249_n1250);
   mult_21_C249_U878 : MUXB2DL port map( A0 => mult_21_C249_n1551, A1 => n284, 
                           SL => mult_21_C249_n1518, Z => mult_21_C249_n946);
   mult_21_C249_U877 : MUXB2DL port map( A0 => mult_21_C249_n1521, A1 => 
                           mult_21_C249_n38, SL => mult_21_C249_n946, Z => 
                           mult_21_C249_n1249);
   mult_21_C249_U876 : MUXB2DL port map( A0 => n287, A1 => mult_21_C249_n1551, 
                           SL => mult_21_C249_n1518, Z => mult_21_C249_n945);
   mult_21_C249_U875 : MUXB2DL port map( A0 => mult_21_C249_n1521, A1 => 
                           mult_21_C249_n38, SL => mult_21_C249_n945, Z => 
                           mult_21_C249_n1248);
   mult_21_C249_U874 : MUXB2DL port map( A0 => n282, A1 => mult_21_C249_n1549, 
                           SL => mult_21_C249_n1518, Z => mult_21_C249_n944);
   mult_21_C249_U873 : MUXB2DL port map( A0 => mult_21_C249_n1521, A1 => 
                           mult_21_C249_n38, SL => mult_21_C249_n944, Z => 
                           mult_21_C249_n1247);
   mult_21_C249_U872 : MUXB2DL port map( A0 => n278, A1 => mult_21_C249_n1547, 
                           SL => mult_21_C249_n1518, Z => mult_21_C249_n943);
   mult_21_C249_U871 : MUXB2DL port map( A0 => mult_21_C249_n1521, A1 => 
                           mult_21_C249_n38, SL => mult_21_C249_n943, Z => 
                           mult_21_C249_n1246);
   mult_21_C249_U870 : MUXB2DL port map( A0 => n279, A1 => mult_21_C249_n1545, 
                           SL => mult_21_C249_n1518, Z => mult_21_C249_n942);
   mult_21_C249_U869 : MUXB2DL port map( A0 => mult_21_C249_n1521, A1 => 
                           mult_21_C249_n38, SL => mult_21_C249_n942, Z => 
                           mult_21_C249_n1245);
   mult_21_C249_U868 : MUXB2DL port map( A0 => n280, A1 => mult_21_C249_n1543, 
                           SL => mult_21_C249_n1518, Z => mult_21_C249_n941);
   mult_21_C249_U867 : MUXB2DL port map( A0 => mult_21_C249_n1521, A1 => 
                           mult_21_C249_n38, SL => mult_21_C249_n941, Z => 
                           mult_21_C249_n1244);
   mult_21_C249_U866 : MUXB2DL port map( A0 => mult_21_C249_n1541, A1 => n280, 
                           SL => mult_21_C249_n1518, Z => mult_21_C249_n940);
   mult_21_C249_U865 : MUXB2DL port map( A0 => mult_21_C249_n1521, A1 => 
                           mult_21_C249_n38, SL => mult_21_C249_n940, Z => 
                           mult_21_C249_n1243);
   mult_21_C249_U864 : MUXB2DL port map( A0 => n285, A1 => mult_21_C249_n1541, 
                           SL => mult_21_C249_n1518, Z => mult_21_C249_n939);
   mult_21_C249_U863 : MUXB2DL port map( A0 => mult_21_C249_n1521, A1 => 
                           mult_21_C249_n38, SL => mult_21_C249_n939, Z => 
                           mult_21_C249_n1242);
   mult_21_C249_U862 : MUXB2DL port map( A0 => n274, A1 => n285, SL => 
                           mult_21_C249_n1518, Z => mult_21_C249_n938);
   mult_21_C249_U861 : MUXB2DL port map( A0 => mult_21_C249_n1521, A1 => 
                           mult_21_C249_n38, SL => mult_21_C249_n938, Z => 
                           mult_21_C249_n1241);
   mult_21_C249_U860 : MUXB2DL port map( A0 => n271, A1 => n274, SL => 
                           mult_21_C249_n1518, Z => mult_21_C249_n937);
   mult_21_C249_U859 : MUXB2DL port map( A0 => mult_21_C249_n1521, A1 => 
                           mult_21_C249_n38, SL => mult_21_C249_n937, Z => 
                           mult_21_C249_n1240);
   mult_21_C249_U858 : MUXB2DL port map( A0 => n272, A1 => n271, SL => 
                           mult_21_C249_n1518, Z => mult_21_C249_n936);
   mult_21_C249_U857 : MUXB2DL port map( A0 => mult_21_C249_n1521, A1 => 
                           mult_21_C249_n38, SL => mult_21_C249_n936, Z => 
                           mult_21_C249_n1239);
   mult_21_C249_U856 : MUXB2DL port map( A0 => n273, A1 => n272, SL => 
                           mult_21_C249_n1518, Z => mult_21_C249_n935);
   mult_21_C249_U855 : MUXB2DL port map( A0 => mult_21_C249_n1521, A1 => 
                           mult_21_C249_n38, SL => mult_21_C249_n935, Z => 
                           mult_21_C249_n1238);
   mult_21_C249_U854 : MUXB2DL port map( A0 => n291, A1 => n273, SL => 
                           mult_21_C249_n1518, Z => mult_21_C249_n934);
   mult_21_C249_U853 : MUXB2DL port map( A0 => mult_21_C249_n1521, A1 => 
                           mult_21_C249_n38, SL => mult_21_C249_n934, Z => 
                           mult_21_C249_n1237);
   mult_21_C249_U852 : MUXB2DL port map( A0 => n292, A1 => n291, SL => 
                           mult_21_C249_n1518, Z => mult_21_C249_n933);
   mult_21_C249_U851 : MUXB2DL port map( A0 => mult_21_C249_n1521, A1 => 
                           mult_21_C249_n38, SL => mult_21_C249_n933, Z => 
                           mult_21_C249_n1236);
   mult_21_C249_U850 : MUXB2DL port map( A0 => n289, A1 => n292, SL => 
                           mult_21_C249_n1518, Z => mult_21_C249_n932);
   mult_21_C249_U849 : MUXB2DL port map( A0 => mult_21_C249_n1521, A1 => 
                           mult_21_C249_n38, SL => mult_21_C249_n932, Z => 
                           mult_21_C249_n1235);
   mult_21_C249_U848 : MUXB2DL port map( A0 => n290, A1 => n289, SL => 
                           mult_21_C249_n1518, Z => mult_21_C249_n931);
   mult_21_C249_U847 : MUXB2DL port map( A0 => mult_21_C249_n1521, A1 => 
                           mult_21_C249_n38, SL => mult_21_C249_n931, Z => 
                           mult_21_C249_n1234);
   mult_21_C249_U846 : MUXB2DL port map( A0 => n293, A1 => n290, SL => 
                           mult_21_C249_n1518, Z => mult_21_C249_n930);
   mult_21_C249_U845 : MUXB2DL port map( A0 => mult_21_C249_n1521, A1 => 
                           mult_21_C249_n38, SL => mult_21_C249_n930, Z => 
                           mult_21_C249_n1233);
   mult_21_C249_U844 : MUXB2DL port map( A0 => n294, A1 => n293, SL => 
                           mult_21_C249_n1518, Z => mult_21_C249_n929);
   mult_21_C249_U843 : MUXB2DL port map( A0 => mult_21_C249_n1521, A1 => 
                           mult_21_C249_n38, SL => mult_21_C249_n929, Z => 
                           mult_21_C249_n1232);
   mult_21_C249_U842 : MUXB2DL port map( A0 => n295, A1 => n294, SL => 
                           mult_21_C249_n1518, Z => mult_21_C249_n928);
   mult_21_C249_U841 : MUXB2DL port map( A0 => mult_21_C249_n1521, A1 => 
                           mult_21_C249_n38, SL => mult_21_C249_n928, Z => 
                           mult_21_C249_n1231);
   mult_21_C249_U840 : MUXB2DL port map( A0 => n296, A1 => n295, SL => 
                           mult_21_C249_n1518, Z => mult_21_C249_n927);
   mult_21_C249_U839 : MUXB2DL port map( A0 => mult_21_C249_n1521, A1 => 
                           mult_21_C249_n38, SL => mult_21_C249_n927, Z => 
                           mult_21_C249_n1230);
   mult_21_C249_U838 : MUXB2DL port map( A0 => n297, A1 => n296, SL => 
                           mult_21_C249_n1518, Z => mult_21_C249_n926);
   mult_21_C249_U837 : MUXB2DL port map( A0 => mult_21_C249_n1521, A1 => 
                           mult_21_C249_n38, SL => mult_21_C249_n926, Z => 
                           mult_21_C249_n1229);
   mult_21_C249_U836 : NOR2M1D1 port map( A1 => mult_21_C249_n1521, A2 => 
                           mult_21_C249_n38, Z => mult_21_C249_n1092);
   mult_21_C249_U835 : NAN2M1D1 port map( A1 => mult_21_C249_n48, A2 => 
                           mult_21_C249_n1556, Z => mult_21_C249_n925);
   mult_21_C249_U834 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n45, SL => mult_21_C249_n925, Z => 
                           mult_21_C249_n1228);
   mult_21_C249_U833 : MUXB2DL port map( A0 => mult_21_C249_n1554, A1 => 
                           mult_21_C249_n1556, SL => mult_21_C249_n48, Z => 
                           mult_21_C249_n924);
   mult_21_C249_U832 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n45, SL => mult_21_C249_n924, Z => 
                           mult_21_C249_n1227);
   mult_21_C249_U831 : MUXB2DL port map( A0 => n284, A1 => mult_21_C249_n1554, 
                           SL => mult_21_C249_n48, Z => mult_21_C249_n923);
   mult_21_C249_U830 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n45, SL => mult_21_C249_n923, Z => 
                           mult_21_C249_n1226);
   mult_21_C249_U829 : MUXB2DL port map( A0 => mult_21_C249_n1551, A1 => n284, 
                           SL => mult_21_C249_n48, Z => mult_21_C249_n922);
   mult_21_C249_U828 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n45, SL => mult_21_C249_n922, Z => 
                           mult_21_C249_n1225);
   mult_21_C249_U827 : MUXB2DL port map( A0 => n287, A1 => mult_21_C249_n1551, 
                           SL => mult_21_C249_n48, Z => mult_21_C249_n921);
   mult_21_C249_U826 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n45, SL => mult_21_C249_n921, Z => 
                           mult_21_C249_n1224);
   mult_21_C249_U825 : MUXB2DL port map( A0 => mult_21_C249_n1547, A1 => n287, 
                           SL => mult_21_C249_n48, Z => mult_21_C249_n920);
   mult_21_C249_U824 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n45, SL => mult_21_C249_n920, Z => 
                           mult_21_C249_n1223);
   mult_21_C249_U823 : MUXB2DL port map( A0 => mult_21_C249_n1545, A1 => 
                           mult_21_C249_n1547, SL => mult_21_C249_n48, Z => 
                           mult_21_C249_n919);
   mult_21_C249_U822 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n45, SL => mult_21_C249_n919, Z => 
                           mult_21_C249_n1222);
   mult_21_C249_U821 : MUXB2DL port map( A0 => n279, A1 => mult_21_C249_n1545, 
                           SL => mult_21_C249_n48, Z => mult_21_C249_n918);
   mult_21_C249_U820 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n45, SL => mult_21_C249_n918, Z => 
                           mult_21_C249_n1221);
   mult_21_C249_U819 : MUXB2DL port map( A0 => n280, A1 => mult_21_C249_n1543, 
                           SL => mult_21_C249_n48, Z => mult_21_C249_n917);
   mult_21_C249_U818 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n45, SL => mult_21_C249_n917, Z => 
                           mult_21_C249_n1220);
   mult_21_C249_U817 : MUXB2DL port map( A0 => mult_21_C249_n1541, A1 => n280, 
                           SL => mult_21_C249_n48, Z => mult_21_C249_n916);
   mult_21_C249_U816 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n45, SL => mult_21_C249_n916, Z => 
                           mult_21_C249_n1219);
   mult_21_C249_U815 : MUXB2DL port map( A0 => n285, A1 => n281, SL => 
                           mult_21_C249_n48, Z => mult_21_C249_n915);
   mult_21_C249_U814 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n45, SL => mult_21_C249_n915, Z => 
                           mult_21_C249_n1218);
   mult_21_C249_U813 : MUXB2DL port map( A0 => n274, A1 => n285, SL => 
                           mult_21_C249_n48, Z => mult_21_C249_n914);
   mult_21_C249_U812 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n45, SL => mult_21_C249_n914, Z => 
                           mult_21_C249_n1217);
   mult_21_C249_U811 : MUXB2DL port map( A0 => n271, A1 => n274, SL => 
                           mult_21_C249_n48, Z => mult_21_C249_n913);
   mult_21_C249_U810 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n45, SL => mult_21_C249_n913, Z => 
                           mult_21_C249_n1216);
   mult_21_C249_U809 : MUXB2DL port map( A0 => n272, A1 => n271, SL => 
                           mult_21_C249_n48, Z => mult_21_C249_n912);
   mult_21_C249_U808 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n45, SL => mult_21_C249_n912, Z => 
                           mult_21_C249_n1215);
   mult_21_C249_U807 : MUXB2DL port map( A0 => n273, A1 => n272, SL => 
                           mult_21_C249_n48, Z => mult_21_C249_n911);
   mult_21_C249_U806 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n45, SL => mult_21_C249_n911, Z => 
                           mult_21_C249_n1214);
   mult_21_C249_U805 : MUXB2DL port map( A0 => n291, A1 => n273, SL => 
                           mult_21_C249_n48, Z => mult_21_C249_n910);
   mult_21_C249_U804 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n45, SL => mult_21_C249_n910, Z => 
                           mult_21_C249_n1213);
   mult_21_C249_U803 : MUXB2DL port map( A0 => n292, A1 => n291, SL => 
                           mult_21_C249_n48, Z => mult_21_C249_n909);
   mult_21_C249_U802 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n45, SL => mult_21_C249_n909, Z => 
                           mult_21_C249_n1212);
   mult_21_C249_U801 : MUXB2DL port map( A0 => n289, A1 => n292, SL => 
                           mult_21_C249_n48, Z => mult_21_C249_n908);
   mult_21_C249_U800 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n45, SL => mult_21_C249_n908, Z => 
                           mult_21_C249_n1211);
   mult_21_C249_U799 : MUXB2DL port map( A0 => n290, A1 => n289, SL => 
                           mult_21_C249_n48, Z => mult_21_C249_n907);
   mult_21_C249_U798 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n45, SL => mult_21_C249_n907, Z => 
                           mult_21_C249_n1210);
   mult_21_C249_U797 : MUXB2DL port map( A0 => n293, A1 => n290, SL => 
                           mult_21_C249_n48, Z => mult_21_C249_n906);
   mult_21_C249_U796 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n45, SL => mult_21_C249_n906, Z => 
                           mult_21_C249_n1209);
   mult_21_C249_U795 : MUXB2DL port map( A0 => n294, A1 => n293, SL => 
                           mult_21_C249_n48, Z => mult_21_C249_n905);
   mult_21_C249_U794 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n45, SL => mult_21_C249_n905, Z => 
                           mult_21_C249_n1208);
   mult_21_C249_U793 : MUXB2DL port map( A0 => n295, A1 => n294, SL => 
                           mult_21_C249_n48, Z => mult_21_C249_n904);
   mult_21_C249_U792 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n45, SL => mult_21_C249_n904, Z => 
                           mult_21_C249_n1207);
   mult_21_C249_U791 : NOR2M1D1 port map( A1 => mult_21_C249_n42, A2 => 
                           mult_21_C249_n45, Z => mult_21_C249_n1091);
   mult_21_C249_U790 : NAN2M1D1 port map( A1 => mult_21_C249_n56, A2 => 
                           mult_21_C249_n1556, Z => mult_21_C249_n903);
   mult_21_C249_U789 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n53, SL => mult_21_C249_n903, Z => 
                           mult_21_C249_n1206);
   mult_21_C249_U788 : MUXB2DL port map( A0 => mult_21_C249_n1554, A1 => 
                           mult_21_C249_n1556, SL => mult_21_C249_n56, Z => 
                           mult_21_C249_n902);
   mult_21_C249_U787 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n53, SL => mult_21_C249_n902, Z => 
                           mult_21_C249_n1205);
   mult_21_C249_U786 : MUXB2DL port map( A0 => n284, A1 => mult_21_C249_n1554, 
                           SL => mult_21_C249_n56, Z => mult_21_C249_n901);
   mult_21_C249_U785 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n53, SL => mult_21_C249_n901, Z => 
                           mult_21_C249_n1204);
   mult_21_C249_U784 : MUXB2DL port map( A0 => mult_21_C249_n1551, A1 => n284, 
                           SL => mult_21_C249_n56, Z => mult_21_C249_n900);
   mult_21_C249_U783 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n53, SL => mult_21_C249_n900, Z => 
                           mult_21_C249_n1203);
   mult_21_C249_U782 : MUXB2DL port map( A0 => mult_21_C249_n1549, A1 => 
                           mult_21_C249_n1551, SL => mult_21_C249_n56, Z => 
                           mult_21_C249_n899);
   mult_21_C249_U781 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n53, SL => mult_21_C249_n899, Z => 
                           mult_21_C249_n1202);
   mult_21_C249_U780 : MUXB2DL port map( A0 => n282, A1 => n287, SL => 
                           mult_21_C249_n56, Z => mult_21_C249_n898);
   mult_21_C249_U779 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n53, SL => mult_21_C249_n898, Z => 
                           mult_21_C249_n1201);
   mult_21_C249_U778 : MUXB2DL port map( A0 => mult_21_C249_n1545, A1 => 
                           mult_21_C249_n1547, SL => mult_21_C249_n56, Z => 
                           mult_21_C249_n897);
   mult_21_C249_U777 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n53, SL => mult_21_C249_n897, Z => 
                           mult_21_C249_n1200);
   mult_21_C249_U776 : MUXB2DL port map( A0 => mult_21_C249_n1543, A1 => 
                           mult_21_C249_n1545, SL => mult_21_C249_n56, Z => 
                           mult_21_C249_n896);
   mult_21_C249_U775 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n53, SL => mult_21_C249_n896, Z => 
                           mult_21_C249_n1199);
   mult_21_C249_U774 : MUXB2DL port map( A0 => n280, A1 => mult_21_C249_n1543, 
                           SL => mult_21_C249_n56, Z => mult_21_C249_n895);
   mult_21_C249_U773 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n53, SL => mult_21_C249_n895, Z => 
                           mult_21_C249_n1198);
   mult_21_C249_U772 : MUXB2DL port map( A0 => mult_21_C249_n1541, A1 => n280, 
                           SL => mult_21_C249_n56, Z => mult_21_C249_n894);
   mult_21_C249_U771 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n53, SL => mult_21_C249_n894, Z => 
                           mult_21_C249_n1197);
   mult_21_C249_U770 : MUXB2DL port map( A0 => n285, A1 => n281, SL => 
                           mult_21_C249_n56, Z => mult_21_C249_n893);
   mult_21_C249_U769 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n53, SL => mult_21_C249_n893, Z => 
                           mult_21_C249_n1196);
   mult_21_C249_U768 : MUXB2DL port map( A0 => n274, A1 => n285, SL => 
                           mult_21_C249_n56, Z => mult_21_C249_n892);
   mult_21_C249_U767 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n53, SL => mult_21_C249_n892, Z => 
                           mult_21_C249_n1195);
   mult_21_C249_U766 : MUXB2DL port map( A0 => n271, A1 => n274, SL => 
                           mult_21_C249_n56, Z => mult_21_C249_n891);
   mult_21_C249_U765 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n53, SL => mult_21_C249_n891, Z => 
                           mult_21_C249_n1194);
   mult_21_C249_U764 : MUXB2DL port map( A0 => n272, A1 => n271, SL => 
                           mult_21_C249_n56, Z => mult_21_C249_n890);
   mult_21_C249_U763 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n53, SL => mult_21_C249_n890, Z => 
                           mult_21_C249_n1193);
   mult_21_C249_U762 : MUXB2DL port map( A0 => n273, A1 => n272, SL => 
                           mult_21_C249_n56, Z => mult_21_C249_n889);
   mult_21_C249_U761 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n53, SL => mult_21_C249_n889, Z => 
                           mult_21_C249_n1192);
   mult_21_C249_U760 : MUXB2DL port map( A0 => n291, A1 => n273, SL => 
                           mult_21_C249_n56, Z => mult_21_C249_n888);
   mult_21_C249_U759 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n53, SL => mult_21_C249_n888, Z => 
                           mult_21_C249_n1191);
   mult_21_C249_U758 : MUXB2DL port map( A0 => n292, A1 => n291, SL => 
                           mult_21_C249_n56, Z => mult_21_C249_n887);
   mult_21_C249_U757 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n53, SL => mult_21_C249_n887, Z => 
                           mult_21_C249_n1190);
   mult_21_C249_U756 : MUXB2DL port map( A0 => n289, A1 => n292, SL => 
                           mult_21_C249_n56, Z => mult_21_C249_n886);
   mult_21_C249_U755 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n53, SL => mult_21_C249_n886, Z => 
                           mult_21_C249_n1189);
   mult_21_C249_U754 : MUXB2DL port map( A0 => n290, A1 => n289, SL => 
                           mult_21_C249_n56, Z => mult_21_C249_n885);
   mult_21_C249_U753 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n53, SL => mult_21_C249_n885, Z => 
                           mult_21_C249_n1188);
   mult_21_C249_U752 : MUXB2DL port map( A0 => n293, A1 => n290, SL => 
                           mult_21_C249_n56, Z => mult_21_C249_n884);
   mult_21_C249_U751 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n53, SL => mult_21_C249_n884, Z => 
                           mult_21_C249_n1187);
   mult_21_C249_U750 : NOR2M1D1 port map( A1 => mult_21_C249_n50, A2 => 
                           mult_21_C249_n53, Z => mult_21_C249_n1090);
   mult_21_C249_U749 : NAN2M1D1 port map( A1 => mult_21_C249_n63, A2 => 
                           mult_21_C249_n1556, Z => mult_21_C249_n883);
   mult_21_C249_U748 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n61, SL => mult_21_C249_n883, Z => 
                           mult_21_C249_n1186);
   mult_21_C249_U747 : MUXB2DL port map( A0 => mult_21_C249_n1554, A1 => n288, 
                           SL => mult_21_C249_n63, Z => mult_21_C249_n882);
   mult_21_C249_U746 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n61, SL => mult_21_C249_n882, Z => 
                           mult_21_C249_n1185);
   mult_21_C249_U745 : MUXB2DL port map( A0 => n284, A1 => mult_21_C249_n1554, 
                           SL => mult_21_C249_n63, Z => mult_21_C249_n881);
   mult_21_C249_U744 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n61, SL => mult_21_C249_n881, Z => 
                           mult_21_C249_n1184);
   mult_21_C249_U743 : MUXB2DL port map( A0 => mult_21_C249_n1551, A1 => n284, 
                           SL => mult_21_C249_n63, Z => mult_21_C249_n880);
   mult_21_C249_U742 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n61, SL => mult_21_C249_n880, Z => 
                           mult_21_C249_n1183);
   mult_21_C249_U741 : MUXB2DL port map( A0 => mult_21_C249_n1549, A1 => n286, 
                           SL => mult_21_C249_n63, Z => mult_21_C249_n879);
   mult_21_C249_U740 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n61, SL => mult_21_C249_n879, Z => 
                           mult_21_C249_n1182);
   mult_21_C249_U739 : MUXB2DL port map( A0 => mult_21_C249_n1547, A1 => 
                           mult_21_C249_n1549, SL => mult_21_C249_n63, Z => 
                           mult_21_C249_n878);
   mult_21_C249_U738 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n61, SL => mult_21_C249_n878, Z => 
                           mult_21_C249_n1181);
   mult_21_C249_U737 : MUXB2DL port map( A0 => n278, A1 => n282, SL => 
                           mult_21_C249_n63, Z => mult_21_C249_n877);
   mult_21_C249_U736 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n61, SL => mult_21_C249_n877, Z => 
                           mult_21_C249_n1180);
   mult_21_C249_U735 : MUXB2DL port map( A0 => n279, A1 => mult_21_C249_n1545, 
                           SL => mult_21_C249_n63, Z => mult_21_C249_n876);
   mult_21_C249_U734 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n61, SL => mult_21_C249_n876, Z => 
                           mult_21_C249_n1179);
   mult_21_C249_U733 : MUXB2DL port map( A0 => n280, A1 => mult_21_C249_n1543, 
                           SL => mult_21_C249_n63, Z => mult_21_C249_n875);
   mult_21_C249_U732 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n61, SL => mult_21_C249_n875, Z => 
                           mult_21_C249_n1178);
   mult_21_C249_U731 : MUXB2DL port map( A0 => mult_21_C249_n1541, A1 => n280, 
                           SL => mult_21_C249_n63, Z => mult_21_C249_n874);
   mult_21_C249_U730 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n61, SL => mult_21_C249_n874, Z => 
                           mult_21_C249_n1177);
   mult_21_C249_U729 : MUXB2DL port map( A0 => n285, A1 => n281, SL => 
                           mult_21_C249_n63, Z => mult_21_C249_n873);
   mult_21_C249_U728 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n61, SL => mult_21_C249_n873, Z => 
                           mult_21_C249_n1176);
   mult_21_C249_U727 : MUXB2DL port map( A0 => n274, A1 => n285, SL => 
                           mult_21_C249_n63, Z => mult_21_C249_n872);
   mult_21_C249_U726 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n61, SL => mult_21_C249_n872, Z => 
                           mult_21_C249_n1175);
   mult_21_C249_U725 : MUXB2DL port map( A0 => n271, A1 => n274, SL => 
                           mult_21_C249_n63, Z => mult_21_C249_n871);
   mult_21_C249_U724 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n61, SL => mult_21_C249_n871, Z => 
                           mult_21_C249_n1174);
   mult_21_C249_U723 : MUXB2DL port map( A0 => n272, A1 => n271, SL => 
                           mult_21_C249_n63, Z => mult_21_C249_n870);
   mult_21_C249_U722 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n61, SL => mult_21_C249_n870, Z => 
                           mult_21_C249_n1173);
   mult_21_C249_U721 : MUXB2DL port map( A0 => n273, A1 => n272, SL => 
                           mult_21_C249_n63, Z => mult_21_C249_n869);
   mult_21_C249_U720 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n61, SL => mult_21_C249_n869, Z => 
                           mult_21_C249_n1172);
   mult_21_C249_U719 : MUXB2DL port map( A0 => n291, A1 => n273, SL => 
                           mult_21_C249_n63, Z => mult_21_C249_n868);
   mult_21_C249_U718 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n61, SL => mult_21_C249_n868, Z => 
                           mult_21_C249_n1171);
   mult_21_C249_U717 : MUXB2DL port map( A0 => n292, A1 => n291, SL => 
                           mult_21_C249_n63, Z => mult_21_C249_n867);
   mult_21_C249_U716 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n61, SL => mult_21_C249_n867, Z => 
                           mult_21_C249_n1170);
   mult_21_C249_U715 : MUXB2DL port map( A0 => n289, A1 => n292, SL => 
                           mult_21_C249_n63, Z => mult_21_C249_n866);
   mult_21_C249_U714 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n61, SL => mult_21_C249_n866, Z => 
                           mult_21_C249_n1169);
   mult_21_C249_U713 : NOR2M1D1 port map( A1 => mult_21_C249_n58, A2 => 
                           mult_21_C249_n61, Z => mult_21_C249_n1089);
   mult_21_C249_U712 : NAN2M1D1 port map( A1 => mult_21_C249_n71, A2 => 
                           mult_21_C249_n1556, Z => mult_21_C249_n865);
   mult_21_C249_U711 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n69, SL => mult_21_C249_n865, Z => 
                           mult_21_C249_n1168);
   mult_21_C249_U710 : MUXB2DL port map( A0 => mult_21_C249_n1553, A1 => n288, 
                           SL => mult_21_C249_n71, Z => mult_21_C249_n864);
   mult_21_C249_U709 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n69, SL => mult_21_C249_n864, Z => 
                           mult_21_C249_n1167);
   mult_21_C249_U708 : MUXB2DL port map( A0 => n284, A1 => mult_21_C249_n1554, 
                           SL => mult_21_C249_n71, Z => mult_21_C249_n863);
   mult_21_C249_U707 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n69, SL => mult_21_C249_n863, Z => 
                           mult_21_C249_n1166);
   mult_21_C249_U706 : MUXB2DL port map( A0 => mult_21_C249_n1551, A1 => n284, 
                           SL => mult_21_C249_n71, Z => mult_21_C249_n862);
   mult_21_C249_U705 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n69, SL => mult_21_C249_n862, Z => 
                           mult_21_C249_n1165);
   mult_21_C249_U704 : MUXB2DL port map( A0 => mult_21_C249_n1549, A1 => 
                           mult_21_C249_n1551, SL => mult_21_C249_n71, Z => 
                           mult_21_C249_n861);
   mult_21_C249_U703 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n69, SL => mult_21_C249_n861, Z => 
                           mult_21_C249_n1164);
   mult_21_C249_U702 : MUXB2DL port map( A0 => mult_21_C249_n1547, A1 => 
                           mult_21_C249_n1549, SL => mult_21_C249_n71, Z => 
                           mult_21_C249_n860);
   mult_21_C249_U701 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n69, SL => mult_21_C249_n860, Z => 
                           mult_21_C249_n1163);
   mult_21_C249_U700 : MUXB2DL port map( A0 => n278, A1 => mult_21_C249_n1547, 
                           SL => mult_21_C249_n71, Z => mult_21_C249_n859);
   mult_21_C249_U699 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n69, SL => mult_21_C249_n859, Z => 
                           mult_21_C249_n1162);
   mult_21_C249_U698 : MUXB2DL port map( A0 => n279, A1 => mult_21_C249_n1545, 
                           SL => mult_21_C249_n71, Z => mult_21_C249_n858);
   mult_21_C249_U697 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n69, SL => mult_21_C249_n858, Z => 
                           mult_21_C249_n1161);
   mult_21_C249_U696 : MUXB2DL port map( A0 => n280, A1 => mult_21_C249_n1543, 
                           SL => mult_21_C249_n71, Z => mult_21_C249_n857);
   mult_21_C249_U695 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n69, SL => mult_21_C249_n857, Z => 
                           mult_21_C249_n1160);
   mult_21_C249_U694 : MUXB2DL port map( A0 => mult_21_C249_n1541, A1 => n280, 
                           SL => mult_21_C249_n71, Z => mult_21_C249_n856);
   mult_21_C249_U693 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n69, SL => mult_21_C249_n856, Z => 
                           mult_21_C249_n1159);
   mult_21_C249_U692 : MUXB2DL port map( A0 => n285, A1 => n281, SL => 
                           mult_21_C249_n71, Z => mult_21_C249_n855);
   mult_21_C249_U691 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n69, SL => mult_21_C249_n855, Z => 
                           mult_21_C249_n1158);
   mult_21_C249_U690 : MUXB2DL port map( A0 => n274, A1 => n285, SL => 
                           mult_21_C249_n71, Z => mult_21_C249_n854);
   mult_21_C249_U689 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n69, SL => mult_21_C249_n854, Z => 
                           mult_21_C249_n1157);
   mult_21_C249_U688 : MUXB2DL port map( A0 => n271, A1 => n274, SL => 
                           mult_21_C249_n71, Z => mult_21_C249_n853);
   mult_21_C249_U687 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n69, SL => mult_21_C249_n853, Z => 
                           mult_21_C249_n1156);
   mult_21_C249_U686 : MUXB2DL port map( A0 => n272, A1 => n271, SL => 
                           mult_21_C249_n71, Z => mult_21_C249_n852);
   mult_21_C249_U685 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n69, SL => mult_21_C249_n852, Z => 
                           mult_21_C249_n1155);
   mult_21_C249_U684 : MUXB2DL port map( A0 => n273, A1 => n272, SL => 
                           mult_21_C249_n71, Z => mult_21_C249_n851);
   mult_21_C249_U683 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n69, SL => mult_21_C249_n851, Z => 
                           mult_21_C249_n1154);
   mult_21_C249_U682 : MUXB2DL port map( A0 => n291, A1 => n273, SL => 
                           mult_21_C249_n71, Z => mult_21_C249_n850);
   mult_21_C249_U681 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n69, SL => mult_21_C249_n850, Z => 
                           mult_21_C249_n1153);
   mult_21_C249_U680 : NOR2M1D1 port map( A1 => mult_21_C249_n66, A2 => 
                           mult_21_C249_n69, Z => mult_21_C249_n1088);
   mult_21_C249_U679 : NAN2M1D1 port map( A1 => mult_21_C249_n78, A2 => n288, Z
                           => mult_21_C249_n849);
   mult_21_C249_U678 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n76, SL => mult_21_C249_n849, Z => 
                           mult_21_C249_n1152);
   mult_21_C249_U677 : MUXB2DL port map( A0 => mult_21_C249_n1553, A1 => 
                           mult_21_C249_n1556, SL => mult_21_C249_n78, Z => 
                           mult_21_C249_n848);
   mult_21_C249_U676 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n76, SL => mult_21_C249_n848, Z => 
                           mult_21_C249_n1151);
   mult_21_C249_U675 : MUXB2DL port map( A0 => n284, A1 => mult_21_C249_n1554, 
                           SL => mult_21_C249_n78, Z => mult_21_C249_n847);
   mult_21_C249_U674 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n76, SL => mult_21_C249_n847, Z => 
                           mult_21_C249_n1150);
   mult_21_C249_U673 : MUXB2DL port map( A0 => n286, A1 => n284, SL => 
                           mult_21_C249_n78, Z => mult_21_C249_n846);
   mult_21_C249_U672 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n76, SL => mult_21_C249_n846, Z => 
                           mult_21_C249_n1149);
   mult_21_C249_U671 : MUXB2DL port map( A0 => n287, A1 => n286, SL => 
                           mult_21_C249_n78, Z => mult_21_C249_n845);
   mult_21_C249_U670 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n76, SL => mult_21_C249_n845, Z => 
                           mult_21_C249_n1148);
   mult_21_C249_U669 : MUXB2DL port map( A0 => n282, A1 => mult_21_C249_n1549, 
                           SL => mult_21_C249_n78, Z => mult_21_C249_n844);
   mult_21_C249_U668 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n76, SL => mult_21_C249_n844, Z => 
                           mult_21_C249_n1147);
   mult_21_C249_U667 : MUXB2DL port map( A0 => n278, A1 => mult_21_C249_n1547, 
                           SL => mult_21_C249_n78, Z => mult_21_C249_n843);
   mult_21_C249_U666 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n76, SL => mult_21_C249_n843, Z => 
                           mult_21_C249_n1146);
   mult_21_C249_U665 : MUXB2DL port map( A0 => n279, A1 => mult_21_C249_n1545, 
                           SL => mult_21_C249_n78, Z => mult_21_C249_n842);
   mult_21_C249_U664 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n76, SL => mult_21_C249_n842, Z => 
                           mult_21_C249_n1145);
   mult_21_C249_U663 : MUXB2DL port map( A0 => n280, A1 => mult_21_C249_n1543, 
                           SL => mult_21_C249_n78, Z => mult_21_C249_n841);
   mult_21_C249_U662 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n76, SL => mult_21_C249_n841, Z => 
                           mult_21_C249_n1144);
   mult_21_C249_U661 : MUXB2DL port map( A0 => mult_21_C249_n1541, A1 => n280, 
                           SL => mult_21_C249_n78, Z => mult_21_C249_n840);
   mult_21_C249_U660 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n76, SL => mult_21_C249_n840, Z => 
                           mult_21_C249_n1143);
   mult_21_C249_U659 : MUXB2DL port map( A0 => n285, A1 => n281, SL => 
                           mult_21_C249_n78, Z => mult_21_C249_n839);
   mult_21_C249_U658 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n76, SL => mult_21_C249_n839, Z => 
                           mult_21_C249_n1142);
   mult_21_C249_U657 : MUXB2DL port map( A0 => n274, A1 => n285, SL => 
                           mult_21_C249_n78, Z => mult_21_C249_n838);
   mult_21_C249_U656 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n76, SL => mult_21_C249_n838, Z => 
                           mult_21_C249_n1141);
   mult_21_C249_U655 : MUXB2DL port map( A0 => n271, A1 => n274, SL => 
                           mult_21_C249_n78, Z => mult_21_C249_n837);
   mult_21_C249_U654 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n76, SL => mult_21_C249_n837, Z => 
                           mult_21_C249_n1140);
   mult_21_C249_U653 : MUXB2DL port map( A0 => n272, A1 => n271, SL => 
                           mult_21_C249_n78, Z => mult_21_C249_n836);
   mult_21_C249_U652 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n76, SL => mult_21_C249_n836, Z => 
                           mult_21_C249_n1139);
   mult_21_C249_U651 : NOR2M1D1 port map( A1 => mult_21_C249_n73, A2 => 
                           mult_21_C249_n76, Z => mult_21_C249_n1087);
   mult_21_C249_U650 : NAN2M1D1 port map( A1 => mult_21_C249_n83, A2 => 
                           mult_21_C249_n1556, Z => mult_21_C249_n835);
   mult_21_C249_U649 : MUXB2DL port map( A0 => mult_21_C249_n79, A1 => 
                           mult_21_C249_n81, SL => mult_21_C249_n835, Z => 
                           mult_21_C249_n1138);
   mult_21_C249_U648 : MUXB2DL port map( A0 => mult_21_C249_n1553, A1 => n288, 
                           SL => mult_21_C249_n83, Z => mult_21_C249_n834);
   mult_21_C249_U647 : MUXB2DL port map( A0 => mult_21_C249_n79, A1 => 
                           mult_21_C249_n81, SL => mult_21_C249_n834, Z => 
                           mult_21_C249_n1137);
   mult_21_C249_U646 : MUXB2DL port map( A0 => n284, A1 => mult_21_C249_n1554, 
                           SL => mult_21_C249_n83, Z => mult_21_C249_n833);
   mult_21_C249_U645 : MUXB2DL port map( A0 => mult_21_C249_n79, A1 => 
                           mult_21_C249_n81, SL => mult_21_C249_n833, Z => 
                           mult_21_C249_n1136);
   mult_21_C249_U644 : MUXB2DL port map( A0 => n286, A1 => n284, SL => 
                           mult_21_C249_n83, Z => mult_21_C249_n832);
   mult_21_C249_U643 : MUXB2DL port map( A0 => mult_21_C249_n79, A1 => 
                           mult_21_C249_n81, SL => mult_21_C249_n832, Z => 
                           mult_21_C249_n1135);
   mult_21_C249_U642 : MUXB2DL port map( A0 => n287, A1 => n286, SL => 
                           mult_21_C249_n83, Z => mult_21_C249_n831);
   mult_21_C249_U641 : MUXB2DL port map( A0 => mult_21_C249_n79, A1 => 
                           mult_21_C249_n81, SL => mult_21_C249_n831, Z => 
                           mult_21_C249_n1134);
   mult_21_C249_U640 : MUXB2DL port map( A0 => n282, A1 => mult_21_C249_n1549, 
                           SL => mult_21_C249_n83, Z => mult_21_C249_n830);
   mult_21_C249_U639 : MUXB2DL port map( A0 => mult_21_C249_n79, A1 => 
                           mult_21_C249_n81, SL => mult_21_C249_n830, Z => 
                           mult_21_C249_n1133);
   mult_21_C249_U638 : MUXB2DL port map( A0 => n278, A1 => mult_21_C249_n1547, 
                           SL => mult_21_C249_n83, Z => mult_21_C249_n829);
   mult_21_C249_U637 : MUXB2DL port map( A0 => mult_21_C249_n79, A1 => 
                           mult_21_C249_n81, SL => mult_21_C249_n829, Z => 
                           mult_21_C249_n1132);
   mult_21_C249_U636 : MUXB2DL port map( A0 => n279, A1 => mult_21_C249_n1545, 
                           SL => mult_21_C249_n83, Z => mult_21_C249_n828);
   mult_21_C249_U635 : MUXB2DL port map( A0 => mult_21_C249_n79, A1 => 
                           mult_21_C249_n81, SL => mult_21_C249_n828, Z => 
                           mult_21_C249_n1131);
   mult_21_C249_U634 : MUXB2DL port map( A0 => n280, A1 => mult_21_C249_n1543, 
                           SL => mult_21_C249_n83, Z => mult_21_C249_n827);
   mult_21_C249_U633 : MUXB2DL port map( A0 => mult_21_C249_n79, A1 => 
                           mult_21_C249_n81, SL => mult_21_C249_n827, Z => 
                           mult_21_C249_n1130);
   mult_21_C249_U632 : MUXB2DL port map( A0 => mult_21_C249_n1541, A1 => n280, 
                           SL => mult_21_C249_n83, Z => mult_21_C249_n826);
   mult_21_C249_U631 : MUXB2DL port map( A0 => mult_21_C249_n79, A1 => 
                           mult_21_C249_n81, SL => mult_21_C249_n826, Z => 
                           mult_21_C249_n1129);
   mult_21_C249_U630 : MUXB2DL port map( A0 => n285, A1 => n281, SL => 
                           mult_21_C249_n83, Z => mult_21_C249_n825);
   mult_21_C249_U629 : MUXB2DL port map( A0 => mult_21_C249_n79, A1 => 
                           mult_21_C249_n81, SL => mult_21_C249_n825, Z => 
                           mult_21_C249_n1128);
   mult_21_C249_U628 : MUXB2DL port map( A0 => n274, A1 => n285, SL => 
                           mult_21_C249_n83, Z => mult_21_C249_n824);
   mult_21_C249_U627 : MUXB2DL port map( A0 => mult_21_C249_n79, A1 => 
                           mult_21_C249_n81, SL => mult_21_C249_n824, Z => 
                           mult_21_C249_n1127);
   mult_21_C249_U626 : NOR2M1D1 port map( A1 => mult_21_C249_n79, A2 => 
                           mult_21_C249_n81, Z => mult_21_C249_n1086);
   mult_21_C249_U625 : NAN2M1D1 port map( A1 => mult_21_C249_n88, A2 => n288, Z
                           => mult_21_C249_n823);
   mult_21_C249_U624 : MUXB2DL port map( A0 => mult_21_C249_n84, A1 => 
                           mult_21_C249_n86, SL => mult_21_C249_n823, Z => 
                           mult_21_C249_n1126);
   mult_21_C249_U623 : MUXB2DL port map( A0 => mult_21_C249_n1553, A1 => n288, 
                           SL => mult_21_C249_n88, Z => mult_21_C249_n822);
   mult_21_C249_U622 : MUXB2DL port map( A0 => mult_21_C249_n84, A1 => 
                           mult_21_C249_n86, SL => mult_21_C249_n822, Z => 
                           mult_21_C249_n1125);
   mult_21_C249_U621 : MUXB2DL port map( A0 => n284, A1 => mult_21_C249_n1554, 
                           SL => mult_21_C249_n88, Z => mult_21_C249_n821);
   mult_21_C249_U620 : MUXB2DL port map( A0 => mult_21_C249_n84, A1 => 
                           mult_21_C249_n86, SL => mult_21_C249_n821, Z => 
                           mult_21_C249_n1124);
   mult_21_C249_U619 : MUXB2DL port map( A0 => mult_21_C249_n1551, A1 => n284, 
                           SL => mult_21_C249_n88, Z => mult_21_C249_n820);
   mult_21_C249_U618 : MUXB2DL port map( A0 => mult_21_C249_n84, A1 => 
                           mult_21_C249_n86, SL => mult_21_C249_n820, Z => 
                           mult_21_C249_n1123);
   mult_21_C249_U617 : MUXB2DL port map( A0 => n287, A1 => n286, SL => 
                           mult_21_C249_n88, Z => mult_21_C249_n819);
   mult_21_C249_U616 : MUXB2DL port map( A0 => mult_21_C249_n84, A1 => 
                           mult_21_C249_n86, SL => mult_21_C249_n819, Z => 
                           mult_21_C249_n1122);
   mult_21_C249_U615 : MUXB2DL port map( A0 => n282, A1 => mult_21_C249_n1549, 
                           SL => mult_21_C249_n88, Z => mult_21_C249_n818);
   mult_21_C249_U614 : MUXB2DL port map( A0 => mult_21_C249_n84, A1 => 
                           mult_21_C249_n86, SL => mult_21_C249_n818, Z => 
                           mult_21_C249_n1121);
   mult_21_C249_U613 : MUXB2DL port map( A0 => n278, A1 => mult_21_C249_n1547, 
                           SL => mult_21_C249_n88, Z => mult_21_C249_n817);
   mult_21_C249_U612 : MUXB2DL port map( A0 => mult_21_C249_n84, A1 => 
                           mult_21_C249_n86, SL => mult_21_C249_n817, Z => 
                           mult_21_C249_n1120);
   mult_21_C249_U611 : MUXB2DL port map( A0 => n279, A1 => mult_21_C249_n1545, 
                           SL => mult_21_C249_n88, Z => mult_21_C249_n816);
   mult_21_C249_U610 : MUXB2DL port map( A0 => mult_21_C249_n84, A1 => 
                           mult_21_C249_n86, SL => mult_21_C249_n816, Z => 
                           mult_21_C249_n1119);
   mult_21_C249_U609 : MUXB2DL port map( A0 => n280, A1 => mult_21_C249_n1543, 
                           SL => mult_21_C249_n88, Z => mult_21_C249_n815);
   mult_21_C249_U608 : MUXB2DL port map( A0 => mult_21_C249_n84, A1 => 
                           mult_21_C249_n86, SL => mult_21_C249_n815, Z => 
                           mult_21_C249_n1118);
   mult_21_C249_U607 : MUXB2DL port map( A0 => mult_21_C249_n1541, A1 => n280, 
                           SL => mult_21_C249_n88, Z => mult_21_C249_n814);
   mult_21_C249_U606 : MUXB2DL port map( A0 => mult_21_C249_n84, A1 => 
                           mult_21_C249_n86, SL => mult_21_C249_n814, Z => 
                           mult_21_C249_n1117);
   mult_21_C249_U605 : NOR2M1D1 port map( A1 => mult_21_C249_n84, A2 => 
                           mult_21_C249_n86, Z => mult_21_C249_n1085);
   mult_21_C249_U604 : NAN2M1D1 port map( A1 => mult_21_C249_n93, A2 => n288, Z
                           => mult_21_C249_n813);
   mult_21_C249_U603 : MUXB2DL port map( A0 => mult_21_C249_n89, A1 => 
                           mult_21_C249_n91, SL => mult_21_C249_n813, Z => 
                           mult_21_C249_n1116);
   mult_21_C249_U602 : MUXB2DL port map( A0 => mult_21_C249_n1553, A1 => n288, 
                           SL => mult_21_C249_n93, Z => mult_21_C249_n812);
   mult_21_C249_U601 : MUXB2DL port map( A0 => mult_21_C249_n89, A1 => 
                           mult_21_C249_n91, SL => mult_21_C249_n812, Z => 
                           mult_21_C249_n1115);
   mult_21_C249_U600 : MUXB2DL port map( A0 => n284, A1 => mult_21_C249_n1553, 
                           SL => mult_21_C249_n93, Z => mult_21_C249_n811);
   mult_21_C249_U599 : MUXB2DL port map( A0 => mult_21_C249_n89, A1 => 
                           mult_21_C249_n91, SL => mult_21_C249_n811, Z => 
                           mult_21_C249_n1114);
   mult_21_C249_U598 : MUXB2DL port map( A0 => mult_21_C249_n1551, A1 => n284, 
                           SL => mult_21_C249_n93, Z => mult_21_C249_n810);
   mult_21_C249_U597 : MUXB2DL port map( A0 => mult_21_C249_n89, A1 => 
                           mult_21_C249_n91, SL => mult_21_C249_n810, Z => 
                           mult_21_C249_n1113);
   mult_21_C249_U596 : MUXB2DL port map( A0 => n287, A1 => n286, SL => 
                           mult_21_C249_n93, Z => mult_21_C249_n809);
   mult_21_C249_U595 : MUXB2DL port map( A0 => mult_21_C249_n89, A1 => 
                           mult_21_C249_n91, SL => mult_21_C249_n809, Z => 
                           mult_21_C249_n1112);
   mult_21_C249_U594 : MUXB2DL port map( A0 => n282, A1 => mult_21_C249_n1549, 
                           SL => mult_21_C249_n93, Z => mult_21_C249_n808);
   mult_21_C249_U593 : MUXB2DL port map( A0 => mult_21_C249_n89, A1 => 
                           mult_21_C249_n91, SL => mult_21_C249_n808, Z => 
                           mult_21_C249_n1111);
   mult_21_C249_U592 : MUXB2DL port map( A0 => n278, A1 => mult_21_C249_n1547, 
                           SL => mult_21_C249_n93, Z => mult_21_C249_n807);
   mult_21_C249_U591 : MUXB2DL port map( A0 => mult_21_C249_n89, A1 => 
                           mult_21_C249_n91, SL => mult_21_C249_n807, Z => 
                           mult_21_C249_n1110);
   mult_21_C249_U590 : MUXB2DL port map( A0 => n279, A1 => mult_21_C249_n1545, 
                           SL => mult_21_C249_n93, Z => mult_21_C249_n806);
   mult_21_C249_U589 : MUXB2DL port map( A0 => mult_21_C249_n89, A1 => 
                           mult_21_C249_n91, SL => mult_21_C249_n806, Z => 
                           mult_21_C249_n1109);
   mult_21_C249_U588 : NOR2M1D1 port map( A1 => mult_21_C249_n89, A2 => 
                           mult_21_C249_n91, Z => mult_21_C249_n1084);
   mult_21_C249_U587 : NAN2M1D1 port map( A1 => mult_21_C249_n98, A2 => 
                           mult_21_C249_n1556, Z => mult_21_C249_n805);
   mult_21_C249_U586 : MUXB2DL port map( A0 => mult_21_C249_n94, A1 => 
                           mult_21_C249_n96, SL => mult_21_C249_n805, Z => 
                           mult_21_C249_n1108);
   mult_21_C249_U585 : MUXB2DL port map( A0 => mult_21_C249_n1553, A1 => n288, 
                           SL => mult_21_C249_n98, Z => mult_21_C249_n804);
   mult_21_C249_U584 : MUXB2DL port map( A0 => mult_21_C249_n94, A1 => 
                           mult_21_C249_n96, SL => mult_21_C249_n804, Z => 
                           mult_21_C249_n1107);
   mult_21_C249_U583 : MUXB2DL port map( A0 => n284, A1 => mult_21_C249_n1554, 
                           SL => mult_21_C249_n98, Z => mult_21_C249_n803);
   mult_21_C249_U582 : MUXB2DL port map( A0 => mult_21_C249_n94, A1 => 
                           mult_21_C249_n96, SL => mult_21_C249_n803, Z => 
                           mult_21_C249_n1106);
   mult_21_C249_U581 : MUXB2DL port map( A0 => mult_21_C249_n1551, A1 => n284, 
                           SL => mult_21_C249_n98, Z => mult_21_C249_n802);
   mult_21_C249_U580 : MUXB2DL port map( A0 => mult_21_C249_n94, A1 => 
                           mult_21_C249_n96, SL => mult_21_C249_n802, Z => 
                           mult_21_C249_n1105);
   mult_21_C249_U579 : MUXB2DL port map( A0 => n287, A1 => n286, SL => 
                           mult_21_C249_n98, Z => mult_21_C249_n801);
   mult_21_C249_U578 : MUXB2DL port map( A0 => mult_21_C249_n94, A1 => 
                           mult_21_C249_n96, SL => mult_21_C249_n801, Z => 
                           mult_21_C249_n1104);
   mult_21_C249_U577 : MUXB2DL port map( A0 => n282, A1 => mult_21_C249_n1549, 
                           SL => mult_21_C249_n98, Z => mult_21_C249_n800);
   mult_21_C249_U576 : MUXB2DL port map( A0 => mult_21_C249_n94, A1 => 
                           mult_21_C249_n96, SL => mult_21_C249_n800, Z => 
                           mult_21_C249_n1103);
   mult_21_C249_U575 : NOR2M1D1 port map( A1 => mult_21_C249_n94, A2 => 
                           mult_21_C249_n96, Z => mult_21_C249_n1083);
   mult_21_C249_U574 : NAN2M1D1 port map( A1 => mult_21_C249_n103, A2 => 
                           mult_21_C249_n1556, Z => mult_21_C249_n799);
   mult_21_C249_U573 : MUXB2DL port map( A0 => mult_21_C249_n99, A1 => 
                           mult_21_C249_n101, SL => mult_21_C249_n799, Z => 
                           mult_21_C249_n1102);
   mult_21_C249_U572 : MUXB2DL port map( A0 => mult_21_C249_n1553, A1 => n288, 
                           SL => mult_21_C249_n103, Z => mult_21_C249_n798);
   mult_21_C249_U571 : MUXB2DL port map( A0 => mult_21_C249_n99, A1 => 
                           mult_21_C249_n101, SL => mult_21_C249_n798, Z => 
                           mult_21_C249_n1101);
   mult_21_C249_U570 : MUXB2DL port map( A0 => n284, A1 => mult_21_C249_n1553, 
                           SL => mult_21_C249_n103, Z => mult_21_C249_n797);
   mult_21_C249_U569 : MUXB2DL port map( A0 => mult_21_C249_n99, A1 => 
                           mult_21_C249_n101, SL => mult_21_C249_n797, Z => 
                           mult_21_C249_n1100);
   mult_21_C249_U568 : MUXB2DL port map( A0 => mult_21_C249_n1551, A1 => n284, 
                           SL => mult_21_C249_n103, Z => mult_21_C249_n796);
   mult_21_C249_U567 : MUXB2DL port map( A0 => mult_21_C249_n99, A1 => 
                           mult_21_C249_n101, SL => mult_21_C249_n796, Z => 
                           mult_21_C249_n1099);
   mult_21_C249_U566 : NOR2M1D1 port map( A1 => mult_21_C249_n99, A2 => 
                           mult_21_C249_n101, Z => mult_21_C249_n1082);
   mult_21_C249_U565 : NAN2M1D1 port map( A1 => mult_21_C249_n106, A2 => 
                           mult_21_C249_n1556, Z => mult_21_C249_n795);
   mult_21_C249_U564 : MUXB2DL port map( A0 => mult_21_C249_n104, A1 => 
                           mult_21_C249_n105, SL => mult_21_C249_n795, Z => 
                           mult_21_C249_n1098);
   mult_21_C249_U563 : MUXB2DL port map( A0 => mult_21_C249_n1553, A1 => n288, 
                           SL => mult_21_C249_n106, Z => mult_21_C249_n794);
   mult_21_C249_U562 : MUXB2DL port map( A0 => mult_21_C249_n104, A1 => 
                           mult_21_C249_n105, SL => mult_21_C249_n794, Z => 
                           mult_21_C249_n1097);
   mult_21_C249_U561 : NOR2M1D1 port map( A1 => mult_21_C249_n104, A2 => 
                           mult_21_C249_n105, Z => mult_21_C249_n1081);
   mult_21_C249_U557 : ADFULD1 port map( A => mult_21_C249_n1334, B => 
                           mult_21_C249_n1364, CI => mult_21_C249_n790, CO => 
                           mult_21_C249_n786, S => mult_21_C249_n787);
   mult_21_C249_U555 : ADFULD1 port map( A => mult_21_C249_n788, B => 
                           mult_21_C249_n1305, CI => mult_21_C249_n785, CO => 
                           mult_21_C249_n782, S => mult_21_C249_n783);
   mult_21_C249_U553 : ADFULD1 port map( A => mult_21_C249_n1304, B => 
                           mult_21_C249_n1362, CI => mult_21_C249_n1332, CO => 
                           mult_21_C249_n778, S => mult_21_C249_n779);
   mult_21_C249_U552 : ADFULD1 port map( A => mult_21_C249_n781, B => 
                           mult_21_C249_n784, CI => mult_21_C249_n779, CO => 
                           mult_21_C249_n776, S => mult_21_C249_n777);
   mult_21_C249_U550 : ADFULD1 port map( A => mult_21_C249_n1277, B => 
                           mult_21_C249_n1303, CI => mult_21_C249_n780, CO => 
                           mult_21_C249_n772, S => mult_21_C249_n773);
   mult_21_C249_U549 : ADFULD1 port map( A => mult_21_C249_n778, B => 
                           mult_21_C249_n775, CI => mult_21_C249_n773, CO => 
                           mult_21_C249_n770, S => mult_21_C249_n771);
   mult_21_C249_U547 : ADFULD1 port map( A => mult_21_C249_n1276, B => 
                           mult_21_C249_n1360, CI => mult_21_C249_n1330, CO => 
                           mult_21_C249_n766, S => mult_21_C249_n767);
   mult_21_C249_U546 : ADFULD1 port map( A => mult_21_C249_n774, B => 
                           mult_21_C249_n1302, CI => mult_21_C249_n769, CO => 
                           mult_21_C249_n764, S => mult_21_C249_n765);
   mult_21_C249_U545 : ADFULD1 port map( A => mult_21_C249_n767, B => 
                           mult_21_C249_n772, CI => mult_21_C249_n765, CO => 
                           mult_21_C249_n762, S => mult_21_C249_n763);
   mult_21_C249_U543 : ADFULD1 port map( A => mult_21_C249_n1275, B => 
                           mult_21_C249_n1301, CI => mult_21_C249_n1251, CO => 
                           mult_21_C249_n758, S => mult_21_C249_n759);
   mult_21_C249_U542 : ADFULD1 port map( A => mult_21_C249_n761, B => 
                           mult_21_C249_n768, CI => mult_21_C249_n766, CO => 
                           mult_21_C249_n756, S => mult_21_C249_n757);
   mult_21_C249_U541 : ADFULD1 port map( A => mult_21_C249_n764, B => 
                           mult_21_C249_n759, CI => mult_21_C249_n757, CO => 
                           mult_21_C249_n754, S => mult_21_C249_n755);
   mult_21_C249_U539 : ADFULD1 port map( A => mult_21_C249_n1250, B => 
                           mult_21_C249_n1358, CI => mult_21_C249_n1328, CO => 
                           mult_21_C249_n750, S => mult_21_C249_n751);
   mult_21_C249_U538 : ADFULD1 port map( A => mult_21_C249_n1274, B => 
                           mult_21_C249_n1300, CI => mult_21_C249_n760, CO => 
                           mult_21_C249_n748, S => mult_21_C249_n749);
   mult_21_C249_U537 : ADFULD1 port map( A => mult_21_C249_n758, B => 
                           mult_21_C249_n753, CI => mult_21_C249_n751, CO => 
                           mult_21_C249_n746, S => mult_21_C249_n747);
   mult_21_C249_U536 : ADFULD1 port map( A => mult_21_C249_n756, B => 
                           mult_21_C249_n749, CI => mult_21_C249_n747, CO => 
                           mult_21_C249_n744, S => mult_21_C249_n745);
   mult_21_C249_U534 : ADFULD1 port map( A => mult_21_C249_n1273, B => 
                           mult_21_C249_n1249, CI => mult_21_C249_n1227, CO => 
                           mult_21_C249_n740, S => mult_21_C249_n741);
   mult_21_C249_U533 : ADFULD1 port map( A => mult_21_C249_n752, B => 
                           mult_21_C249_n1299, CI => mult_21_C249_n743, CO => 
                           mult_21_C249_n738, S => mult_21_C249_n739);
   mult_21_C249_U532 : ADFULD1 port map( A => mult_21_C249_n748, B => 
                           mult_21_C249_n750, CI => mult_21_C249_n741, CO => 
                           mult_21_C249_n736, S => mult_21_C249_n737);
   mult_21_C249_U531 : ADFULD1 port map( A => mult_21_C249_n746, B => 
                           mult_21_C249_n739, CI => mult_21_C249_n737, CO => 
                           mult_21_C249_n734, S => mult_21_C249_n735);
   mult_21_C249_U529 : ADFULD1 port map( A => mult_21_C249_n1248, B => 
                           mult_21_C249_n1356, CI => mult_21_C249_n1326, CO => 
                           mult_21_C249_n730, S => mult_21_C249_n731);
   mult_21_C249_U528 : ADFULD1 port map( A => mult_21_C249_n1272, B => 
                           mult_21_C249_n1298, CI => mult_21_C249_n1226, CO => 
                           mult_21_C249_n728, S => mult_21_C249_n729);
   mult_21_C249_U527 : ADFULD1 port map( A => mult_21_C249_n733, B => 
                           mult_21_C249_n742, CI => mult_21_C249_n740, CO => 
                           mult_21_C249_n726, S => mult_21_C249_n727);
   mult_21_C249_U526 : ADFULD1 port map( A => mult_21_C249_n729, B => 
                           mult_21_C249_n731, CI => mult_21_C249_n738, CO => 
                           mult_21_C249_n724, S => mult_21_C249_n725);
   mult_21_C249_U525 : ADFULD1 port map( A => mult_21_C249_n736, B => 
                           mult_21_C249_n727, CI => mult_21_C249_n725, CO => 
                           mult_21_C249_n722, S => mult_21_C249_n723);
   mult_21_C249_U523 : ADFULD1 port map( A => mult_21_C249_n1205, B => 
                           mult_21_C249_n1297, CI => mult_21_C249_n1225, CO => 
                           mult_21_C249_n718, S => mult_21_C249_n719);
   mult_21_C249_U522 : ADFULD1 port map( A => mult_21_C249_n1247, B => 
                           mult_21_C249_n1271, CI => mult_21_C249_n732, CO => 
                           mult_21_C249_n716, S => mult_21_C249_n717);
   mult_21_C249_U521 : ADFULD1 port map( A => mult_21_C249_n730, B => 
                           mult_21_C249_n721, CI => mult_21_C249_n728, CO => 
                           mult_21_C249_n714, S => mult_21_C249_n715);
   mult_21_C249_U520 : ADFULD1 port map( A => mult_21_C249_n717, B => 
                           mult_21_C249_n719, CI => mult_21_C249_n726, CO => 
                           mult_21_C249_n712, S => mult_21_C249_n713);
   mult_21_C249_U519 : ADFULD1 port map( A => mult_21_C249_n724, B => 
                           mult_21_C249_n715, CI => mult_21_C249_n713, CO => 
                           mult_21_C249_n710, S => mult_21_C249_n711);
   mult_21_C249_U517 : ADFULD1 port map( A => mult_21_C249_n1204, B => 
                           mult_21_C249_n1354, CI => mult_21_C249_n1324, CO => 
                           mult_21_C249_n706, S => mult_21_C249_n707);
   mult_21_C249_U516 : ADFULD1 port map( A => mult_21_C249_n1246, B => 
                           mult_21_C249_n1296, CI => mult_21_C249_n1224, CO => 
                           mult_21_C249_n704, S => mult_21_C249_n705);
   mult_21_C249_U515 : ADFULD1 port map( A => mult_21_C249_n720, B => 
                           mult_21_C249_n1270, CI => mult_21_C249_n709, CO => 
                           mult_21_C249_n702, S => mult_21_C249_n703);
   mult_21_C249_U514 : ADFULD1 port map( A => mult_21_C249_n716, B => 
                           mult_21_C249_n718, CI => mult_21_C249_n707, CO => 
                           mult_21_C249_n700, S => mult_21_C249_n701);
   mult_21_C249_U513 : ADFULD1 port map( A => mult_21_C249_n703, B => 
                           mult_21_C249_n705, CI => mult_21_C249_n714, CO => 
                           mult_21_C249_n698, S => mult_21_C249_n699);
   mult_21_C249_U512 : ADFULD1 port map( A => mult_21_C249_n712, B => 
                           mult_21_C249_n701, CI => mult_21_C249_n699, CO => 
                           mult_21_C249_n696, S => mult_21_C249_n697);
   mult_21_C249_U510 : ADFULD1 port map( A => mult_21_C249_n1185, B => 
                           mult_21_C249_n1269, CI => mult_21_C249_n1223, CO => 
                           mult_21_C249_n692, S => mult_21_C249_n693);
   mult_21_C249_U509 : ADFULD1 port map( A => mult_21_C249_n1203, B => 
                           mult_21_C249_n1295, CI => mult_21_C249_n1245, CO => 
                           mult_21_C249_n690, S => mult_21_C249_n691);
   mult_21_C249_U508 : ADFULD1 port map( A => mult_21_C249_n695, B => 
                           mult_21_C249_n708, CI => mult_21_C249_n706, CO => 
                           mult_21_C249_n688, S => mult_21_C249_n689);
   mult_21_C249_U507 : ADFULD1 port map( A => mult_21_C249_n691, B => 
                           mult_21_C249_n704, CI => mult_21_C249_n693, CO => 
                           mult_21_C249_n686, S => mult_21_C249_n687);
   mult_21_C249_U506 : ADFULD1 port map( A => mult_21_C249_n700, B => 
                           mult_21_C249_n702, CI => mult_21_C249_n689, CO => 
                           mult_21_C249_n684, S => mult_21_C249_n685);
   mult_21_C249_U505 : ADFULD1 port map( A => mult_21_C249_n698, B => 
                           mult_21_C249_n687, CI => mult_21_C249_n685, CO => 
                           mult_21_C249_n682, S => mult_21_C249_n683);
   mult_21_C249_U503 : ADFULD1 port map( A => mult_21_C249_n1202, B => 
                           mult_21_C249_n1352, CI => mult_21_C249_n1322, CO => 
                           mult_21_C249_n678, S => mult_21_C249_n679);
   mult_21_C249_U502 : ADFULD1 port map( A => mult_21_C249_n1184, B => 
                           mult_21_C249_n1268, CI => mult_21_C249_n1222, CO => 
                           mult_21_C249_n676, S => mult_21_C249_n677);
   mult_21_C249_U501 : ADFULD1 port map( A => mult_21_C249_n1244, B => 
                           mult_21_C249_n1294, CI => mult_21_C249_n694, CO => 
                           mult_21_C249_n674, S => mult_21_C249_n675);
   mult_21_C249_U500 : ADFULD1 port map( A => mult_21_C249_n692, B => 
                           mult_21_C249_n681, CI => mult_21_C249_n690, CO => 
                           mult_21_C249_n672, S => mult_21_C249_n673);
   mult_21_C249_U499 : ADFULD1 port map( A => mult_21_C249_n677, B => 
                           mult_21_C249_n679, CI => mult_21_C249_n675, CO => 
                           mult_21_C249_n670, S => mult_21_C249_n671);
   mult_21_C249_U498 : ADFULD1 port map( A => mult_21_C249_n686, B => 
                           mult_21_C249_n688, CI => mult_21_C249_n673, CO => 
                           mult_21_C249_n668, S => mult_21_C249_n669);
   mult_21_C249_U497 : ADFULD1 port map( A => mult_21_C249_n684, B => 
                           mult_21_C249_n671, CI => mult_21_C249_n669, CO => 
                           mult_21_C249_n666, S => mult_21_C249_n667);
   mult_21_C249_U495 : ADFULD1 port map( A => mult_21_C249_n1167, B => 
                           mult_21_C249_n1201, CI => mult_21_C249_n1221, CO => 
                           mult_21_C249_n662, S => mult_21_C249_n663);
   mult_21_C249_U494 : ADFULD1 port map( A => mult_21_C249_n1243, B => 
                           mult_21_C249_n1183, CI => mult_21_C249_n1267, CO => 
                           mult_21_C249_n660, S => mult_21_C249_n661);
   mult_21_C249_U493 : ADFULD1 port map( A => mult_21_C249_n680, B => 
                           mult_21_C249_n1293, CI => mult_21_C249_n665, CO => 
                           mult_21_C249_n658, S => mult_21_C249_n659);
   mult_21_C249_U492 : ADFULD1 port map( A => mult_21_C249_n676, B => 
                           mult_21_C249_n678, CI => mult_21_C249_n674, CO => 
                           mult_21_C249_n656, S => mult_21_C249_n657);
   mult_21_C249_U491 : ADFULD1 port map( A => mult_21_C249_n663, B => 
                           mult_21_C249_n661, CI => mult_21_C249_n672, CO => 
                           mult_21_C249_n654, S => mult_21_C249_n655);
   mult_21_C249_U490 : ADFULD1 port map( A => mult_21_C249_n670, B => 
                           mult_21_C249_n659, CI => mult_21_C249_n657, CO => 
                           mult_21_C249_n652, S => mult_21_C249_n653);
   mult_21_C249_U489 : ADFULD1 port map( A => mult_21_C249_n668, B => 
                           mult_21_C249_n655, CI => mult_21_C249_n653, CO => 
                           mult_21_C249_n650, S => mult_21_C249_n651);
   mult_21_C249_U487 : ADFULD1 port map( A => mult_21_C249_n1200, B => 
                           mult_21_C249_n1350, CI => mult_21_C249_n1320, CO => 
                           mult_21_C249_n646, S => mult_21_C249_n647);
   mult_21_C249_U486 : ADFULD1 port map( A => mult_21_C249_n1166, B => 
                           mult_21_C249_n1266, CI => mult_21_C249_n1220, CO => 
                           mult_21_C249_n644, S => mult_21_C249_n645);
   mult_21_C249_U485 : ADFULD1 port map( A => mult_21_C249_n1182, B => 
                           mult_21_C249_n1292, CI => mult_21_C249_n1242, CO => 
                           mult_21_C249_n642, S => mult_21_C249_n643);
   mult_21_C249_U484 : ADFULD1 port map( A => mult_21_C249_n649, B => 
                           mult_21_C249_n664, CI => mult_21_C249_n662, CO => 
                           mult_21_C249_n640, S => mult_21_C249_n641);
   mult_21_C249_U483 : ADFULD1 port map( A => mult_21_C249_n647, B => 
                           mult_21_C249_n660, CI => mult_21_C249_n643, CO => 
                           mult_21_C249_n638, S => mult_21_C249_n639);
   mult_21_C249_U482 : ADFULD1 port map( A => mult_21_C249_n658, B => 
                           mult_21_C249_n645, CI => mult_21_C249_n656, CO => 
                           mult_21_C249_n636, S => mult_21_C249_n637);
   mult_21_C249_U481 : ADFULD1 port map( A => mult_21_C249_n639, B => 
                           mult_21_C249_n641, CI => mult_21_C249_n654, CO => 
                           mult_21_C249_n634, S => mult_21_C249_n635);
   mult_21_C249_U480 : ADFULD1 port map( A => mult_21_C249_n652, B => 
                           mult_21_C249_n637, CI => mult_21_C249_n635, CO => 
                           mult_21_C249_n632, S => mult_21_C249_n633);
   mult_21_C249_U478 : ADFULD1 port map( A => mult_21_C249_n1151, B => 
                           mult_21_C249_n1199, CI => mult_21_C249_n1219, CO => 
                           mult_21_C249_n628, S => mult_21_C249_n629);
   mult_21_C249_U477 : ADFULD1 port map( A => mult_21_C249_n1291, B => 
                           mult_21_C249_n1181, CI => mult_21_C249_n1165, CO => 
                           mult_21_C249_n626, S => mult_21_C249_n627);
   mult_21_C249_U476 : ADFULD1 port map( A => mult_21_C249_n1241, B => 
                           mult_21_C249_n1265, CI => mult_21_C249_n648, CO => 
                           mult_21_C249_n624, S => mult_21_C249_n625);
   mult_21_C249_U475 : ADFULD1 port map( A => mult_21_C249_n646, B => 
                           mult_21_C249_n631, CI => mult_21_C249_n642, CO => 
                           mult_21_C249_n622, S => mult_21_C249_n623);
   mult_21_C249_U474 : ADFULD1 port map( A => mult_21_C249_n627, B => 
                           mult_21_C249_n644, CI => mult_21_C249_n629, CO => 
                           mult_21_C249_n620, S => mult_21_C249_n621);
   mult_21_C249_U473 : ADFULD1 port map( A => mult_21_C249_n640, B => 
                           mult_21_C249_n625, CI => mult_21_C249_n638, CO => 
                           mult_21_C249_n618, S => mult_21_C249_n619);
   mult_21_C249_U472 : ADFULD1 port map( A => mult_21_C249_n621, B => 
                           mult_21_C249_n623, CI => mult_21_C249_n636, CO => 
                           mult_21_C249_n616, S => mult_21_C249_n617);
   mult_21_C249_U471 : ADFULD1 port map( A => mult_21_C249_n634, B => 
                           mult_21_C249_n619, CI => mult_21_C249_n617, CO => 
                           mult_21_C249_n614, S => mult_21_C249_n615);
   mult_21_C249_U469 : ADFULD1 port map( A => mult_21_C249_n1164, B => 
                           mult_21_C249_n1348, CI => mult_21_C249_n1318, CO => 
                           mult_21_C249_n610, S => mult_21_C249_n611);
   mult_21_C249_U468 : ADFULD1 port map( A => mult_21_C249_n1290, B => 
                           mult_21_C249_n1198, CI => mult_21_C249_n1218, CO => 
                           mult_21_C249_n608, S => mult_21_C249_n609);
   mult_21_C249_U467 : ADFULD1 port map( A => mult_21_C249_n1150, B => 
                           mult_21_C249_n1264, CI => mult_21_C249_n1180, CO => 
                           mult_21_C249_n606, S => mult_21_C249_n607);
   mult_21_C249_U466 : ADFULD1 port map( A => mult_21_C249_n630, B => 
                           mult_21_C249_n1240, CI => mult_21_C249_n613, CO => 
                           mult_21_C249_n604, S => mult_21_C249_n605);
   mult_21_C249_U465 : ADFULD1 port map( A => mult_21_C249_n626, B => 
                           mult_21_C249_n628, CI => mult_21_C249_n624, CO => 
                           mult_21_C249_n602, S => mult_21_C249_n603);
   mult_21_C249_U464 : ADFULD1 port map( A => mult_21_C249_n609, B => 
                           mult_21_C249_n611, CI => mult_21_C249_n607, CO => 
                           mult_21_C249_n600, S => mult_21_C249_n601);
   mult_21_C249_U463 : ADFULD1 port map( A => mult_21_C249_n622, B => 
                           mult_21_C249_n605, CI => mult_21_C249_n620, CO => 
                           mult_21_C249_n598, S => mult_21_C249_n599);
   mult_21_C249_U462 : ADFULD1 port map( A => mult_21_C249_n601, B => 
                           mult_21_C249_n603, CI => mult_21_C249_n618, CO => 
                           mult_21_C249_n596, S => mult_21_C249_n597);
   mult_21_C249_U461 : ADFULD1 port map( A => mult_21_C249_n616, B => 
                           mult_21_C249_n599, CI => mult_21_C249_n597, CO => 
                           mult_21_C249_n594, S => mult_21_C249_n595);
   mult_21_C249_U459 : ADFULD1 port map( A => mult_21_C249_n1137, B => 
                           mult_21_C249_n1179, CI => mult_21_C249_n1217, CO => 
                           mult_21_C249_n590, S => mult_21_C249_n591);
   mult_21_C249_U458 : ADFULD1 port map( A => mult_21_C249_n1289, B => 
                           mult_21_C249_n1163, CI => mult_21_C249_n1149, CO => 
                           mult_21_C249_n588, S => mult_21_C249_n589);
   mult_21_C249_U457 : ADFULD1 port map( A => mult_21_C249_n1197, B => 
                           mult_21_C249_n1263, CI => mult_21_C249_n1239, CO => 
                           mult_21_C249_n586, S => mult_21_C249_n587);
   mult_21_C249_U456 : ADFULD1 port map( A => mult_21_C249_n593, B => 
                           mult_21_C249_n612, CI => mult_21_C249_n610, CO => 
                           mult_21_C249_n584, S => mult_21_C249_n585);
   mult_21_C249_U455 : ADFULD1 port map( A => mult_21_C249_n606, B => 
                           mult_21_C249_n608, CI => mult_21_C249_n587, CO => 
                           mult_21_C249_n582, S => mult_21_C249_n583);
   mult_21_C249_U454 : ADFULD1 port map( A => mult_21_C249_n591, B => 
                           mult_21_C249_n589, CI => mult_21_C249_n604, CO => 
                           mult_21_C249_n580, S => mult_21_C249_n581);
   mult_21_C249_U453 : ADFULD1 port map( A => mult_21_C249_n585, B => 
                           mult_21_C249_n602, CI => mult_21_C249_n600, CO => 
                           mult_21_C249_n578, S => mult_21_C249_n579);
   mult_21_C249_U452 : ADFULD1 port map( A => mult_21_C249_n581, B => 
                           mult_21_C249_n583, CI => mult_21_C249_n598, CO => 
                           mult_21_C249_n576, S => mult_21_C249_n577);
   mult_21_C249_U451 : ADFULD1 port map( A => mult_21_C249_n596, B => 
                           mult_21_C249_n579, CI => mult_21_C249_n577, CO => 
                           mult_21_C249_n574, S => mult_21_C249_n575);
   mult_21_C249_U449 : ADFULD1 port map( A => mult_21_C249_n1136, B => 
                           mult_21_C249_n1346, CI => mult_21_C249_n1316, CO => 
                           mult_21_C249_n570, S => mult_21_C249_n571);
   mult_21_C249_U448 : ADFULD1 port map( A => mult_21_C249_n1288, B => 
                           mult_21_C249_n1178, CI => mult_21_C249_n1216, CO => 
                           mult_21_C249_n568, S => mult_21_C249_n569);
   mult_21_C249_U447 : ADFULD1 port map( A => mult_21_C249_n1148, B => 
                           mult_21_C249_n1262, CI => mult_21_C249_n1162, CO => 
                           mult_21_C249_n566, S => mult_21_C249_n567);
   mult_21_C249_U446 : ADFULD1 port map( A => mult_21_C249_n1196, B => 
                           mult_21_C249_n1238, CI => mult_21_C249_n592, CO => 
                           mult_21_C249_n564, S => mult_21_C249_n565);
   mult_21_C249_U445 : ADFULD1 port map( A => mult_21_C249_n590, B => 
                           mult_21_C249_n573, CI => mult_21_C249_n588, CO => 
                           mult_21_C249_n562, S => mult_21_C249_n563);
   mult_21_C249_U444 : ADFULD1 port map( A => mult_21_C249_n571, B => 
                           mult_21_C249_n586, CI => mult_21_C249_n567, CO => 
                           mult_21_C249_n560, S => mult_21_C249_n561);
   mult_21_C249_U443 : ADFULD1 port map( A => mult_21_C249_n565, B => 
                           mult_21_C249_n569, CI => mult_21_C249_n584, CO => 
                           mult_21_C249_n558, S => mult_21_C249_n559);
   mult_21_C249_U442 : ADFULD1 port map( A => mult_21_C249_n563, B => 
                           mult_21_C249_n582, CI => mult_21_C249_n580, CO => 
                           mult_21_C249_n556, S => mult_21_C249_n557);
   mult_21_C249_U441 : ADFULD1 port map( A => mult_21_C249_n559, B => 
                           mult_21_C249_n561, CI => mult_21_C249_n578, CO => 
                           mult_21_C249_n554, S => mult_21_C249_n555);
   mult_21_C249_U440 : ADFULD1 port map( A => mult_21_C249_n576, B => 
                           mult_21_C249_n557, CI => mult_21_C249_n555, CO => 
                           mult_21_C249_n552, S => mult_21_C249_n553);
   mult_21_C249_U438 : ADFULD1 port map( A => mult_21_C249_n1125, B => 
                           mult_21_C249_n1177, CI => mult_21_C249_n1215, CO => 
                           mult_21_C249_n548, S => mult_21_C249_n549);
   mult_21_C249_U437 : ADFULD1 port map( A => mult_21_C249_n1287, B => 
                           mult_21_C249_n1161, CI => mult_21_C249_n1261, CO => 
                           mult_21_C249_n546, S => mult_21_C249_n547);
   mult_21_C249_U436 : ADFULD1 port map( A => mult_21_C249_n1135, B => 
                           mult_21_C249_n1237, CI => mult_21_C249_n1147, CO => 
                           mult_21_C249_n544, S => mult_21_C249_n545);
   mult_21_C249_U435 : ADFULD1 port map( A => mult_21_C249_n572, B => 
                           mult_21_C249_n1195, CI => mult_21_C249_n551, CO => 
                           mult_21_C249_n542, S => mult_21_C249_n543);
   mult_21_C249_U434 : ADFULD1 port map( A => mult_21_C249_n566, B => 
                           mult_21_C249_n570, CI => mult_21_C249_n568, CO => 
                           mult_21_C249_n540, S => mult_21_C249_n541);
   mult_21_C249_U433 : ADFULD1 port map( A => mult_21_C249_n549, B => 
                           mult_21_C249_n564, CI => mult_21_C249_n547, CO => 
                           mult_21_C249_n538, S => mult_21_C249_n539);
   mult_21_C249_U432 : ADFULD1 port map( A => mult_21_C249_n562, B => 
                           mult_21_C249_n545, CI => mult_21_C249_n543, CO => 
                           mult_21_C249_n536, S => mult_21_C249_n537);
   mult_21_C249_U431 : ADFULD1 port map( A => mult_21_C249_n541, B => 
                           mult_21_C249_n560, CI => mult_21_C249_n558, CO => 
                           mult_21_C249_n534, S => mult_21_C249_n535);
   mult_21_C249_U430 : ADFULD1 port map( A => mult_21_C249_n556, B => 
                           mult_21_C249_n539, CI => mult_21_C249_n537, CO => 
                           mult_21_C249_n532, S => mult_21_C249_n533);
   mult_21_C249_U429 : ADFULD1 port map( A => mult_21_C249_n554, B => 
                           mult_21_C249_n535, CI => mult_21_C249_n533, CO => 
                           mult_21_C249_n530, S => mult_21_C249_n531);
   mult_21_C249_U427 : ADFULD1 port map( A => mult_21_C249_n1146, B => 
                           mult_21_C249_n1344, CI => mult_21_C249_n1314, CO => 
                           mult_21_C249_n526, S => mult_21_C249_n527);
   mult_21_C249_U426 : ADFULD1 port map( A => mult_21_C249_n1124, B => 
                           mult_21_C249_n1176, CI => mult_21_C249_n1214, CO => 
                           mult_21_C249_n524, S => mult_21_C249_n525);
   mult_21_C249_U425 : ADFULD1 port map( A => mult_21_C249_n1134, B => 
                           mult_21_C249_n1286, CI => mult_21_C249_n1160, CO => 
                           mult_21_C249_n522, S => mult_21_C249_n523);
   mult_21_C249_U424 : ADFULD1 port map( A => mult_21_C249_n1194, B => 
                           mult_21_C249_n1260, CI => mult_21_C249_n1236, CO => 
                           mult_21_C249_n520, S => mult_21_C249_n521);
   mult_21_C249_U423 : ADFULD1 port map( A => mult_21_C249_n529, B => 
                           mult_21_C249_n550, CI => mult_21_C249_n548, CO => 
                           mult_21_C249_n518, S => mult_21_C249_n519);
   mult_21_C249_U422 : ADFULD1 port map( A => mult_21_C249_n544, B => 
                           mult_21_C249_n546, CI => mult_21_C249_n527, CO => 
                           mult_21_C249_n516, S => mult_21_C249_n517);
   mult_21_C249_U421 : ADFULD1 port map( A => mult_21_C249_n525, B => 
                           mult_21_C249_n521, CI => mult_21_C249_n523, CO => 
                           mult_21_C249_n514, S => mult_21_C249_n515);
   mult_21_C249_U420 : ADFULD1 port map( A => mult_21_C249_n540, B => 
                           mult_21_C249_n542, CI => mult_21_C249_n519, CO => 
                           mult_21_C249_n512, S => mult_21_C249_n513);
   mult_21_C249_U419 : ADFULD1 port map( A => mult_21_C249_n517, B => 
                           mult_21_C249_n538, CI => mult_21_C249_n515, CO => 
                           mult_21_C249_n510, S => mult_21_C249_n511);
   mult_21_C249_U418 : ADFULD1 port map( A => mult_21_C249_n513, B => 
                           mult_21_C249_n536, CI => mult_21_C249_n534, CO => 
                           mult_21_C249_n508, S => mult_21_C249_n509);
   mult_21_C249_U417 : ADFULD1 port map( A => mult_21_C249_n532, B => 
                           mult_21_C249_n511, CI => mult_21_C249_n509, CO => 
                           mult_21_C249_n506, S => mult_21_C249_n507);
   mult_21_C249_U415 : ADFULD1 port map( A => mult_21_C249_n1115, B => 
                           mult_21_C249_n1175, CI => mult_21_C249_n1213, CO => 
                           mult_21_C249_n502, S => mult_21_C249_n503);
   mult_21_C249_U414 : ADFULD1 port map( A => mult_21_C249_n1123, B => 
                           mult_21_C249_n1145, CI => mult_21_C249_n1133, CO => 
                           mult_21_C249_n500, S => mult_21_C249_n501);
   mult_21_C249_U413 : ADFULD1 port map( A => mult_21_C249_n1159, B => 
                           mult_21_C249_n1285, CI => mult_21_C249_n1193, CO => 
                           mult_21_C249_n498, S => mult_21_C249_n499);
   mult_21_C249_U412 : ADFULD1 port map( A => mult_21_C249_n1235, B => 
                           mult_21_C249_n1259, CI => mult_21_C249_n528, CO => 
                           mult_21_C249_n496, S => mult_21_C249_n497);
   mult_21_C249_U411 : ADFULD1 port map( A => mult_21_C249_n526, B => 
                           mult_21_C249_n505, CI => mult_21_C249_n520, CO => 
                           mult_21_C249_n494, S => mult_21_C249_n495);
   mult_21_C249_U410 : ADFULD1 port map( A => mult_21_C249_n522, B => 
                           mult_21_C249_n524, CI => mult_21_C249_n499, CO => 
                           mult_21_C249_n492, S => mult_21_C249_n493);
   mult_21_C249_U409 : ADFULD1 port map( A => mult_21_C249_n501, B => 
                           mult_21_C249_n503, CI => mult_21_C249_n497, CO => 
                           mult_21_C249_n490, S => mult_21_C249_n491);
   mult_21_C249_U408 : ADFULD1 port map( A => mult_21_C249_n516, B => 
                           mult_21_C249_n518, CI => mult_21_C249_n495, CO => 
                           mult_21_C249_n488, S => mult_21_C249_n489);
   mult_21_C249_U407 : ADFULD1 port map( A => mult_21_C249_n493, B => 
                           mult_21_C249_n514, CI => mult_21_C249_n491, CO => 
                           mult_21_C249_n486, S => mult_21_C249_n487);
   mult_21_C249_U406 : ADFULD1 port map( A => mult_21_C249_n510, B => 
                           mult_21_C249_n512, CI => mult_21_C249_n489, CO => 
                           mult_21_C249_n484, S => mult_21_C249_n485);
   mult_21_C249_U405 : ADFULD1 port map( A => mult_21_C249_n508, B => 
                           mult_21_C249_n487, CI => mult_21_C249_n485, CO => 
                           mult_21_C249_n482, S => mult_21_C249_n483);
   mult_21_C249_U403 : ADFULD1 port map( A => mult_21_C249_n1114, B => 
                           mult_21_C249_n1342, CI => mult_21_C249_n1312, CO => 
                           mult_21_C249_n478, S => mult_21_C249_n479);
   mult_21_C249_U402 : ADFULD1 port map( A => mult_21_C249_n1284, B => 
                           mult_21_C249_n1174, CI => mult_21_C249_n1212, CO => 
                           mult_21_C249_n476, S => mult_21_C249_n477);
   mult_21_C249_U401 : ADFULD1 port map( A => mult_21_C249_n1258, B => 
                           mult_21_C249_n1132, CI => mult_21_C249_n1122, CO => 
                           mult_21_C249_n474, S => mult_21_C249_n475);
   mult_21_C249_U400 : ADFULD1 port map( A => mult_21_C249_n1144, B => 
                           mult_21_C249_n1234, CI => mult_21_C249_n1158, CO => 
                           mult_21_C249_n472, S => mult_21_C249_n473);
   mult_21_C249_U399 : ADFULD1 port map( A => mult_21_C249_n504, B => 
                           mult_21_C249_n1192, CI => mult_21_C249_n481, CO => 
                           mult_21_C249_n470, S => mult_21_C249_n471);
   mult_21_C249_U398 : ADFULD1 port map( A => mult_21_C249_n498, B => 
                           mult_21_C249_n502, CI => mult_21_C249_n496, CO => 
                           mult_21_C249_n468, S => mult_21_C249_n469);
   mult_21_C249_U397 : ADFULD1 port map( A => mult_21_C249_n479, B => 
                           mult_21_C249_n500, CI => mult_21_C249_n473, CO => 
                           mult_21_C249_n466, S => mult_21_C249_n467);
   mult_21_C249_U396 : ADFULD1 port map( A => mult_21_C249_n475, B => 
                           mult_21_C249_n477, CI => mult_21_C249_n471, CO => 
                           mult_21_C249_n464, S => mult_21_C249_n465);
   mult_21_C249_U395 : ADFULD1 port map( A => mult_21_C249_n492, B => 
                           mult_21_C249_n494, CI => mult_21_C249_n490, CO => 
                           mult_21_C249_n462, S => mult_21_C249_n463);
   mult_21_C249_U394 : ADFULD1 port map( A => mult_21_C249_n467, B => 
                           mult_21_C249_n469, CI => mult_21_C249_n465, CO => 
                           mult_21_C249_n460, S => mult_21_C249_n461);
   mult_21_C249_U393 : ADFULD1 port map( A => mult_21_C249_n486, B => 
                           mult_21_C249_n488, CI => mult_21_C249_n463, CO => 
                           mult_21_C249_n458, S => mult_21_C249_n459);
   mult_21_C249_U392 : ADFULD1 port map( A => mult_21_C249_n484, B => 
                           mult_21_C249_n461, CI => mult_21_C249_n459, CO => 
                           mult_21_C249_n456, S => mult_21_C249_n457);
   mult_21_C249_U390 : ADFULD1 port map( A => mult_21_C249_n1107, B => 
                           mult_21_C249_n1157, CI => mult_21_C249_n1211, CO => 
                           mult_21_C249_n452, S => mult_21_C249_n453);
   mult_21_C249_U389 : ADFULD1 port map( A => mult_21_C249_n1283, B => 
                           mult_21_C249_n1143, CI => mult_21_C249_n1257, CO => 
                           mult_21_C249_n450, S => mult_21_C249_n451);
   mult_21_C249_U388 : ADFULD1 port map( A => mult_21_C249_n1113, B => 
                           mult_21_C249_n1233, CI => mult_21_C249_n1121, CO => 
                           mult_21_C249_n448, S => mult_21_C249_n449);
   mult_21_C249_U387 : ADFULD1 port map( A => mult_21_C249_n1131, B => 
                           mult_21_C249_n1191, CI => mult_21_C249_n1173, CO => 
                           mult_21_C249_n446, S => mult_21_C249_n447);
   mult_21_C249_U386 : ADFULD1 port map( A => mult_21_C249_n455, B => 
                           mult_21_C249_n480, CI => mult_21_C249_n478, CO => 
                           mult_21_C249_n444, S => mult_21_C249_n445);
   mult_21_C249_U385 : ADFULD1 port map( A => mult_21_C249_n474, B => 
                           mult_21_C249_n472, CI => mult_21_C249_n476, CO => 
                           mult_21_C249_n442, S => mult_21_C249_n443);
   mult_21_C249_U384 : ADFULD1 port map( A => mult_21_C249_n453, B => 
                           mult_21_C249_n447, CI => mult_21_C249_n470, CO => 
                           mult_21_C249_n440, S => mult_21_C249_n441);
   mult_21_C249_U383 : ADFULD1 port map( A => mult_21_C249_n449, B => 
                           mult_21_C249_n451, CI => mult_21_C249_n468, CO => 
                           mult_21_C249_n438, S => mult_21_C249_n439);
   mult_21_C249_U382 : ADFULD1 port map( A => mult_21_C249_n466, B => 
                           mult_21_C249_n445, CI => mult_21_C249_n443, CO => 
                           mult_21_C249_n436, S => mult_21_C249_n437);
   mult_21_C249_U381 : ADFULD1 port map( A => mult_21_C249_n441, B => 
                           mult_21_C249_n464, CI => mult_21_C249_n462, CO => 
                           mult_21_C249_n434, S => mult_21_C249_n435);
   mult_21_C249_U380 : ADFULD1 port map( A => mult_21_C249_n437, B => 
                           mult_21_C249_n439, CI => mult_21_C249_n460, CO => 
                           mult_21_C249_n432, S => mult_21_C249_n433);
   mult_21_C249_U379 : ADFULD1 port map( A => mult_21_C249_n458, B => 
                           mult_21_C249_n435, CI => mult_21_C249_n433, CO => 
                           mult_21_C249_n430, S => mult_21_C249_n431);
   mult_21_C249_U377 : ADFULD1 port map( A => mult_21_C249_n1106, B => 
                           mult_21_C249_n1340, CI => mult_21_C249_n1310, CO => 
                           mult_21_C249_n426, S => mult_21_C249_n427);
   mult_21_C249_U376 : ADFULD1 port map( A => mult_21_C249_n1282, B => 
                           mult_21_C249_n1156, CI => mult_21_C249_n1210, CO => 
                           mult_21_C249_n424, S => mult_21_C249_n425);
   mult_21_C249_U375 : ADFULD1 port map( A => mult_21_C249_n1112, B => 
                           mult_21_C249_n1130, CI => mult_21_C249_n1120, CO => 
                           mult_21_C249_n422, S => mult_21_C249_n423);
   mult_21_C249_U374 : ADFULD1 port map( A => mult_21_C249_n1142, B => 
                           mult_21_C249_n1256, CI => mult_21_C249_n1172, CO => 
                           mult_21_C249_n420, S => mult_21_C249_n421);
   mult_21_C249_U373 : ADFULD1 port map( A => mult_21_C249_n1232, B => 
                           mult_21_C249_n1190, CI => mult_21_C249_n454, CO => 
                           mult_21_C249_n418, S => mult_21_C249_n419);
   mult_21_C249_U372 : ADFULD1 port map( A => mult_21_C249_n452, B => 
                           mult_21_C249_n429, CI => mult_21_C249_n450, CO => 
                           mult_21_C249_n416, S => mult_21_C249_n417);
   mult_21_C249_U371 : ADFULD1 port map( A => mult_21_C249_n448, B => 
                           mult_21_C249_n446, CI => mult_21_C249_n427, CO => 
                           mult_21_C249_n414, S => mult_21_C249_n415);
   mult_21_C249_U370 : ADFULD1 port map( A => mult_21_C249_n421, B => 
                           mult_21_C249_n423, CI => mult_21_C249_n425, CO => 
                           mult_21_C249_n412, S => mult_21_C249_n413);
   mult_21_C249_U369 : ADFULD1 port map( A => mult_21_C249_n444, B => 
                           mult_21_C249_n419, CI => mult_21_C249_n442, CO => 
                           mult_21_C249_n410, S => mult_21_C249_n411);
   mult_21_C249_U368 : ADFULD1 port map( A => mult_21_C249_n440, B => 
                           mult_21_C249_n417, CI => mult_21_C249_n415, CO => 
                           mult_21_C249_n408, S => mult_21_C249_n409);
   mult_21_C249_U367 : ADFULD1 port map( A => mult_21_C249_n438, B => 
                           mult_21_C249_n413, CI => mult_21_C249_n411, CO => 
                           mult_21_C249_n406, S => mult_21_C249_n407);
   mult_21_C249_U366 : ADFULD1 port map( A => mult_21_C249_n409, B => 
                           mult_21_C249_n436, CI => mult_21_C249_n434, CO => 
                           mult_21_C249_n404, S => mult_21_C249_n405);
   mult_21_C249_U365 : ADFULD1 port map( A => mult_21_C249_n432, B => 
                           mult_21_C249_n407, CI => mult_21_C249_n405, CO => 
                           mult_21_C249_n402, S => mult_21_C249_n403);
   mult_21_C249_U363 : ADFULD1 port map( A => mult_21_C249_n1101, B => 
                           mult_21_C249_n1155, CI => mult_21_C249_n1209, CO => 
                           mult_21_C249_n398, S => mult_21_C249_n399);
   mult_21_C249_U362 : ADFULD1 port map( A => mult_21_C249_n1281, B => 
                           mult_21_C249_n1129, CI => mult_21_C249_n1105, CO => 
                           mult_21_C249_n396, S => mult_21_C249_n397);
   mult_21_C249_U361 : ADFULD1 port map( A => mult_21_C249_n1255, B => 
                           mult_21_C249_n1119, CI => mult_21_C249_n1111, CO => 
                           mult_21_C249_n394, S => mult_21_C249_n395);
   mult_21_C249_U360 : ADFULD1 port map( A => mult_21_C249_n1141, B => 
                           mult_21_C249_n1231, CI => mult_21_C249_n1171, CO => 
                           mult_21_C249_n392, S => mult_21_C249_n393);
   mult_21_C249_U359 : ADFULD1 port map( A => mult_21_C249_n428, B => 
                           mult_21_C249_n1189, CI => mult_21_C249_n401, CO => 
                           mult_21_C249_n390, S => mult_21_C249_n391);
   mult_21_C249_U358 : ADFULD1 port map( A => mult_21_C249_n424, B => 
                           mult_21_C249_n426, CI => mult_21_C249_n420, CO => 
                           mult_21_C249_n388, S => mult_21_C249_n389);
   mult_21_C249_U357 : ADFULD1 port map( A => mult_21_C249_n418, B => 
                           mult_21_C249_n422, CI => mult_21_C249_n393, CO => 
                           mult_21_C249_n386, S => mult_21_C249_n387);
   mult_21_C249_U356 : ADFULD1 port map( A => mult_21_C249_n395, B => 
                           mult_21_C249_n397, CI => mult_21_C249_n399, CO => 
                           mult_21_C249_n384, S => mult_21_C249_n385);
   mult_21_C249_U355 : ADFULD1 port map( A => mult_21_C249_n391, B => 
                           mult_21_C249_n416, CI => mult_21_C249_n414, CO => 
                           mult_21_C249_n382, S => mult_21_C249_n383);
   mult_21_C249_U354 : ADFULD1 port map( A => mult_21_C249_n412, B => 
                           mult_21_C249_n389, CI => mult_21_C249_n387, CO => 
                           mult_21_C249_n380, S => mult_21_C249_n381);
   mult_21_C249_U353 : ADFULD1 port map( A => mult_21_C249_n410, B => 
                           mult_21_C249_n385, CI => mult_21_C249_n383, CO => 
                           mult_21_C249_n378, S => mult_21_C249_n379);
   mult_21_C249_U352 : ADFULD1 port map( A => mult_21_C249_n381, B => 
                           mult_21_C249_n408, CI => mult_21_C249_n406, CO => 
                           mult_21_C249_n376, S => mult_21_C249_n377);
   mult_21_C249_U351 : ADFULD1 port map( A => mult_21_C249_n404, B => 
                           mult_21_C249_n379, CI => mult_21_C249_n377, CO => 
                           mult_21_C249_n374, S => mult_21_C249_n375);
   mult_21_C249_U349 : ADFULD1 port map( A => mult_21_C249_n1100, B => 
                           mult_21_C249_n1338, CI => mult_21_C249_n1308, CO => 
                           mult_21_C249_n370, S => mult_21_C249_n371);
   mult_21_C249_U348 : ADFULD1 port map( A => mult_21_C249_n1280, B => 
                           mult_21_C249_n1154, CI => mult_21_C249_n1208, CO => 
                           mult_21_C249_n368, S => mult_21_C249_n369);
   mult_21_C249_U347 : ADFULD1 port map( A => mult_21_C249_n1254, B => 
                           mult_21_C249_n1128, CI => mult_21_C249_n1230, CO => 
                           mult_21_C249_n366, S => mult_21_C249_n367);
   mult_21_C249_U346 : ADFULD1 port map( A => mult_21_C249_n1104, B => 
                           mult_21_C249_n1188, CI => mult_21_C249_n1110, CO => 
                           mult_21_C249_n364, S => mult_21_C249_n365);
   mult_21_C249_U345 : ADFULD1 port map( A => mult_21_C249_n1170, B => 
                           mult_21_C249_n1118, CI => mult_21_C249_n1140, CO => 
                           mult_21_C249_n362, S => mult_21_C249_n363);
   mult_21_C249_U344 : ADFULD1 port map( A => mult_21_C249_n373, B => 
                           mult_21_C249_n400, CI => mult_21_C249_n392, CO => 
                           mult_21_C249_n360, S => mult_21_C249_n361);
   mult_21_C249_U343 : ADFULD1 port map( A => mult_21_C249_n398, B => 
                           mult_21_C249_n394, CI => mult_21_C249_n396, CO => 
                           mult_21_C249_n358, S => mult_21_C249_n359);
   mult_21_C249_U342 : ADFULD1 port map( A => mult_21_C249_n369, B => 
                           mult_21_C249_n371, CI => mult_21_C249_n367, CO => 
                           mult_21_C249_n356, S => mult_21_C249_n357);
   mult_21_C249_U341 : ADFULD1 port map( A => mult_21_C249_n365, B => 
                           mult_21_C249_n363, CI => mult_21_C249_n390, CO => 
                           mult_21_C249_n354, S => mult_21_C249_n355);
   mult_21_C249_U340 : ADFULD1 port map( A => mult_21_C249_n361, B => 
                           mult_21_C249_n388, CI => mult_21_C249_n386, CO => 
                           mult_21_C249_n352, S => mult_21_C249_n353);
   mult_21_C249_U339 : ADFULD1 port map( A => mult_21_C249_n359, B => 
                           mult_21_C249_n384, CI => mult_21_C249_n357, CO => 
                           mult_21_C249_n350, S => mult_21_C249_n351);
   mult_21_C249_U338 : ADFULD1 port map( A => mult_21_C249_n382, B => 
                           mult_21_C249_n355, CI => mult_21_C249_n380, CO => 
                           mult_21_C249_n348, S => mult_21_C249_n349);
   mult_21_C249_U337 : ADFULD1 port map( A => mult_21_C249_n351, B => 
                           mult_21_C249_n353, CI => mult_21_C249_n378, CO => 
                           mult_21_C249_n346, S => mult_21_C249_n347);
   mult_21_C249_U336 : ADFULD1 port map( A => mult_21_C249_n376, B => 
                           mult_21_C249_n349, CI => mult_21_C249_n347, CO => 
                           mult_21_C249_n344, S => mult_21_C249_n345);
   mult_21_C249_U334 : EXOR3D1 port map( A1 => mult_21_C249_n1097, A2 => 
                           mult_21_C249_n1279, A3 => mult_21_C249_n1207, Z => 
                           mult_21_C249_n342);
   mult_21_C249_U333 : EXOR3D1 port map( A1 => mult_21_C249_n1253, A2 => 
                           mult_21_C249_n1127, A3 => mult_21_C249_n1099, Z => 
                           mult_21_C249_n341);
   mult_21_C249_U332 : EXOR3D1 port map( A1 => mult_21_C249_n1103, A2 => 
                           mult_21_C249_n1117, A3 => mult_21_C249_n1109, Z => 
                           mult_21_C249_n340);
   mult_21_C249_U331 : EXOR3D1 port map( A1 => mult_21_C249_n1139, A2 => 
                           mult_21_C249_n1229, A3 => mult_21_C249_n1153, Z => 
                           mult_21_C249_n339);
   mult_21_C249_U330 : EXOR3D1 port map( A1 => mult_21_C249_n1187, A2 => 
                           mult_21_C249_n1169, A3 => mult_21_C249_n372, Z => 
                           mult_21_C249_n338);
   mult_21_C249_U329 : EXOR3D1 port map( A1 => mult_21_C249_n368, A2 => 
                           mult_21_C249_n370, A3 => mult_21_C249_n364, Z => 
                           mult_21_C249_n337);
   mult_21_C249_U328 : EXOR3D1 port map( A1 => mult_21_C249_n366, A2 => 
                           mult_21_C249_n343, A3 => mult_21_C249_n362, Z => 
                           mult_21_C249_n336);
   mult_21_C249_U327 : EXOR3D1 port map( A1 => mult_21_C249_n342, A2 => 
                           mult_21_C249_n338, A3 => mult_21_C249_n341, Z => 
                           mult_21_C249_n335);
   mult_21_C249_U326 : EXOR3D1 port map( A1 => mult_21_C249_n339, A2 => 
                           mult_21_C249_n340, A3 => mult_21_C249_n360, Z => 
                           mult_21_C249_n334);
   mult_21_C249_U325 : EXOR3D1 port map( A1 => mult_21_C249_n337, A2 => 
                           mult_21_C249_n358, A3 => mult_21_C249_n336, Z => 
                           mult_21_C249_n333);
   mult_21_C249_U324 : EXOR3D1 port map( A1 => mult_21_C249_n354, A2 => 
                           mult_21_C249_n356, A3 => mult_21_C249_n335, Z => 
                           mult_21_C249_n332);
   mult_21_C249_U323 : EXOR3D1 port map( A1 => mult_21_C249_n352, A2 => 
                           mult_21_C249_n334, A3 => mult_21_C249_n333, Z => 
                           mult_21_C249_n331);
   mult_21_C249_U322 : EXOR3D1 port map( A1 => mult_21_C249_n332, A2 => 
                           mult_21_C249_n350, A3 => mult_21_C249_n348, Z => 
                           mult_21_C249_n330);
   mult_21_C249_U321 : EXOR3D1 port map( A1 => mult_21_C249_n346, A2 => 
                           mult_21_C249_n331, A3 => mult_21_C249_n330, Z => 
                           mult_21_C249_n329);
   mult_21_C249_U313 : EXOR2D1 port map( A1 => mult_21_C249_n303, A2 => 
                           mult_21_C249_n305, Z => N3362);
   mult_21_C249_U305 : EXNOR2D1 port map( A1 => mult_21_C249_n176, A2 => 
                           mult_21_C249_n302, Z => N3363);
   mult_21_C249_U300 : OAI21D1 port map( A1 => mult_21_C249_n297, A2 => 
                           mult_21_C249_n295, B => mult_21_C249_n296, Z => 
                           mult_21_C249_n294);
   mult_21_C249_U299 : EXOR2D1 port map( A1 => mult_21_C249_n297, A2 => 
                           mult_21_C249_n175, Z => N3364);
   mult_21_C249_U291 : EXNOR2D1 port map( A1 => mult_21_C249_n174, A2 => 
                           mult_21_C249_n294, Z => N3365);
   mult_21_C249_U286 : OAI21D1 port map( A1 => mult_21_C249_n289, A2 => 
                           mult_21_C249_n287, B => mult_21_C249_n288, Z => 
                           mult_21_C249_n286);
   mult_21_C249_U284 : EXOR2D1 port map( A1 => mult_21_C249_n173, A2 => 
                           mult_21_C249_n289, Z => N3366);
   mult_21_C249_U279 : OAI21D1 port map( A1 => mult_21_C249_n285, A2 => 
                           mult_21_C249_n283, B => mult_21_C249_n284, Z => 
                           mult_21_C249_n282);
   mult_21_C249_U278 : EXOR2D1 port map( A1 => mult_21_C249_n172, A2 => 
                           mult_21_C249_n285, Z => N3367);
   mult_21_C249_U273 : OAI21D1 port map( A1 => mult_21_C249_n280, A2 => 
                           mult_21_C249_n284, B => mult_21_C249_n281, Z => 
                           mult_21_C249_n279);
   mult_21_C249_U271 : AOI21D1 port map( A1 => mult_21_C249_n278, A2 => 
                           mult_21_C249_n286, B => mult_21_C249_n279, Z => 
                           mult_21_C249_n277);
   mult_21_C249_U269 : EXNOR2D1 port map( A1 => mult_21_C249_n282, A2 => 
                           mult_21_C249_n171, Z => N3368);
   mult_21_C249_U262 : AOI21D1 port map( A1 => mult_21_C249_n276, A2 => 
                           mult_21_C249_n1529, B => mult_21_C249_n273, Z => 
                           mult_21_C249_n271);
   mult_21_C249_U261 : EXNOR2D1 port map( A1 => mult_21_C249_n276, A2 => 
                           mult_21_C249_n170, Z => N3369);
   mult_21_C249_U254 : AOI21D1 port map( A1 => mult_21_C249_n1526, A2 => 
                           mult_21_C249_n273, B => mult_21_C249_n268, Z => 
                           mult_21_C249_n266);
   mult_21_C249_U252 : OAI21D1 port map( A1 => mult_21_C249_n265, A2 => 
                           mult_21_C249_n277, B => mult_21_C249_n266, Z => 
                           mult_21_C249_n264);
   mult_21_C249_U250 : EXOR2D1 port map( A1 => mult_21_C249_n271, A2 => 
                           mult_21_C249_n169, Z => N3370);
   mult_21_C249_U245 : OAI21D1 port map( A1 => mult_21_C249_n263, A2 => 
                           mult_21_C249_n261, B => mult_21_C249_n262, Z => 
                           mult_21_C249_n260);
   mult_21_C249_U244 : EXOR2D1 port map( A1 => mult_21_C249_n263, A2 => 
                           mult_21_C249_n168, Z => N3371);
   mult_21_C249_U239 : OAI21D1 port map( A1 => mult_21_C249_n258, A2 => 
                           mult_21_C249_n262, B => mult_21_C249_n259, Z => 
                           mult_21_C249_n257);
   mult_21_C249_U237 : AOI21D1 port map( A1 => mult_21_C249_n256, A2 => 
                           mult_21_C249_n264, B => mult_21_C249_n257, Z => 
                           mult_21_C249_n255);
   mult_21_C249_U235 : EXNOR2D1 port map( A1 => mult_21_C249_n260, A2 => 
                           mult_21_C249_n167, Z => N3372);
   mult_21_C249_U228 : AOI21D1 port map( A1 => mult_21_C249_n254, A2 => 
                           mult_21_C249_n1531, B => mult_21_C249_n251, Z => 
                           mult_21_C249_n249);
   mult_21_C249_U227 : EXNOR2D1 port map( A1 => mult_21_C249_n254, A2 => 
                           mult_21_C249_n166, Z => N3373);
   mult_21_C249_U220 : AOI21D1 port map( A1 => mult_21_C249_n1532, A2 => 
                           mult_21_C249_n251, B => mult_21_C249_n246, Z => 
                           mult_21_C249_n244);
   mult_21_C249_U218 : OAI21D1 port map( A1 => mult_21_C249_n255, A2 => 
                           mult_21_C249_n243, B => mult_21_C249_n244, Z => 
                           mult_21_C249_n242);
   mult_21_C249_U216 : EXOR2D1 port map( A1 => mult_21_C249_n249, A2 => 
                           mult_21_C249_n165, Z => N3374);
   mult_21_C249_U211 : OAI21D1 port map( A1 => mult_21_C249_n241, A2 => 
                           mult_21_C249_n239, B => mult_21_C249_n240, Z => 
                           mult_21_C249_n238);
   mult_21_C249_U210 : EXOR2D1 port map( A1 => mult_21_C249_n241, A2 => 
                           mult_21_C249_n164, Z => N3375);
   mult_21_C249_U205 : OAI21D1 port map( A1 => mult_21_C249_n236, A2 => 
                           mult_21_C249_n240, B => mult_21_C249_n237, Z => 
                           mult_21_C249_n235);
   mult_21_C249_U203 : AOI21D1 port map( A1 => mult_21_C249_n242, A2 => 
                           mult_21_C249_n234, B => mult_21_C249_n235, Z => 
                           mult_21_C249_n233);
   mult_21_C249_U201 : EXNOR2D1 port map( A1 => mult_21_C249_n238, A2 => 
                           mult_21_C249_n163, Z => N3376);
   mult_21_C249_U194 : AOI21D1 port map( A1 => mult_21_C249_n232, A2 => 
                           mult_21_C249_n313, B => mult_21_C249_n229, Z => 
                           mult_21_C249_n227);
   mult_21_C249_U193 : EXNOR2D1 port map( A1 => mult_21_C249_n232, A2 => 
                           mult_21_C249_n162, Z => N3377);
   mult_21_C249_U188 : OAI21D1 port map( A1 => mult_21_C249_n225, A2 => 
                           mult_21_C249_n231, B => mult_21_C249_n226, Z => 
                           mult_21_C249_n224);
   mult_21_C249_U186 : AOI21D1 port map( A1 => mult_21_C249_n232, A2 => 
                           mult_21_C249_n223, B => mult_21_C249_n224, Z => 
                           mult_21_C249_n222);
   mult_21_C249_U185 : EXOR2D1 port map( A1 => mult_21_C249_n227, A2 => 
                           mult_21_C249_n161, Z => N3378);
   mult_21_C249_U178 : AOI21D1 port map( A1 => mult_21_C249_n224, A2 => 
                           mult_21_C249_n1530, B => mult_21_C249_n219, Z => 
                           mult_21_C249_n217);
   mult_21_C249_U176 : OAI21D1 port map( A1 => mult_21_C249_n233, A2 => 
                           mult_21_C249_n216, B => mult_21_C249_n217, Z => 
                           mult_21_C249_n215);
   mult_21_C249_U174 : EXOR2D1 port map( A1 => mult_21_C249_n222, A2 => 
                           mult_21_C249_n160, Z => N3379);
   mult_21_C249_U165 : OAI21D1 port map( A1 => mult_21_C249_n214, A2 => 
                           mult_21_C249_n208, B => mult_21_C249_n209, Z => 
                           mult_21_C249_n207);
   mult_21_C249_U164 : EXOR2D1 port map( A1 => mult_21_C249_n214, A2 => 
                           mult_21_C249_n159, Z => N3380);
   mult_21_C249_U157 : AOI21D1 port map( A1 => mult_21_C249_n1527, A2 => 
                           mult_21_C249_n211, B => mult_21_C249_n204, Z => 
                           mult_21_C249_n202);
   mult_21_C249_U155 : OAI21D1 port map( A1 => mult_21_C249_n214, A2 => 
                           mult_21_C249_n201, B => mult_21_C249_n202, Z => 
                           mult_21_C249_n200);
   mult_21_C249_U154 : EXNOR2D1 port map( A1 => mult_21_C249_n207, A2 => 
                           mult_21_C249_n158, Z => N3381);
   mult_21_C249_U147 : AOI21D1 port map( A1 => mult_21_C249_n200, A2 => 
                           mult_21_C249_n1528, B => mult_21_C249_n197, Z => 
                           mult_21_C249_n195);
   mult_21_C249_U146 : EXNOR2D1 port map( A1 => mult_21_C249_n200, A2 => 
                           mult_21_C249_n157, Z => N3382);
   mult_21_C249_U137 : OAI21D1 port map( A1 => mult_21_C249_n202, A2 => 
                           mult_21_C249_n189, B => mult_21_C249_n190, Z => 
                           mult_21_C249_n188);
   mult_21_C249_U134 : EXOR2D1 port map( A1 => mult_21_C249_n195, A2 => 
                           mult_21_C249_n156, Z => N3383);
   mult_21_C249_U132 : ADFULD1 port map( A => mult_21_C249_n531, B => 
                           mult_21_C249_n552, CI => mult_21_C249_n1523, CO => 
                           mult_21_C249_n185, S => N3384);
   mult_21_C249_U131 : ADFULD1 port map( A => mult_21_C249_n507, B => 
                           mult_21_C249_n530, CI => mult_21_C249_n185, CO => 
                           mult_21_C249_n184, S => N3385);
   mult_21_C249_U130 : ADFULD1 port map( A => mult_21_C249_n483, B => 
                           mult_21_C249_n506, CI => mult_21_C249_n184, CO => 
                           mult_21_C249_n183, S => N3386);
   mult_21_C249_U129 : ADFULD1 port map( A => mult_21_C249_n457, B => 
                           mult_21_C249_n482, CI => mult_21_C249_n183, CO => 
                           mult_21_C249_n182, S => N3387);
   mult_21_C249_U128 : ADFULD1 port map( A => mult_21_C249_n431, B => 
                           mult_21_C249_n456, CI => mult_21_C249_n182, CO => 
                           mult_21_C249_n181, S => N3388);
   mult_21_C249_U127 : ADFULD1 port map( A => mult_21_C249_n403, B => 
                           mult_21_C249_n430, CI => mult_21_C249_n181, CO => 
                           mult_21_C249_n180, S => N3389);
   mult_21_C249_U126 : ADFULD1 port map( A => mult_21_C249_n375, B => 
                           mult_21_C249_n402, CI => mult_21_C249_n180, CO => 
                           mult_21_C249_n179, S => N3390);
   mult_21_C249_U125 : ADFULD1 port map( A => mult_21_C249_n345, B => 
                           mult_21_C249_n374, CI => mult_21_C249_n179, CO => 
                           mult_21_C249_n178, S => N3391);

end flat_filter_none_5;
