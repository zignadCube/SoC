-------------------------------------------------------------------------------
-- File         : tvc_forcer_ent.vhd
-- Description  : "forcer" entity to be instantiated in a TVC
-- Author       : Sabih Gerez, University of Twente
-- Creation date: September 1, 2017
-------------------------------------------------------------------------------
-- $Rev: 1$
-- $Author: gerezsh$
-- $Date: Fri Sep  9 19:24:38 CEST 2022$
-- $Log$
-------------------------------------------------------------------------------


entity tvc_forcer is
  port (request_id: in integer);
end tvc_forcer;
