
library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

package CONV_PACK_gp_custom is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_gp_custom;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_gp_custom.all;

architecture hier_filter_none_20 of gp_custom_DW_mult_tc_4 is

   component AOI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component MUXB2DL
      port( A0, A1, SL : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal n42, n50, n58, n66, n73, n80, n84, n89, n94, n99, n104, n156, n157, 
      n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, 
      n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, 
      n182, n183, n184, n185, n186, n202, n203, n204, n205, n206, n207, n208, 
      n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, 
      n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, 
      n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, 
      n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, 
      n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, 
      n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, 
      n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
      n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, 
      n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, 
      n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, 
      n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, 
      n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, 
      n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, 
      n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, 
      n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, 
      n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, 
      n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, 
      n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, 
      n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, 
      n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, 
      n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, 
      n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, 
      n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, 
      n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, 
      n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, 
      n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, 
      n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
      n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, 
      n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, 
      n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, 
      n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
      n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, 
      n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, 
      n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, 
      n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, 
      n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, 
      n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, 
      n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, 
      n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, 
      n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, 
      n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, 
      n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, 
      n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, 
      n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, 
      n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, 
      n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, 
      n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, 
      n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, 
      n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, 
      n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, 
      n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, 
      n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, 
      n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, 
      n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, 
      n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, 
      n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, 
      n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, 
      n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, 
      n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, 
      n917, n918, n919, n920, n921, n922, n923, n939, n940, n941, n942, n943, 
      n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n955, n956, 
      n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, 
      n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, 
      n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, 
      n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, 
      n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, 
      n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, 
      n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, 
      n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, 
      n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, 
      n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, 
      n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, 
      n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, 
      n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, 
      n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, 
      n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, 
      n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, 
      n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, 
      n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, 
      n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, 
      n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, 
      n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, 
      n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, 
      n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, 
      n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, 
      n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, 
      n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, 
      n1224, n1225, n1226, n1375, n1376, n1377, n1378, n1379, n1380, n1381, 
      n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, 
      n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, 
      n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, 
      n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, 
      n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, 
      n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, 
      n1442, n1443, n1444, n1445, n1446, n1447, n1448 : std_logic;

begin
   
   U125 : ADFULD1 port map( A => n203, B => n232, CI => n157, CO => n156, S => 
                           product(30));
   U126 : ADFULD1 port map( A => n233, B => n260, CI => n158, CO => n157, S => 
                           product(29));
   U127 : ADFULD1 port map( A => n261, B => n288, CI => n159, CO => n158, S => 
                           product(28));
   U128 : ADFULD1 port map( A => n289, B => n314, CI => n160, CO => n159, S => 
                           product(27));
   U129 : ADFULD1 port map( A => n315, B => n340, CI => n161, CO => n160, S => 
                           product(26));
   U130 : ADFULD1 port map( A => n341, B => n364, CI => n162, CO => n161, S => 
                           product(25));
   U131 : ADFULD1 port map( A => n365, B => n388, CI => n163, CO => n162, S => 
                           product(24));
   U132 : ADFULD1 port map( A => n389, B => n410, CI => n164, CO => n163, S => 
                           product(23));
   U133 : ADFULD1 port map( A => n411, B => n432, CI => n165, CO => n164, S => 
                           product(22));
   U134 : ADFULD1 port map( A => n433, B => n452, CI => n166, CO => n165, S => 
                           product(21));
   U135 : ADFULD1 port map( A => n453, B => n472, CI => n167, CO => n166, S => 
                           product(20));
   U136 : ADFULD1 port map( A => n473, B => n490, CI => n168, CO => n167, S => 
                           product(19));
   U137 : ADFULD1 port map( A => n491, B => n508, CI => n169, CO => n168, S => 
                           product(18));
   U138 : ADFULD1 port map( A => n509, B => n524, CI => n170, CO => n169, S => 
                           product(17));
   U139 : ADFULD1 port map( A => n525, B => n540, CI => n171, CO => n170, S => 
                           product(16));
   U140 : ADFULD1 port map( A => n541, B => n554, CI => n172, CO => n171, S => 
                           product(15));
   U141 : ADFULD1 port map( A => n555, B => n568, CI => n173, CO => n172, S => 
                           product(14));
   U142 : ADFULD1 port map( A => n569, B => n580, CI => n174, CO => n173, S => 
                           product(13));
   U143 : ADFULD1 port map( A => n581, B => n592, CI => n175, CO => n174, S => 
                           product(12));
   U144 : ADFULD1 port map( A => n593, B => n602, CI => n176, CO => n175, S => 
                           product(11));
   U145 : ADFULD1 port map( A => n603, B => n612, CI => n177, CO => n176, S => 
                           product(10));
   U146 : ADFULD1 port map( A => n613, B => n620, CI => n178, CO => n177, S => 
                           product(9));
   U147 : ADFULD1 port map( A => n621, B => n628, CI => n179, CO => n178, S => 
                           product(8));
   U148 : ADFULD1 port map( A => n629, B => n634, CI => n180, CO => n179, S => 
                           product(7));
   U149 : ADFULD1 port map( A => n635, B => n640, CI => n181, CO => n180, S => 
                           product(6));
   U150 : ADFULD1 port map( A => n641, B => n644, CI => n182, CO => n181, S => 
                           product(5));
   U151 : ADFULD1 port map( A => n645, B => n648, CI => n183, CO => n182, S => 
                           product(4));
   U152 : ADFULD1 port map( A => n649, B => n1193, CI => n184, CO => n183, S =>
                           product(3));
   U153 : ADFULD1 port map( A => n651, B => n1194, CI => n185, CO => n184, S =>
                           product(2));
   U154 : ADHALFDL port map( A => n186, B => n1225, CO => n185, S => product(1)
                           );
   U155 : ADHALFDL port map( A => n1226, B => a(1), CO => n186, S => product(0)
                           );
   U171 : ADFULD1 port map( A => n234, B => n207, CI => n205, CO => n202, S => 
                           n203);
   U172 : ADFULD1 port map( A => n209, B => n211, CI => n236, CO => n204, S => 
                           n205);
   U173 : ADFULD1 port map( A => n240, B => n213, CI => n238, CO => n206, S => 
                           n207);
   U174 : ADFULD1 port map( A => n217, B => n242, CI => n215, CO => n208, S => 
                           n209);
   U175 : ADFULD1 port map( A => n244, B => n246, CI => n219, CO => n210, S => 
                           n211);
   U176 : ADFULD1 port map( A => n225, B => n223, CI => n248, CO => n212, S => 
                           n213);
   U177 : ADFULD1 port map( A => n221, B => n229, CI => n227, CO => n214, S => 
                           n215);
   U178 : ADFULD1 port map( A => n256, B => n252, CI => n254, CO => n216, S => 
                           n217);
   U179 : ADFULD1 port map( A => n258, B => n1088, CI => n250, CO => n218, S =>
                           n219);
   U180 : ADFULD1 port map( A => n1046, B => n1112, CI => n1066, CO => n220, S 
                           => n221);
   U181 : ADFULD1 port map( A => n986, B => n976, CI => n998, CO => n222, S => 
                           n223);
   U182 : ADFULD1 port map( A => n962, B => n1138, CI => n968, CO => n224, S =>
                           n225);
   U183 : ADFULD1 port map( A => n1166, B => n1012, CI => n231, CO => n226, S 
                           => n227);
   U184 : ADFULD1 port map( A => n1028, B => n956, CI => n958, CO => n228, S =>
                           n229);
   U185 : ADHALFDL port map( A => n1196, B => n939, CO => n230, S => n231);
   U186 : ADFULD1 port map( A => n262, B => n237, CI => n235, CO => n232, S => 
                           n233);
   U187 : ADFULD1 port map( A => n239, B => n266, CI => n264, CO => n234, S => 
                           n235);
   U188 : ADFULD1 port map( A => n268, B => n243, CI => n241, CO => n236, S => 
                           n237);
   U189 : ADFULD1 port map( A => n270, B => n247, CI => n245, CO => n238, S => 
                           n239);
   U190 : ADFULD1 port map( A => n274, B => n249, CI => n272, CO => n240, S => 
                           n241);
   U191 : ADFULD1 port map( A => n253, B => n255, CI => n257, CO => n242, S => 
                           n243);
   U192 : ADFULD1 port map( A => n280, B => n276, CI => n251, CO => n244, S => 
                           n245);
   U193 : ADFULD1 port map( A => n278, B => n284, CI => n282, CO => n246, S => 
                           n247);
   U194 : ADFULD1 port map( A => n1047, B => n1013, CI => n259, CO => n248, S 
                           => n249);
   U195 : ADFULD1 port map( A => n977, B => n1067, CI => n999, CO => n250, S =>
                           n251);
   U196 : ADFULD1 port map( A => n959, B => n969, CI => n963, CO => n252, S => 
                           n253);
   U197 : ADFULD1 port map( A => n1113, B => n987, CI => n1089, CO => n254, S 
                           => n255);
   U198 : ADFULD1 port map( A => n1167, B => n1029, CI => n1139, CO => n256, S 
                           => n257);
   U199 : ADHALFDL port map( A => n286, B => n1197, CO => n258, S => n259);
   U200 : ADFULD1 port map( A => n290, B => n265, CI => n263, CO => n260, S => 
                           n261);
   U201 : ADFULD1 port map( A => n267, B => n294, CI => n292, CO => n262, S => 
                           n263);
   U202 : ADFULD1 port map( A => n296, B => n271, CI => n269, CO => n264, S => 
                           n265);
   U203 : ADFULD1 port map( A => n275, B => n298, CI => n273, CO => n266, S => 
                           n267);
   U204 : ADFULD1 port map( A => n302, B => n281, CI => n300, CO => n268, S => 
                           n269);
   U205 : ADFULD1 port map( A => n283, B => n277, CI => n279, CO => n270, S => 
                           n271);
   U206 : ADFULD1 port map( A => n310, B => n308, CI => n285, CO => n272, S => 
                           n273);
   U207 : ADFULD1 port map( A => n304, B => n312, CI => n306, CO => n274, S => 
                           n275);
   U208 : ADFULD1 port map( A => n1014, B => n1068, CI => n1048, CO => n276, S 
                           => n277);
   U209 : ADFULD1 port map( A => n978, B => n1090, CI => n988, CO => n278, S =>
                           n279);
   U210 : ADFULD1 port map( A => n964, B => n1114, CI => n970, CO => n280, S =>
                           n281);
   U211 : ADFULD1 port map( A => n1140, B => n1000, CI => n287, CO => n282, S 
                           => n283);
   U212 : ADFULD1 port map( A => n1030, B => n960, CI => n1168, CO => n284, S 
                           => n285);
   U213 : ADHALFDL port map( A => n1198, B => n940, CO => n286, S => n287);
   U214 : ADFULD1 port map( A => n316, B => n293, CI => n291, CO => n288, S => 
                           n289);
   U215 : ADFULD1 port map( A => n318, B => n297, CI => n295, CO => n290, S => 
                           n291);
   U216 : ADFULD1 port map( A => n299, B => n322, CI => n320, CO => n292, S => 
                           n293);
   U217 : ADFULD1 port map( A => n324, B => n303, CI => n301, CO => n294, S => 
                           n295);
   U218 : ADFULD1 port map( A => n307, B => n309, CI => n326, CO => n296, S => 
                           n297);
   U219 : ADFULD1 port map( A => n305, B => n328, CI => n311, CO => n298, S => 
                           n299);
   U220 : ADFULD1 port map( A => n332, B => n330, CI => n334, CO => n300, S => 
                           n301);
   U221 : ADFULD1 port map( A => n313, B => n1091, CI => n336, CO => n302, S =>
                           n303);
   U222 : ADFULD1 port map( A => n1015, B => n1115, CI => n1069, CO => n304, S 
                           => n305);
   U223 : ADFULD1 port map( A => n1141, B => n1001, CI => n989, CO => n306, S 
                           => n307);
   U224 : ADFULD1 port map( A => n979, B => n1049, CI => n1169, CO => n308, S 
                           => n309);
   U225 : ADFULD1 port map( A => n965, B => n1031, CI => n971, CO => n310, S =>
                           n311);
   U226 : ADHALFDL port map( A => n338, B => n1199, CO => n312, S => n313);
   U227 : ADFULD1 port map( A => n342, B => n319, CI => n317, CO => n314, S => 
                           n315);
   U228 : ADFULD1 port map( A => n344, B => n346, CI => n321, CO => n316, S => 
                           n317);
   U229 : ADFULD1 port map( A => n325, B => n327, CI => n323, CO => n318, S => 
                           n319);
   U230 : ADFULD1 port map( A => n350, B => n352, CI => n348, CO => n320, S => 
                           n321);
   U231 : ADFULD1 port map( A => n333, B => n335, CI => n329, CO => n322, S => 
                           n323);
   U232 : ADFULD1 port map( A => n337, B => n358, CI => n331, CO => n324, S => 
                           n325);
   U233 : ADFULD1 port map( A => n354, B => n360, CI => n356, CO => n326, S => 
                           n327);
   U234 : ADFULD1 port map( A => n1092, B => n1116, CI => n362, CO => n328, S 
                           => n329);
   U235 : ADFULD1 port map( A => n1016, B => n1142, CI => n1070, CO => n330, S 
                           => n331);
   U236 : ADFULD1 port map( A => n990, B => n1170, CI => n1002, CO => n332, S 
                           => n333);
   U237 : ADFULD1 port map( A => n980, B => n1032, CI => n339, CO => n334, S =>
                           n335);
   U238 : ADFULD1 port map( A => n1050, B => n966, CI => n972, CO => n336, S =>
                           n337);
   U239 : ADHALFDL port map( A => n1200, B => n941, CO => n338, S => n339);
   U240 : ADFULD1 port map( A => n366, B => n345, CI => n343, CO => n340, S => 
                           n341);
   U241 : ADFULD1 port map( A => n347, B => n370, CI => n368, CO => n342, S => 
                           n343);
   U242 : ADFULD1 port map( A => n351, B => n372, CI => n349, CO => n344, S => 
                           n345);
   U243 : ADFULD1 port map( A => n374, B => n376, CI => n353, CO => n346, S => 
                           n347);
   U244 : ADFULD1 port map( A => n361, B => n357, CI => n359, CO => n348, S => 
                           n349);
   U245 : ADFULD1 port map( A => n378, B => n380, CI => n355, CO => n350, S => 
                           n351);
   U246 : ADFULD1 port map( A => n384, B => n363, CI => n382, CO => n352, S => 
                           n353);
   U247 : ADFULD1 port map( A => n1033, B => n1093, CI => n1071, CO => n354, S 
                           => n355);
   U248 : ADFULD1 port map( A => n991, B => n1117, CI => n1017, CO => n356, S 
                           => n357);
   U249 : ADFULD1 port map( A => n973, B => n1003, CI => n981, CO => n358, S =>
                           n359);
   U250 : ADFULD1 port map( A => n1171, B => n1051, CI => n1143, CO => n360, S 
                           => n361);
   U251 : ADHALFDL port map( A => n386, B => n1201, CO => n362, S => n363);
   U252 : ADFULD1 port map( A => n390, B => n369, CI => n367, CO => n364, S => 
                           n365);
   U253 : ADFULD1 port map( A => n371, B => n394, CI => n392, CO => n366, S => 
                           n367);
   U254 : ADFULD1 port map( A => n375, B => n396, CI => n373, CO => n368, S => 
                           n369);
   U255 : ADFULD1 port map( A => n398, B => n400, CI => n377, CO => n370, S => 
                           n371);
   U256 : ADFULD1 port map( A => n383, B => n379, CI => n381, CO => n372, S => 
                           n373);
   U257 : ADFULD1 port map( A => n402, B => n404, CI => n385, CO => n374, S => 
                           n375);
   U258 : ADFULD1 port map( A => n408, B => n1072, CI => n406, CO => n376, S =>
                           n377);
   U259 : ADFULD1 port map( A => n1004, B => n1094, CI => n1034, CO => n378, S 
                           => n379);
   U260 : ADFULD1 port map( A => n992, B => n1144, CI => n1118, CO => n380, S 
                           => n381);
   U261 : ADFULD1 port map( A => n982, B => n1018, CI => n387, CO => n382, S =>
                           n383);
   U262 : ADFULD1 port map( A => n1052, B => n974, CI => n1172, CO => n384, S 
                           => n385);
   U263 : ADHALFDL port map( A => n1202, B => n942, CO => n386, S => n387);
   U264 : ADFULD1 port map( A => n412, B => n393, CI => n391, CO => n388, S => 
                           n389);
   U265 : ADFULD1 port map( A => n395, B => n397, CI => n414, CO => n390, S => 
                           n391);
   U266 : ADFULD1 port map( A => n399, B => n418, CI => n416, CO => n392, S => 
                           n393);
   U267 : ADFULD1 port map( A => n401, B => n407, CI => n420, CO => n394, S => 
                           n395);
   U268 : ADFULD1 port map( A => n403, B => n424, CI => n405, CO => n396, S => 
                           n397);
   U269 : ADFULD1 port map( A => n426, B => n428, CI => n422, CO => n398, S => 
                           n399);
   U270 : ADFULD1 port map( A => n1073, B => n1095, CI => n409, CO => n400, S 
                           => n401);
   U271 : ADFULD1 port map( A => n1005, B => n1119, CI => n1019, CO => n402, S 
                           => n403);
   U272 : ADFULD1 port map( A => n1173, B => n1035, CI => n1145, CO => n404, S 
                           => n405);
   U273 : ADFULD1 port map( A => n983, B => n1053, CI => n993, CO => n406, S =>
                           n407);
   U274 : ADHALFDL port map( A => n430, B => n1203, CO => n408, S => n409);
   U275 : ADFULD1 port map( A => n434, B => n415, CI => n413, CO => n410, S => 
                           n411);
   U276 : ADFULD1 port map( A => n417, B => n419, CI => n436, CO => n412, S => 
                           n413);
   U277 : ADFULD1 port map( A => n421, B => n440, CI => n438, CO => n414, S => 
                           n415);
   U278 : ADFULD1 port map( A => n427, B => n425, CI => n442, CO => n416, S => 
                           n417);
   U279 : ADFULD1 port map( A => n429, B => n444, CI => n423, CO => n418, S => 
                           n419);
   U280 : ADFULD1 port map( A => n448, B => n450, CI => n446, CO => n420, S => 
                           n421);
   U281 : ADFULD1 port map( A => n1074, B => n1120, CI => n1096, CO => n422, S 
                           => n423);
   U282 : ADFULD1 port map( A => n1006, B => n1146, CI => n1020, CO => n424, S 
                           => n425);
   U283 : ADFULD1 port map( A => n1174, B => n1036, CI => n431, CO => n426, S 
                           => n427);
   U284 : ADFULD1 port map( A => n1054, B => n984, CI => n994, CO => n428, S =>
                           n429);
   U285 : ADHALFDL port map( A => n1204, B => n943, CO => n430, S => n431);
   U286 : ADFULD1 port map( A => n454, B => n437, CI => n435, CO => n432, S => 
                           n433);
   U287 : ADFULD1 port map( A => n439, B => n441, CI => n456, CO => n434, S => 
                           n435);
   U288 : ADFULD1 port map( A => n443, B => n460, CI => n458, CO => n436, S => 
                           n437);
   U289 : ADFULD1 port map( A => n449, B => n445, CI => n447, CO => n438, S => 
                           n439);
   U290 : ADFULD1 port map( A => n464, B => n466, CI => n462, CO => n440, S => 
                           n441);
   U291 : ADFULD1 port map( A => n451, B => n1037, CI => n468, CO => n442, S =>
                           n443);
   U292 : ADFULD1 port map( A => n995, B => n1075, CI => n1007, CO => n444, S 
                           => n445);
   U293 : ADFULD1 port map( A => n1121, B => n1021, CI => n1097, CO => n446, S 
                           => n447);
   U294 : ADFULD1 port map( A => n1175, B => n1055, CI => n1147, CO => n448, S 
                           => n449);
   U295 : ADHALFDL port map( A => n470, B => n1205, CO => n450, S => n451);
   U296 : ADFULD1 port map( A => n474, B => n457, CI => n455, CO => n452, S => 
                           n453);
   U297 : ADFULD1 port map( A => n459, B => n461, CI => n476, CO => n454, S => 
                           n455);
   U298 : ADFULD1 port map( A => n480, B => n463, CI => n478, CO => n456, S => 
                           n457);
   U299 : ADFULD1 port map( A => n465, B => n469, CI => n467, CO => n458, S => 
                           n459);
   U300 : ADFULD1 port map( A => n482, B => n486, CI => n484, CO => n460, S => 
                           n461);
   U301 : ADFULD1 port map( A => n1098, B => n1122, CI => n488, CO => n462, S 
                           => n463);
   U302 : ADFULD1 port map( A => n1022, B => n1148, CI => n1056, CO => n464, S 
                           => n465);
   U303 : ADFULD1 port map( A => n1008, B => n1038, CI => n471, CO => n466, S 
                           => n467);
   U304 : ADFULD1 port map( A => n1076, B => n996, CI => n1176, CO => n468, S 
                           => n469);
   U305 : ADHALFDL port map( A => n1206, B => n944, CO => n470, S => n471);
   U306 : ADFULD1 port map( A => n492, B => n477, CI => n475, CO => n472, S => 
                           n473);
   U307 : ADFULD1 port map( A => n479, B => n481, CI => n494, CO => n474, S => 
                           n475);
   U308 : ADFULD1 port map( A => n498, B => n487, CI => n496, CO => n476, S => 
                           n477);
   U309 : ADFULD1 port map( A => n483, B => n500, CI => n485, CO => n478, S => 
                           n479);
   U310 : ADFULD1 port map( A => n504, B => n489, CI => n502, CO => n480, S => 
                           n481);
   U311 : ADFULD1 port map( A => n1057, B => n1149, CI => n1123, CO => n482, S 
                           => n483);
   U312 : ADFULD1 port map( A => n1177, B => n1099, CI => n1039, CO => n484, S 
                           => n485);
   U313 : ADFULD1 port map( A => n1009, B => n1077, CI => n1023, CO => n486, S 
                           => n487);
   U314 : ADHALFDL port map( A => n506, B => n1207, CO => n488, S => n489);
   U315 : ADFULD1 port map( A => n510, B => n495, CI => n493, CO => n490, S => 
                           n491);
   U316 : ADFULD1 port map( A => n497, B => n499, CI => n512, CO => n492, S => 
                           n493);
   U317 : ADFULD1 port map( A => n516, B => n503, CI => n514, CO => n494, S => 
                           n495);
   U318 : ADFULD1 port map( A => n505, B => n518, CI => n501, CO => n496, S => 
                           n497);
   U319 : ADFULD1 port map( A => n522, B => n1124, CI => n520, CO => n498, S =>
                           n499);
   U320 : ADFULD1 port map( A => n1040, B => n1150, CI => n1058, CO => n500, S 
                           => n501);
   U321 : ADFULD1 port map( A => n1178, B => n1100, CI => n507, CO => n502, S 
                           => n503);
   U322 : ADFULD1 port map( A => n1078, B => n1010, CI => n1024, CO => n504, S 
                           => n505);
   U323 : ADHALFDL port map( A => n1208, B => n945, CO => n506, S => n507);
   U324 : ADFULD1 port map( A => n526, B => n513, CI => n511, CO => n508, S => 
                           n509);
   U325 : ADFULD1 port map( A => n528, B => n530, CI => n515, CO => n510, S => 
                           n511);
   U326 : ADFULD1 port map( A => n521, B => n519, CI => n517, CO => n512, S => 
                           n513);
   U327 : ADFULD1 port map( A => n534, B => n536, CI => n532, CO => n514, S => 
                           n515);
   U328 : ADFULD1 port map( A => n1101, B => n1125, CI => n523, CO => n516, S 
                           => n517);
   U329 : ADFULD1 port map( A => n1025, B => n1041, CI => n1059, CO => n518, S 
                           => n519);
   U330 : ADFULD1 port map( A => n1179, B => n1079, CI => n1151, CO => n520, S 
                           => n521);
   U331 : ADHALFDL port map( A => n538, B => n1209, CO => n522, S => n523);
   U332 : ADFULD1 port map( A => n542, B => n529, CI => n527, CO => n524, S => 
                           n525);
   U333 : ADFULD1 port map( A => n544, B => n546, CI => n531, CO => n526, S => 
                           n527);
   U334 : ADFULD1 port map( A => n533, B => n537, CI => n535, CO => n528, S => 
                           n529);
   U335 : ADFULD1 port map( A => n550, B => n552, CI => n548, CO => n530, S => 
                           n531);
   U336 : ADFULD1 port map( A => n1080, B => n1152, CI => n1126, CO => n532, S 
                           => n533);
   U337 : ADFULD1 port map( A => n1042, B => n1060, CI => n539, CO => n534, S 
                           => n535);
   U338 : ADFULD1 port map( A => n1102, B => n1026, CI => n1180, CO => n536, S 
                           => n537);
   U339 : ADHALFDL port map( A => n1210, B => n946, CO => n538, S => n539);
   U340 : ADFULD1 port map( A => n556, B => n545, CI => n543, CO => n540, S => 
                           n541);
   U341 : ADFULD1 port map( A => n547, B => n551, CI => n558, CO => n542, S => 
                           n543);
   U342 : ADFULD1 port map( A => n560, B => n562, CI => n549, CO => n544, S => 
                           n545);
   U343 : ADFULD1 port map( A => n553, B => n1153, CI => n564, CO => n546, S =>
                           n547);
   U344 : ADFULD1 port map( A => n1181, B => n1081, CI => n1127, CO => n548, S 
                           => n549);
   U345 : ADFULD1 port map( A => n1043, B => n1103, CI => n1061, CO => n550, S 
                           => n551);
   U346 : ADHALFDL port map( A => n566, B => n1211, CO => n552, S => n553);
   U347 : ADFULD1 port map( A => n570, B => n559, CI => n557, CO => n554, S => 
                           n555);
   U348 : ADFULD1 port map( A => n561, B => n563, CI => n572, CO => n556, S => 
                           n557);
   U349 : ADFULD1 port map( A => n574, B => n576, CI => n565, CO => n558, S => 
                           n559);
   U350 : ADFULD1 port map( A => n1062, B => n1128, CI => n578, CO => n560, S 
                           => n561);
   U351 : ADFULD1 port map( A => n1154, B => n1082, CI => n567, CO => n562, S 
                           => n563);
   U352 : ADFULD1 port map( A => n1104, B => n1044, CI => n1182, CO => n564, S 
                           => n565);
   U353 : ADHALFDL port map( A => n1212, B => n947, CO => n566, S => n567);
   U354 : ADFULD1 port map( A => n582, B => n573, CI => n571, CO => n568, S => 
                           n569);
   U355 : ADFULD1 port map( A => n577, B => n575, CI => n584, CO => n570, S => 
                           n571);
   U356 : ADFULD1 port map( A => n588, B => n579, CI => n586, CO => n572, S => 
                           n573);
   U357 : ADFULD1 port map( A => n1063, B => n1129, CI => n1083, CO => n574, S 
                           => n575);
   U358 : ADFULD1 port map( A => n1183, B => n1105, CI => n1155, CO => n576, S 
                           => n577);
   U359 : ADHALFDL port map( A => n590, B => n1213, CO => n578, S => n579);
   U360 : ADFULD1 port map( A => n585, B => n594, CI => n583, CO => n580, S => 
                           n581);
   U361 : ADFULD1 port map( A => n587, B => n589, CI => n596, CO => n582, S => 
                           n583);
   U362 : ADFULD1 port map( A => n600, B => n1106, CI => n598, CO => n584, S =>
                           n585);
   U363 : ADFULD1 port map( A => n1084, B => n1156, CI => n591, CO => n586, S 
                           => n587);
   U364 : ADFULD1 port map( A => n1130, B => n1064, CI => n1184, CO => n588, S 
                           => n589);
   U365 : ADHALFDL port map( A => n1214, B => n948, CO => n590, S => n591);
   U366 : ADFULD1 port map( A => n604, B => n597, CI => n595, CO => n592, S => 
                           n593);
   U367 : ADFULD1 port map( A => n606, B => n608, CI => n599, CO => n594, S => 
                           n595);
   U368 : ADFULD1 port map( A => n1107, B => n1157, CI => n601, CO => n596, S 
                           => n597);
   U369 : ADFULD1 port map( A => n1085, B => n1131, CI => n1185, CO => n598, S 
                           => n599);
   U370 : ADHALFDL port map( A => n610, B => n1215, CO => n600, S => n601);
   U371 : ADFULD1 port map( A => n614, B => n607, CI => n605, CO => n602, S => 
                           n603);
   U372 : ADFULD1 port map( A => n616, B => n618, CI => n609, CO => n604, S => 
                           n605);
   U373 : ADFULD1 port map( A => n1108, B => n1158, CI => n611, CO => n606, S 
                           => n607);
   U374 : ADFULD1 port map( A => n1132, B => n1086, CI => n1186, CO => n608, S 
                           => n609);
   U375 : ADHALFDL port map( A => n1216, B => n949, CO => n610, S => n611);
   U376 : ADFULD1 port map( A => n617, B => n622, CI => n615, CO => n612, S => 
                           n613);
   U377 : ADFULD1 port map( A => n619, B => n1187, CI => n624, CO => n614, S =>
                           n615);
   U378 : ADFULD1 port map( A => n1109, B => n1133, CI => n1159, CO => n616, S 
                           => n617);
   U379 : ADHALFDL port map( A => n626, B => n1217, CO => n618, S => n619);
   U380 : ADFULD1 port map( A => n625, B => n630, CI => n623, CO => n620, S => 
                           n621);
   U381 : ADFULD1 port map( A => n627, B => n1160, CI => n632, CO => n622, S =>
                           n623);
   U382 : ADFULD1 port map( A => n1188, B => n1110, CI => n1134, CO => n624, S 
                           => n625);
   U383 : ADHALFDL port map( A => n1218, B => n950, CO => n626, S => n627);
   U384 : ADFULD1 port map( A => n636, B => n633, CI => n631, CO => n628, S => 
                           n629);
   U385 : ADFULD1 port map( A => n1135, B => n1189, CI => n1161, CO => n630, S 
                           => n631);
   U386 : ADHALFDL port map( A => n638, B => n1219, CO => n632, S => n633);
   U387 : ADFULD1 port map( A => n642, B => n639, CI => n637, CO => n634, S => 
                           n635);
   U388 : ADFULD1 port map( A => n1190, B => n1136, CI => n1162, CO => n636, S 
                           => n637);
   U389 : ADHALFDL port map( A => n1220, B => n951, CO => n638, S => n639);
   U390 : ADFULD1 port map( A => n1163, B => n1191, CI => n643, CO => n640, S 
                           => n641);
   U391 : ADHALFDL port map( A => n646, B => n1221, CO => n642, S => n643);
   U392 : ADFULD1 port map( A => n1192, B => n1164, CI => n647, CO => n644, S 
                           => n645);
   U393 : ADHALFDL port map( A => n1222, B => n952, CO => n646, S => n647);
   U394 : ADHALFDL port map( A => n650, B => n1223, CO => n648, S => n649);
   U395 : ADHALFDL port map( A => n1224, B => n953, CO => n650, S => n651);
   U397 : MUXB2DL port map( A0 => n104, A1 => n1417, SL => n652, Z => n955);
   U399 : MUXB2DL port map( A0 => n104, A1 => n1417, SL => n653, Z => n956);
   U402 : MUXB2DL port map( A0 => n99, A1 => n1416, SL => n654, Z => n957);
   U404 : MUXB2DL port map( A0 => n99, A1 => n1416, SL => n655, Z => n958);
   U406 : MUXB2DL port map( A0 => n99, A1 => n1416, SL => n656, Z => n959);
   U408 : MUXB2DL port map( A0 => n99, A1 => n1416, SL => n657, Z => n960);
   U411 : MUXB2DL port map( A0 => n94, A1 => n1413, SL => n658, Z => n961);
   U413 : MUXB2DL port map( A0 => n94, A1 => n1413, SL => n659, Z => n962);
   U415 : MUXB2DL port map( A0 => n94, A1 => n1413, SL => n660, Z => n963);
   U417 : MUXB2DL port map( A0 => n94, A1 => n1413, SL => n661, Z => n964);
   U419 : MUXB2DL port map( A0 => n94, A1 => n1413, SL => n662, Z => n965);
   U421 : MUXB2DL port map( A0 => n94, A1 => n1413, SL => n663, Z => n966);
   U424 : MUXB2DL port map( A0 => n89, A1 => n1411, SL => n664, Z => n967);
   U426 : MUXB2DL port map( A0 => n89, A1 => n1411, SL => n665, Z => n968);
   U428 : MUXB2DL port map( A0 => n89, A1 => n1411, SL => n666, Z => n969);
   U430 : MUXB2DL port map( A0 => n89, A1 => n1411, SL => n667, Z => n970);
   U432 : MUXB2DL port map( A0 => n89, A1 => n1411, SL => n668, Z => n971);
   U434 : MUXB2DL port map( A0 => n89, A1 => n1411, SL => n669, Z => n972);
   U436 : MUXB2DL port map( A0 => n89, A1 => n1411, SL => n670, Z => n973);
   U438 : MUXB2DL port map( A0 => n89, A1 => n1411, SL => n671, Z => n974);
   U441 : MUXB2DL port map( A0 => n84, A1 => n1409, SL => n672, Z => n975);
   U443 : MUXB2DL port map( A0 => n84, A1 => n1409, SL => n673, Z => n976);
   U445 : MUXB2DL port map( A0 => n84, A1 => n1409, SL => n674, Z => n977);
   U447 : MUXB2DL port map( A0 => n84, A1 => n1409, SL => n675, Z => n978);
   U449 : MUXB2DL port map( A0 => n84, A1 => n1409, SL => n676, Z => n979);
   U451 : MUXB2DL port map( A0 => n84, A1 => n1409, SL => n677, Z => n980);
   U453 : MUXB2DL port map( A0 => n84, A1 => n1409, SL => n678, Z => n981);
   U455 : MUXB2DL port map( A0 => n84, A1 => n1409, SL => n679, Z => n982);
   U457 : MUXB2DL port map( A0 => n84, A1 => n1409, SL => n680, Z => n983);
   U459 : MUXB2DL port map( A0 => n84, A1 => n1409, SL => n681, Z => n984);
   U462 : MUXB2DL port map( A0 => n80, A1 => n1407, SL => n682, Z => n985);
   U464 : MUXB2DL port map( A0 => n80, A1 => n1407, SL => n683, Z => n986);
   U466 : MUXB2DL port map( A0 => n80, A1 => n1407, SL => n684, Z => n987);
   U468 : MUXB2DL port map( A0 => n80, A1 => n1407, SL => n685, Z => n988);
   U470 : MUXB2DL port map( A0 => n80, A1 => n1407, SL => n686, Z => n989);
   U472 : MUXB2DL port map( A0 => n80, A1 => n1407, SL => n687, Z => n990);
   U474 : MUXB2DL port map( A0 => n80, A1 => n1407, SL => n688, Z => n991);
   U476 : MUXB2DL port map( A0 => n80, A1 => n1407, SL => n689, Z => n992);
   U478 : MUXB2DL port map( A0 => n80, A1 => n1407, SL => n690, Z => n993);
   U480 : MUXB2DL port map( A0 => n80, A1 => n1407, SL => n691, Z => n994);
   U482 : MUXB2DL port map( A0 => n80, A1 => n1407, SL => n692, Z => n995);
   U484 : MUXB2DL port map( A0 => n80, A1 => n1407, SL => n693, Z => n996);
   U487 : MUXB2DL port map( A0 => n73, A1 => n1405, SL => n694, Z => n997);
   U489 : MUXB2DL port map( A0 => n73, A1 => n1405, SL => n695, Z => n998);
   U491 : MUXB2DL port map( A0 => n73, A1 => n1405, SL => n696, Z => n999);
   U493 : MUXB2DL port map( A0 => n73, A1 => n1405, SL => n697, Z => n1000);
   U495 : MUXB2DL port map( A0 => n73, A1 => n1405, SL => n698, Z => n1001);
   U497 : MUXB2DL port map( A0 => n73, A1 => n1405, SL => n699, Z => n1002);
   U499 : MUXB2DL port map( A0 => n73, A1 => n1405, SL => n700, Z => n1003);
   U501 : MUXB2DL port map( A0 => n73, A1 => n1405, SL => n701, Z => n1004);
   U503 : MUXB2DL port map( A0 => n73, A1 => n1405, SL => n702, Z => n1005);
   U505 : MUXB2DL port map( A0 => n73, A1 => n1405, SL => n703, Z => n1006);
   U507 : MUXB2DL port map( A0 => n73, A1 => n1405, SL => n704, Z => n1007);
   U509 : MUXB2DL port map( A0 => n73, A1 => n1405, SL => n705, Z => n1008);
   U511 : MUXB2DL port map( A0 => n73, A1 => n1405, SL => n706, Z => n1009);
   U513 : MUXB2DL port map( A0 => n73, A1 => n1405, SL => n707, Z => n1010);
   U516 : MUXB2DL port map( A0 => n66, A1 => n1403, SL => n708, Z => n1011);
   U518 : MUXB2DL port map( A0 => n66, A1 => n1403, SL => n709, Z => n1012);
   U520 : MUXB2DL port map( A0 => n66, A1 => n1403, SL => n710, Z => n1013);
   U522 : MUXB2DL port map( A0 => n66, A1 => n1403, SL => n711, Z => n1014);
   U524 : MUXB2DL port map( A0 => n66, A1 => n1403, SL => n712, Z => n1015);
   U526 : MUXB2DL port map( A0 => n66, A1 => n1403, SL => n713, Z => n1016);
   U528 : MUXB2DL port map( A0 => n66, A1 => n1403, SL => n714, Z => n1017);
   U530 : MUXB2DL port map( A0 => n66, A1 => n1403, SL => n715, Z => n1018);
   U532 : MUXB2DL port map( A0 => n66, A1 => n1403, SL => n716, Z => n1019);
   U534 : MUXB2DL port map( A0 => n66, A1 => n1403, SL => n717, Z => n1020);
   U536 : MUXB2DL port map( A0 => n66, A1 => n1403, SL => n718, Z => n1021);
   U538 : MUXB2DL port map( A0 => n66, A1 => n1403, SL => n719, Z => n1022);
   U540 : MUXB2DL port map( A0 => n66, A1 => n1403, SL => n720, Z => n1023);
   U542 : MUXB2DL port map( A0 => n66, A1 => n1403, SL => n721, Z => n1024);
   U544 : MUXB2DL port map( A0 => n66, A1 => n1403, SL => n722, Z => n1025);
   U546 : MUXB2DL port map( A0 => n66, A1 => n1403, SL => n723, Z => n1026);
   U549 : MUXB2DL port map( A0 => n58, A1 => n1401, SL => n724, Z => n1027);
   U551 : MUXB2DL port map( A0 => n58, A1 => n1401, SL => n725, Z => n1028);
   U553 : MUXB2DL port map( A0 => n58, A1 => n1401, SL => n726, Z => n1029);
   U555 : MUXB2DL port map( A0 => n58, A1 => n1401, SL => n727, Z => n1030);
   U557 : MUXB2DL port map( A0 => n58, A1 => n1401, SL => n728, Z => n1031);
   U559 : MUXB2DL port map( A0 => n58, A1 => n1401, SL => n729, Z => n1032);
   U561 : MUXB2DL port map( A0 => n58, A1 => n1401, SL => n730, Z => n1033);
   U563 : MUXB2DL port map( A0 => n58, A1 => n1401, SL => n731, Z => n1034);
   U565 : MUXB2DL port map( A0 => n58, A1 => n1401, SL => n732, Z => n1035);
   U567 : MUXB2DL port map( A0 => n58, A1 => n1401, SL => n733, Z => n1036);
   U569 : MUXB2DL port map( A0 => n58, A1 => n1401, SL => n734, Z => n1037);
   U571 : MUXB2DL port map( A0 => n58, A1 => n1401, SL => n735, Z => n1038);
   U573 : MUXB2DL port map( A0 => n58, A1 => n1401, SL => n736, Z => n1039);
   U575 : MUXB2DL port map( A0 => n58, A1 => n1401, SL => n737, Z => n1040);
   U577 : MUXB2DL port map( A0 => n58, A1 => n1401, SL => n738, Z => n1041);
   U579 : MUXB2DL port map( A0 => n58, A1 => n1401, SL => n739, Z => n1042);
   U581 : MUXB2DL port map( A0 => n58, A1 => n1401, SL => n740, Z => n1043);
   U583 : MUXB2DL port map( A0 => n58, A1 => n1401, SL => n741, Z => n1044);
   U586 : MUXB2DL port map( A0 => n50, A1 => n1399, SL => n742, Z => n1045);
   U588 : MUXB2DL port map( A0 => n50, A1 => n1399, SL => n743, Z => n1046);
   U590 : MUXB2DL port map( A0 => n50, A1 => n1399, SL => n744, Z => n1047);
   U592 : MUXB2DL port map( A0 => n50, A1 => n1399, SL => n745, Z => n1048);
   U594 : MUXB2DL port map( A0 => n50, A1 => n1399, SL => n746, Z => n1049);
   U596 : MUXB2DL port map( A0 => n50, A1 => n1399, SL => n747, Z => n1050);
   U598 : MUXB2DL port map( A0 => n50, A1 => n1399, SL => n748, Z => n1051);
   U600 : MUXB2DL port map( A0 => n50, A1 => n1399, SL => n749, Z => n1052);
   U602 : MUXB2DL port map( A0 => n50, A1 => n1399, SL => n750, Z => n1053);
   U604 : MUXB2DL port map( A0 => n50, A1 => n1399, SL => n751, Z => n1054);
   U606 : MUXB2DL port map( A0 => n50, A1 => n1399, SL => n752, Z => n1055);
   U608 : MUXB2DL port map( A0 => n50, A1 => n1399, SL => n753, Z => n1056);
   U610 : MUXB2DL port map( A0 => n50, A1 => n1399, SL => n754, Z => n1057);
   U612 : MUXB2DL port map( A0 => n50, A1 => n1399, SL => n755, Z => n1058);
   U614 : MUXB2DL port map( A0 => n50, A1 => n1399, SL => n756, Z => n1059);
   U616 : MUXB2DL port map( A0 => n50, A1 => n1399, SL => n757, Z => n1060);
   U618 : MUXB2DL port map( A0 => n50, A1 => n1399, SL => n758, Z => n1061);
   U620 : MUXB2DL port map( A0 => n50, A1 => n1399, SL => n759, Z => n1062);
   U622 : MUXB2DL port map( A0 => n50, A1 => n1399, SL => n760, Z => n1063);
   U624 : MUXB2DL port map( A0 => n50, A1 => n1399, SL => n761, Z => n1064);
   U627 : MUXB2DL port map( A0 => n42, A1 => n1397, SL => n762, Z => n1065);
   U629 : MUXB2DL port map( A0 => n42, A1 => n1397, SL => n763, Z => n1066);
   U631 : MUXB2DL port map( A0 => n42, A1 => n1397, SL => n764, Z => n1067);
   U633 : MUXB2DL port map( A0 => n42, A1 => n1397, SL => n765, Z => n1068);
   U635 : MUXB2DL port map( A0 => n42, A1 => n1397, SL => n766, Z => n1069);
   U637 : MUXB2DL port map( A0 => n42, A1 => n1397, SL => n767, Z => n1070);
   U639 : MUXB2DL port map( A0 => n42, A1 => n1397, SL => n768, Z => n1071);
   U641 : MUXB2DL port map( A0 => n42, A1 => n1397, SL => n769, Z => n1072);
   U643 : MUXB2DL port map( A0 => n42, A1 => n1397, SL => n770, Z => n1073);
   U645 : MUXB2DL port map( A0 => n42, A1 => n1397, SL => n771, Z => n1074);
   U647 : MUXB2DL port map( A0 => n42, A1 => n1397, SL => n772, Z => n1075);
   U649 : MUXB2DL port map( A0 => n42, A1 => n1397, SL => n773, Z => n1076);
   U651 : MUXB2DL port map( A0 => n42, A1 => n1397, SL => n774, Z => n1077);
   U653 : MUXB2DL port map( A0 => n42, A1 => n1397, SL => n775, Z => n1078);
   U655 : MUXB2DL port map( A0 => n42, A1 => n1397, SL => n776, Z => n1079);
   U657 : MUXB2DL port map( A0 => n42, A1 => n1397, SL => n777, Z => n1080);
   U659 : MUXB2DL port map( A0 => n42, A1 => n1397, SL => n778, Z => n1081);
   U661 : MUXB2DL port map( A0 => n42, A1 => n1397, SL => n779, Z => n1082);
   U663 : MUXB2DL port map( A0 => n42, A1 => n1397, SL => n780, Z => n1083);
   U665 : MUXB2DL port map( A0 => n42, A1 => n1397, SL => n781, Z => n1084);
   U667 : MUXB2DL port map( A0 => n42, A1 => n1397, SL => n782, Z => n1085);
   U669 : MUXB2DL port map( A0 => n42, A1 => n1397, SL => n783, Z => n1086);
   U672 : MUXB2DL port map( A0 => n1382, A1 => n1395, SL => n784, Z => n1087);
   U674 : MUXB2DL port map( A0 => n1382, A1 => n1395, SL => n785, Z => n1088);
   U676 : MUXB2DL port map( A0 => n1382, A1 => n1395, SL => n786, Z => n1089);
   U678 : MUXB2DL port map( A0 => n1382, A1 => n1395, SL => n787, Z => n1090);
   U680 : MUXB2DL port map( A0 => n1382, A1 => n1395, SL => n788, Z => n1091);
   U682 : MUXB2DL port map( A0 => n1382, A1 => n1395, SL => n789, Z => n1092);
   U684 : MUXB2DL port map( A0 => n1382, A1 => n1395, SL => n790, Z => n1093);
   U686 : MUXB2DL port map( A0 => n1382, A1 => n1395, SL => n791, Z => n1094);
   U688 : MUXB2DL port map( A0 => n1382, A1 => n1395, SL => n792, Z => n1095);
   U690 : MUXB2DL port map( A0 => n1382, A1 => n1395, SL => n793, Z => n1096);
   U692 : MUXB2DL port map( A0 => n1382, A1 => n1395, SL => n794, Z => n1097);
   U694 : MUXB2DL port map( A0 => n1382, A1 => n1395, SL => n795, Z => n1098);
   U696 : MUXB2DL port map( A0 => n1382, A1 => n1395, SL => n796, Z => n1099);
   U698 : MUXB2DL port map( A0 => n1382, A1 => n1395, SL => n797, Z => n1100);
   U700 : MUXB2DL port map( A0 => n1382, A1 => n1395, SL => n798, Z => n1101);
   U702 : MUXB2DL port map( A0 => n1382, A1 => n1395, SL => n799, Z => n1102);
   U704 : MUXB2DL port map( A0 => n1382, A1 => n1395, SL => n800, Z => n1103);
   U706 : MUXB2DL port map( A0 => n1382, A1 => n1395, SL => n801, Z => n1104);
   U708 : MUXB2DL port map( A0 => n1382, A1 => n1395, SL => n802, Z => n1105);
   U710 : MUXB2DL port map( A0 => n1382, A1 => n1395, SL => n803, Z => n1106);
   U712 : MUXB2DL port map( A0 => n1382, A1 => n1395, SL => n804, Z => n1107);
   U714 : MUXB2DL port map( A0 => n1382, A1 => n1395, SL => n805, Z => n1108);
   U716 : MUXB2DL port map( A0 => n1382, A1 => n1395, SL => n806, Z => n1109);
   U718 : MUXB2DL port map( A0 => n1382, A1 => n1395, SL => n807, Z => n1110);
   U721 : MUXB2DL port map( A0 => n1381, A1 => n1393, SL => n808, Z => n1111);
   U723 : MUXB2DL port map( A0 => n1381, A1 => n1393, SL => n809, Z => n1112);
   U725 : MUXB2DL port map( A0 => n1381, A1 => n1393, SL => n810, Z => n1113);
   U727 : MUXB2DL port map( A0 => n1381, A1 => n1393, SL => n811, Z => n1114);
   U729 : MUXB2DL port map( A0 => n1381, A1 => n1393, SL => n812, Z => n1115);
   U731 : MUXB2DL port map( A0 => n1381, A1 => n1393, SL => n813, Z => n1116);
   U733 : MUXB2DL port map( A0 => n1381, A1 => n1393, SL => n814, Z => n1117);
   U735 : MUXB2DL port map( A0 => n1381, A1 => n1393, SL => n815, Z => n1118);
   U737 : MUXB2DL port map( A0 => n1381, A1 => n1393, SL => n816, Z => n1119);
   U739 : MUXB2DL port map( A0 => n1381, A1 => n1393, SL => n817, Z => n1120);
   U741 : MUXB2DL port map( A0 => n1381, A1 => n1393, SL => n818, Z => n1121);
   U743 : MUXB2DL port map( A0 => n1381, A1 => n1393, SL => n819, Z => n1122);
   U745 : MUXB2DL port map( A0 => n1381, A1 => n1393, SL => n820, Z => n1123);
   U747 : MUXB2DL port map( A0 => n1381, A1 => n1393, SL => n821, Z => n1124);
   U749 : MUXB2DL port map( A0 => n1381, A1 => n1393, SL => n822, Z => n1125);
   U751 : MUXB2DL port map( A0 => n1381, A1 => n1393, SL => n823, Z => n1126);
   U753 : MUXB2DL port map( A0 => n1381, A1 => n1393, SL => n824, Z => n1127);
   U755 : MUXB2DL port map( A0 => n1381, A1 => n1393, SL => n825, Z => n1128);
   U757 : MUXB2DL port map( A0 => n1381, A1 => n1393, SL => n826, Z => n1129);
   U759 : MUXB2DL port map( A0 => n1381, A1 => n1393, SL => n827, Z => n1130);
   U761 : MUXB2DL port map( A0 => n1381, A1 => n1393, SL => n828, Z => n1131);
   U763 : MUXB2DL port map( A0 => n1381, A1 => n1393, SL => n829, Z => n1132);
   U765 : MUXB2DL port map( A0 => n1381, A1 => n1393, SL => n830, Z => n1133);
   U767 : MUXB2DL port map( A0 => n1381, A1 => n1393, SL => n831, Z => n1134);
   U769 : MUXB2DL port map( A0 => n1381, A1 => n1393, SL => n832, Z => n1135);
   U771 : MUXB2DL port map( A0 => n1381, A1 => n1393, SL => n833, Z => n1136);
   U774 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n834, Z => n1137);
   U776 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n835, Z => n1138);
   U778 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n836, Z => n1139);
   U780 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n837, Z => n1140);
   U782 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n838, Z => n1141);
   U784 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n839, Z => n1142);
   U786 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n840, Z => n1143);
   U788 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n841, Z => n1144);
   U790 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n842, Z => n1145);
   U792 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n843, Z => n1146);
   U794 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n844, Z => n1147);
   U796 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n845, Z => n1148);
   U798 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n846, Z => n1149);
   U800 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n847, Z => n1150);
   U802 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n848, Z => n1151);
   U804 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n849, Z => n1152);
   U806 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n850, Z => n1153);
   U808 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n851, Z => n1154);
   U810 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n852, Z => n1155);
   U812 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n853, Z => n1156);
   U814 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n854, Z => n1157);
   U816 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n855, Z => n1158);
   U818 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n856, Z => n1159);
   U820 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n857, Z => n1160);
   U822 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n858, Z => n1161);
   U824 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n859, Z => n1162);
   U826 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n860, Z => n1163);
   U828 : MUXB2DL port map( A0 => n1380, A1 => n1391, SL => n861, Z => n1164);
   U831 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n862, Z => n1165);
   U833 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n863, Z => n1166);
   U835 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n864, Z => n1167);
   U837 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n865, Z => n1168);
   U839 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n866, Z => n1169);
   U841 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n867, Z => n1170);
   U843 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n868, Z => n1171);
   U845 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n869, Z => n1172);
   U847 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n870, Z => n1173);
   U849 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n871, Z => n1174);
   U851 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n872, Z => n1175);
   U853 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n873, Z => n1176);
   U855 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n874, Z => n1177);
   U857 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n875, Z => n1178);
   U859 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n876, Z => n1179);
   U861 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n877, Z => n1180);
   U863 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n878, Z => n1181);
   U865 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n879, Z => n1182);
   U867 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n880, Z => n1183);
   U869 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n881, Z => n1184);
   U871 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n882, Z => n1185);
   U873 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n883, Z => n1186);
   U875 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n884, Z => n1187);
   U877 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n885, Z => n1188);
   U879 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n886, Z => n1189);
   U881 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n887, Z => n1190);
   U883 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n888, Z => n1191);
   U885 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n889, Z => n1192);
   U887 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n890, Z => n1193);
   U889 : MUXB2DL port map( A0 => n1379, A1 => n1390, SL => n891, Z => n1194);
   U892 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n892, Z => n1195);
   U894 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n893, Z => n1196);
   U896 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n894, Z => n1197);
   U898 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n895, Z => n1198);
   U900 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n896, Z => n1199);
   U902 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n897, Z => n1200);
   U904 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n898, Z => n1201);
   U906 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n899, Z => n1202);
   U908 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n900, Z => n1203);
   U910 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n901, Z => n1204);
   U912 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n902, Z => n1205);
   U914 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n903, Z => n1206);
   U916 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n904, Z => n1207);
   U918 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n905, Z => n1208);
   U920 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n906, Z => n1209);
   U922 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n907, Z => n1210);
   U924 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n908, Z => n1211);
   U926 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n909, Z => n1212);
   U928 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n910, Z => n1213);
   U930 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n911, Z => n1214);
   U932 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n912, Z => n1215);
   U934 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n913, Z => n1216);
   U936 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n914, Z => n1217);
   U938 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n915, Z => n1218);
   U940 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n916, Z => n1219);
   U942 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n917, Z => n1220);
   U944 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n918, Z => n1221);
   U946 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n919, Z => n1222);
   U948 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n920, Z => n1223);
   U950 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n921, Z => n1224);
   U952 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n922, Z => n1225);
   U954 : MUXB2DL port map( A0 => n1378, A1 => n1389, SL => n923, Z => n1226);
   U1021 : EXOR2D1 port map( A1 => a(4), A2 => a(3), Z => n1375);
   U1022 : EXOR2D1 port map( A1 => a(6), A2 => a(5), Z => n1376);
   U1023 : EXOR2D1 port map( A1 => a(8), A2 => a(7), Z => n1377);
   U1024 : NAN2D1 port map( A1 => a(0), A2 => n1389, Z => n1378);
   U1025 : OAI21D1 port map( A1 => a(2), A2 => a(1), B => n1392, Z => n1379);
   U1026 : OAI21D1 port map( A1 => a(4), A2 => a(3), B => n1394, Z => n1380);
   U1027 : OAI21D1 port map( A1 => a(6), A2 => a(5), B => n1396, Z => n1381);
   U1028 : OAI21D1 port map( A1 => a(8), A2 => a(7), B => n1398, Z => n1382);
   U1029 : INVD1 port map( A => n1383, Z => n1384);
   U1030 : INVD1 port map( A => n953, Z => n1390);
   U1031 : INVD1 port map( A => n952, Z => n1391);
   U1032 : INVD1 port map( A => n951, Z => n1393);
   U1033 : INVD1 port map( A => n950, Z => n1395);
   U1034 : INVD1 port map( A => n949, Z => n1397);
   U1035 : INVD1 port map( A => n948, Z => n1399);
   U1036 : INVD1 port map( A => n947, Z => n1401);
   U1037 : INVD1 port map( A => n946, Z => n1403);
   U1038 : INVD1 port map( A => n945, Z => n1405);
   U1039 : INVD1 port map( A => n944, Z => n1407);
   U1040 : INVD1 port map( A => n943, Z => n1409);
   U1041 : INVD1 port map( A => n942, Z => n1411);
   U1042 : INVD1 port map( A => n941, Z => n1413);
   U1043 : INVD1 port map( A => n940, Z => n1416);
   U1044 : INVD1 port map( A => n939, Z => n1417);
   U1045 : INVD1 port map( A => a(1), Z => n1389);
   U1046 : EXNOR2D1 port map( A1 => a(2), A2 => a(1), Z => n1383);
   U1047 : INVD1 port map( A => n1388, Z => n1387);
   U1048 : INVD1 port map( A => n1386, Z => n1385);
   U1049 : INVD1 port map( A => a(3), Z => n1392);
   U1050 : INVD1 port map( A => a(5), Z => n1394);
   U1051 : INVD1 port map( A => a(7), Z => n1396);
   U1052 : INVD1 port map( A => a(9), Z => n1398);
   U1053 : EXOR2D1 port map( A1 => a(10), A2 => a(9), Z => n1438);
   U1054 : INVD1 port map( A => a(11), Z => n1400);
   U1055 : OAI21D1 port map( A1 => a(9), A2 => a(10), B => n1400, Z => n42);
   U1056 : EXOR2D1 port map( A1 => a(12), A2 => a(11), Z => n1439);
   U1057 : INVD1 port map( A => a(13), Z => n1402);
   U1058 : OAI21D1 port map( A1 => a(12), A2 => a(11), B => n1402, Z => n50);
   U1059 : EXOR2D1 port map( A1 => a(14), A2 => a(13), Z => n1440);
   U1060 : INVD1 port map( A => a(15), Z => n1404);
   U1061 : OAI21D1 port map( A1 => a(14), A2 => a(13), B => n1404, Z => n58);
   U1062 : EXOR2D1 port map( A1 => a(16), A2 => a(15), Z => n1441);
   U1063 : INVD1 port map( A => a(17), Z => n1406);
   U1064 : OAI21D1 port map( A1 => a(16), A2 => a(15), B => n1406, Z => n66);
   U1065 : EXOR2D1 port map( A1 => a(18), A2 => a(17), Z => n1442);
   U1066 : INVD1 port map( A => a(19), Z => n1408);
   U1067 : OAI21D1 port map( A1 => a(18), A2 => a(17), B => n1408, Z => n73);
   U1068 : EXOR2D1 port map( A1 => a(20), A2 => a(19), Z => n1443);
   U1069 : INVD1 port map( A => a(21), Z => n1410);
   U1070 : OAI21D1 port map( A1 => a(20), A2 => a(19), B => n1410, Z => n80);
   U1071 : EXOR2D1 port map( A1 => a(22), A2 => a(21), Z => n1444);
   U1072 : INVD1 port map( A => a(23), Z => n1412);
   U1073 : OAI21D1 port map( A1 => a(22), A2 => a(21), B => n1412, Z => n84);
   U1074 : INVD1 port map( A => a(25), Z => n1414);
   U1075 : INVD1 port map( A => a(27), Z => n1415);
   U1076 : INVD1 port map( A => a(29), Z => n1418);
   U1077 : MUXB2DL port map( A0 => b(29), A1 => b(28), SL => n1383, Z => n862);
   U1078 : INVD1 port map( A => b(1), Z => n1388);
   U1079 : INVD1 port map( A => b(3), Z => n1386);
   U1080 : INVD1 port map( A => a(31), Z => n1419);
   U1081 : EXOR3D1 port map( A1 => n1420, A2 => n1421, A3 => n1422, Z => 
                           product(31));
   U1082 : EXOR3D1 port map( A1 => n208, A2 => n206, A3 => n1423, Z => n1422);
   U1083 : EXOR2D1 port map( A1 => n214, A2 => n212, Z => n1423);
   U1084 : EXOR2D1 port map( A1 => n202, A2 => n156, Z => n1421);
   U1085 : EXOR3D1 port map( A1 => n1424, A2 => n1425, A3 => n1426, Z => n1420)
                           ;
   U1086 : EXOR3D1 port map( A1 => n957, A2 => n955, A3 => n1427, Z => n1426);
   U1087 : EXNOR2D1 port map( A1 => n997, A2 => n975, Z => n1427);
   U1088 : EXOR3D1 port map( A1 => n1428, A2 => n204, A3 => n1429, Z => n1425);
   U1089 : EXOR3D1 port map( A1 => n1087, A2 => n1065, A3 => n1430, Z => n1429)
                           ;
   U1090 : EXNOR2D1 port map( A1 => n210, A2 => n1111, Z => n1430);
   U1091 : EXOR3D1 port map( A1 => n961, A2 => n218, A3 => n1431, Z => n1428);
   U1092 : EXOR2D1 port map( A1 => n985, A2 => n967, Z => n1431);
   U1093 : EXOR3D1 port map( A1 => n1432, A2 => n1433, A3 => n1434, Z => n1424)
                           ;
   U1094 : EXOR3D1 port map( A1 => n1027, A2 => n1011, A3 => n1435, Z => n1434)
                           ;
   U1095 : EXOR3D1 port map( A1 => n1165, A2 => n1137, A3 => n1045, Z => n1435)
                           ;
   U1096 : EXOR3D1 port map( A1 => n216, A2 => n1195, A3 => n1436, Z => n1433);
   U1097 : EXOR2D1 port map( A1 => n222, A2 => n220, Z => n1436);
   U1098 : EXOR3D1 port map( A1 => n226, A2 => n224, A3 => n1437, Z => n1432);
   U1099 : EXOR2D1 port map( A1 => n230, A2 => n228, Z => n1437);
   U1100 : OAI21D1 port map( A1 => a(28), A2 => a(27), B => n1418, Z => n99);
   U1101 : AOI21D1 port map( A1 => a(25), A2 => a(26), B => n1415, Z => n941);
   U1102 : OAI21D1 port map( A1 => a(26), A2 => a(25), B => n1415, Z => n94);
   U1103 : NAN2D1 port map( A1 => b(0), A2 => a(0), Z => n923);
   U1104 : MUXB2DL port map( A0 => b(0), A1 => n1387, SL => a(0), Z => n922);
   U1105 : MUXB2DL port map( A0 => n1387, A1 => b(2), SL => a(0), Z => n921);
   U1106 : MUXB2DL port map( A0 => b(2), A1 => n1385, SL => a(0), Z => n920);
   U1107 : MUXB2DL port map( A0 => n1385, A1 => b(4), SL => a(0), Z => n919);
   U1108 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => a(0), Z => n918);
   U1109 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => a(0), Z => n917);
   U1110 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => a(0), Z => n916);
   U1111 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => a(0), Z => n915);
   U1112 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => a(0), Z => n914);
   U1113 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => a(0), Z => n913);
   U1114 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => a(0), Z => n912);
   U1115 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => a(0), Z => n911);
   U1116 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => a(0), Z => n910);
   U1117 : AOI21D1 port map( A1 => a(23), A2 => a(24), B => n1414, Z => n942);
   U1118 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => a(0), Z => n909);
   U1119 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => a(0), Z => n908);
   U1120 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => a(0), Z => n907);
   U1121 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => a(0), Z => n906);
   U1122 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => a(0), Z => n905);
   U1123 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => a(0), Z => n904);
   U1124 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => a(0), Z => n903);
   U1125 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => a(0), Z => n902);
   U1126 : MUXB2DL port map( A0 => b(21), A1 => b(22), SL => a(0), Z => n901);
   U1127 : MUXB2DL port map( A0 => b(22), A1 => b(23), SL => a(0), Z => n900);
   U1128 : MUXB2DL port map( A0 => b(23), A1 => b(24), SL => a(0), Z => n899);
   U1129 : MUXB2DL port map( A0 => b(24), A1 => b(25), SL => a(0), Z => n898);
   U1130 : MUXB2DL port map( A0 => b(25), A1 => b(26), SL => a(0), Z => n897);
   U1131 : MUXB2DL port map( A0 => b(26), A1 => b(27), SL => a(0), Z => n896);
   U1132 : MUXB2DL port map( A0 => b(27), A1 => b(28), SL => a(0), Z => n895);
   U1133 : MUXB2DL port map( A0 => b(28), A1 => b(29), SL => a(0), Z => n894);
   U1134 : MUXB2DL port map( A0 => b(29), A1 => b(30), SL => a(0), Z => n893);
   U1135 : MUXB2DL port map( A0 => b(30), A1 => b(31), SL => a(0), Z => n892);
   U1136 : NAN2D1 port map( A1 => b(0), A2 => n1384, Z => n891);
   U1137 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1384, Z => n890);
   U1138 : OAI21D1 port map( A1 => a(24), A2 => a(23), B => n1414, Z => n89);
   U1139 : MUXB2DL port map( A0 => n1387, A1 => b(2), SL => n1384, Z => n889);
   U1140 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1384, Z => n888);
   U1141 : MUXB2DL port map( A0 => n1385, A1 => b(4), SL => n1384, Z => n887);
   U1142 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1384, Z => n886);
   U1143 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1384, Z => n885);
   U1144 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1384, Z => n884);
   U1145 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1384, Z => n883);
   U1146 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1384, Z => n882);
   U1147 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1384, Z => n881);
   U1148 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1384, Z => n880);
   U1149 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1384, Z => n879);
   U1150 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1384, Z => n878);
   U1151 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1384, Z => n877);
   U1152 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1384, Z => n876);
   U1153 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1384, Z => n875);
   U1154 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1384, Z => n874);
   U1155 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1384, Z => n873);
   U1156 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1384, Z => n872);
   U1157 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => n1384, Z => n871);
   U1158 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => n1384, Z => n870);
   U1159 : MUXB2DL port map( A0 => b(21), A1 => b(22), SL => n1384, Z => n869);
   U1160 : MUXB2DL port map( A0 => b(22), A1 => b(23), SL => n1384, Z => n868);
   U1161 : MUXB2DL port map( A0 => b(23), A1 => b(24), SL => n1384, Z => n867);
   U1162 : MUXB2DL port map( A0 => b(24), A1 => b(25), SL => n1384, Z => n866);
   U1163 : MUXB2DL port map( A0 => b(25), A1 => b(26), SL => n1384, Z => n865);
   U1164 : MUXB2DL port map( A0 => b(26), A1 => b(27), SL => n1384, Z => n864);
   U1165 : MUXB2DL port map( A0 => b(27), A1 => b(28), SL => n1384, Z => n863);
   U1166 : NAN2D1 port map( A1 => b(0), A2 => n1375, Z => n861);
   U1167 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1375, Z => n860);
   U1168 : AOI21D1 port map( A1 => a(21), A2 => a(22), B => n1412, Z => n943);
   U1169 : MUXB2DL port map( A0 => n1387, A1 => b(2), SL => n1375, Z => n859);
   U1170 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1375, Z => n858);
   U1171 : MUXB2DL port map( A0 => n1385, A1 => b(4), SL => n1375, Z => n857);
   U1172 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1375, Z => n856);
   U1173 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1375, Z => n855);
   U1174 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1375, Z => n854);
   U1175 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1375, Z => n853);
   U1176 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1375, Z => n852);
   U1177 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1375, Z => n851);
   U1178 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1375, Z => n850);
   U1179 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1375, Z => n849);
   U1180 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1375, Z => n848);
   U1181 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1375, Z => n847);
   U1182 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1375, Z => n846);
   U1183 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1375, Z => n845);
   U1184 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1375, Z => n844);
   U1185 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1375, Z => n843);
   U1186 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1375, Z => n842);
   U1187 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => n1375, Z => n841);
   U1188 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => n1375, Z => n840);
   U1189 : MUXB2DL port map( A0 => b(21), A1 => b(22), SL => n1375, Z => n839);
   U1190 : MUXB2DL port map( A0 => b(22), A1 => b(23), SL => n1375, Z => n838);
   U1191 : MUXB2DL port map( A0 => b(23), A1 => b(24), SL => n1375, Z => n837);
   U1192 : MUXB2DL port map( A0 => b(24), A1 => b(25), SL => n1375, Z => n836);
   U1193 : MUXB2DL port map( A0 => b(25), A1 => b(26), SL => n1375, Z => n835);
   U1194 : MUXB2DL port map( A0 => b(26), A1 => b(27), SL => n1375, Z => n834);
   U1195 : NAN2D1 port map( A1 => b(0), A2 => n1376, Z => n833);
   U1196 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1376, Z => n832);
   U1197 : MUXB2DL port map( A0 => n1387, A1 => b(2), SL => n1376, Z => n831);
   U1198 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1376, Z => n830);
   U1199 : MUXB2DL port map( A0 => n1385, A1 => b(4), SL => n1376, Z => n829);
   U1200 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1376, Z => n828);
   U1201 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1376, Z => n827);
   U1202 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1376, Z => n826);
   U1203 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1376, Z => n825);
   U1204 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1376, Z => n824);
   U1205 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1376, Z => n823);
   U1206 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1376, Z => n822);
   U1207 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1376, Z => n821);
   U1208 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1376, Z => n820);
   U1209 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1376, Z => n819);
   U1210 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1376, Z => n818);
   U1211 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1376, Z => n817);
   U1212 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1376, Z => n816);
   U1213 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1376, Z => n815);
   U1214 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1376, Z => n814);
   U1215 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => n1376, Z => n813);
   U1216 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => n1376, Z => n812);
   U1217 : MUXB2DL port map( A0 => b(21), A1 => b(22), SL => n1376, Z => n811);
   U1218 : MUXB2DL port map( A0 => b(22), A1 => b(23), SL => n1376, Z => n810);
   U1219 : AOI21D1 port map( A1 => a(19), A2 => a(20), B => n1410, Z => n944);
   U1220 : MUXB2DL port map( A0 => b(23), A1 => b(24), SL => n1376, Z => n809);
   U1221 : MUXB2DL port map( A0 => b(24), A1 => b(25), SL => n1376, Z => n808);
   U1222 : NAN2D1 port map( A1 => b(0), A2 => n1377, Z => n807);
   U1223 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1377, Z => n806);
   U1224 : MUXB2DL port map( A0 => b(1), A1 => b(2), SL => n1377, Z => n805);
   U1225 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1377, Z => n804);
   U1226 : MUXB2DL port map( A0 => n1385, A1 => b(4), SL => n1377, Z => n803);
   U1227 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1377, Z => n802);
   U1228 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1377, Z => n801);
   U1229 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1377, Z => n800);
   U1230 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1377, Z => n799);
   U1231 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1377, Z => n798);
   U1232 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1377, Z => n797);
   U1233 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1377, Z => n796);
   U1234 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1377, Z => n795);
   U1235 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1377, Z => n794);
   U1236 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1377, Z => n793);
   U1237 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1377, Z => n792);
   U1238 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1377, Z => n791);
   U1239 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1377, Z => n790);
   U1240 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1377, Z => n789);
   U1241 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1377, Z => n788);
   U1242 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => n1377, Z => n787);
   U1243 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => n1377, Z => n786);
   U1244 : MUXB2DL port map( A0 => b(21), A1 => b(22), SL => n1377, Z => n785);
   U1245 : MUXB2DL port map( A0 => b(22), A1 => b(23), SL => n1377, Z => n784);
   U1246 : NAN2D1 port map( A1 => b(0), A2 => n1438, Z => n783);
   U1247 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1438, Z => n782);
   U1248 : MUXB2DL port map( A0 => n1387, A1 => b(2), SL => n1438, Z => n781);
   U1249 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1438, Z => n780);
   U1250 : MUXB2DL port map( A0 => b(3), A1 => b(4), SL => n1438, Z => n779);
   U1251 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1438, Z => n778);
   U1252 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1438, Z => n777);
   U1253 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1438, Z => n776);
   U1254 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1438, Z => n775);
   U1255 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1438, Z => n774);
   U1256 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1438, Z => n773);
   U1257 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1438, Z => n772);
   U1258 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1438, Z => n771);
   U1259 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1438, Z => n770);
   U1260 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1438, Z => n769);
   U1261 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1438, Z => n768);
   U1262 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1438, Z => n767);
   U1263 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1438, Z => n766);
   U1264 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1438, Z => n765);
   U1265 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1438, Z => n764);
   U1266 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => n1438, Z => n763);
   U1267 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => n1438, Z => n762);
   U1268 : NAN2D1 port map( A1 => b(0), A2 => n1439, Z => n761);
   U1269 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1439, Z => n760);
   U1270 : MUXB2DL port map( A0 => b(1), A1 => b(2), SL => n1439, Z => n759);
   U1271 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1439, Z => n758);
   U1272 : MUXB2DL port map( A0 => n1385, A1 => b(4), SL => n1439, Z => n757);
   U1273 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1439, Z => n756);
   U1274 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1439, Z => n755);
   U1275 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1439, Z => n754);
   U1276 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1439, Z => n753);
   U1277 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1439, Z => n752);
   U1278 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1439, Z => n751);
   U1279 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1439, Z => n750);
   U1280 : AOI21D1 port map( A1 => a(17), A2 => a(18), B => n1408, Z => n945);
   U1281 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1439, Z => n749);
   U1282 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1439, Z => n748);
   U1283 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1439, Z => n747);
   U1284 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1439, Z => n746);
   U1285 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1439, Z => n745);
   U1286 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1439, Z => n744);
   U1287 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1439, Z => n743);
   U1288 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1439, Z => n742);
   U1289 : NAN2D1 port map( A1 => b(0), A2 => n1440, Z => n741);
   U1290 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1440, Z => n740);
   U1291 : MUXB2DL port map( A0 => n1387, A1 => b(2), SL => n1440, Z => n739);
   U1292 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1440, Z => n738);
   U1293 : MUXB2DL port map( A0 => n1385, A1 => b(4), SL => n1440, Z => n737);
   U1294 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1440, Z => n736);
   U1295 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1440, Z => n735);
   U1296 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1440, Z => n734);
   U1297 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1440, Z => n733);
   U1298 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1440, Z => n732);
   U1299 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1440, Z => n731);
   U1300 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1440, Z => n730);
   U1301 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1440, Z => n729);
   U1302 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1440, Z => n728);
   U1303 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1440, Z => n727);
   U1304 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1440, Z => n726);
   U1305 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1440, Z => n725);
   U1306 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1440, Z => n724);
   U1307 : NAN2D1 port map( A1 => b(0), A2 => n1441, Z => n723);
   U1308 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1441, Z => n722);
   U1309 : MUXB2DL port map( A0 => n1387, A1 => b(2), SL => n1441, Z => n721);
   U1310 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1441, Z => n720);
   U1311 : MUXB2DL port map( A0 => n1385, A1 => b(4), SL => n1441, Z => n719);
   U1312 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1441, Z => n718);
   U1313 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1441, Z => n717);
   U1314 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1441, Z => n716);
   U1315 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1441, Z => n715);
   U1316 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1441, Z => n714);
   U1317 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1441, Z => n713);
   U1318 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1441, Z => n712);
   U1319 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1441, Z => n711);
   U1320 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1441, Z => n710);
   U1321 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1441, Z => n709);
   U1322 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1441, Z => n708);
   U1323 : NAN2D1 port map( A1 => b(0), A2 => n1442, Z => n707);
   U1324 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1442, Z => n706);
   U1325 : MUXB2DL port map( A0 => n1387, A1 => b(2), SL => n1442, Z => n705);
   U1326 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1442, Z => n704);
   U1327 : MUXB2DL port map( A0 => n1385, A1 => b(4), SL => n1442, Z => n703);
   U1328 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1442, Z => n702);
   U1329 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1442, Z => n701);
   U1330 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1442, Z => n700);
   U1331 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1442, Z => n699);
   U1332 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1442, Z => n698);
   U1333 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1442, Z => n697);
   U1334 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1442, Z => n696);
   U1335 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1442, Z => n695);
   U1336 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1442, Z => n694);
   U1337 : NAN2D1 port map( A1 => b(0), A2 => n1443, Z => n693);
   U1338 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1443, Z => n692);
   U1339 : MUXB2DL port map( A0 => n1387, A1 => b(2), SL => n1443, Z => n691);
   U1340 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1443, Z => n690);
   U1341 : MUXB2DL port map( A0 => n1385, A1 => b(4), SL => n1443, Z => n689);
   U1342 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1443, Z => n688);
   U1343 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1443, Z => n687);
   U1344 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1443, Z => n686);
   U1345 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1443, Z => n685);
   U1346 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1443, Z => n684);
   U1347 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1443, Z => n683);
   U1348 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1443, Z => n682);
   U1349 : NAN2D1 port map( A1 => b(0), A2 => n1444, Z => n681);
   U1350 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1444, Z => n680);
   U1351 : AOI21D1 port map( A1 => a(15), A2 => a(16), B => n1406, Z => n946);
   U1352 : MUXB2DL port map( A0 => n1387, A1 => b(2), SL => n1444, Z => n679);
   U1353 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1444, Z => n678);
   U1354 : MUXB2DL port map( A0 => n1385, A1 => b(4), SL => n1444, Z => n677);
   U1355 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1444, Z => n676);
   U1356 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1444, Z => n675);
   U1357 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1444, Z => n674);
   U1358 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1444, Z => n673);
   U1359 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1444, Z => n672);
   U1360 : NAN2D1 port map( A1 => b(0), A2 => n1445, Z => n671);
   U1361 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1445, Z => n670);
   U1362 : MUXB2DL port map( A0 => n1387, A1 => b(2), SL => n1445, Z => n669);
   U1363 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1445, Z => n668);
   U1364 : MUXB2DL port map( A0 => n1385, A1 => b(4), SL => n1445, Z => n667);
   U1365 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1445, Z => n666);
   U1366 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1445, Z => n665);
   U1367 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1445, Z => n664);
   U1368 : EXOR2D1 port map( A1 => a(24), A2 => a(23), Z => n1445);
   U1369 : NAN2D1 port map( A1 => b(0), A2 => n1446, Z => n663);
   U1370 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1446, Z => n662);
   U1371 : MUXB2DL port map( A0 => n1387, A1 => b(2), SL => n1446, Z => n661);
   U1372 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1446, Z => n660);
   U1373 : MUXB2DL port map( A0 => n1385, A1 => b(4), SL => n1446, Z => n659);
   U1374 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1446, Z => n658);
   U1375 : EXOR2D1 port map( A1 => a(26), A2 => a(25), Z => n1446);
   U1376 : NAN2D1 port map( A1 => b(0), A2 => n1447, Z => n657);
   U1377 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1447, Z => n656);
   U1378 : MUXB2DL port map( A0 => n1387, A1 => b(2), SL => n1447, Z => n655);
   U1379 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1447, Z => n654);
   U1380 : EXOR2D1 port map( A1 => a(28), A2 => a(27), Z => n1447);
   U1381 : NAN2D1 port map( A1 => b(0), A2 => n1448, Z => n653);
   U1382 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1448, Z => n652);
   U1383 : EXOR2D1 port map( A1 => a(30), A2 => a(29), Z => n1448);
   U1384 : AOI21D1 port map( A1 => a(13), A2 => a(14), B => n1404, Z => n947);
   U1385 : AOI21D1 port map( A1 => a(11), A2 => a(12), B => n1402, Z => n948);
   U1386 : AOI21D1 port map( A1 => a(9), A2 => a(10), B => n1400, Z => n949);
   U1387 : AOI21D1 port map( A1 => a(7), A2 => a(8), B => n1398, Z => n950);
   U1388 : AOI21D1 port map( A1 => a(5), A2 => a(6), B => n1396, Z => n951);
   U1389 : AOI21D1 port map( A1 => a(3), A2 => a(4), B => n1394, Z => n952);
   U1390 : AOI21D1 port map( A1 => a(1), A2 => a(2), B => n1392, Z => n953);
   U1391 : AOI21D1 port map( A1 => a(29), A2 => a(30), B => n1419, Z => n939);
   U1392 : OAI21D1 port map( A1 => a(30), A2 => a(29), B => n1419, Z => n104);
   U1393 : AOI21D1 port map( A1 => a(27), A2 => a(28), B => n1418, Z => n940);

end hier_filter_none_20;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_gp_custom.all;

architecture hier_filter_none_20 of gp_custom_DW_mult_tc_3 is

   component AOI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component MUXB2DL
      port( A0, A1, SL : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal n42, n50, n58, n66, n73, n80, n84, n89, n94, n99, n104, n156, n157, 
      n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, 
      n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, 
      n182, n183, n184, n185, n186, n202, n203, n204, n205, n206, n207, n208, 
      n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, 
      n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, 
      n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, 
      n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, 
      n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, 
      n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, 
      n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
      n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, 
      n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, 
      n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, 
      n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, 
      n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, 
      n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, 
      n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, 
      n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, 
      n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, 
      n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, 
      n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, 
      n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, 
      n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, 
      n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, 
      n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, 
      n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, 
      n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, 
      n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, 
      n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, 
      n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
      n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, 
      n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, 
      n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, 
      n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
      n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, 
      n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, 
      n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, 
      n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, 
      n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, 
      n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, 
      n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, 
      n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, 
      n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, 
      n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, 
      n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, 
      n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, 
      n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, 
      n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, 
      n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, 
      n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, 
      n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, 
      n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, 
      n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, 
      n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, 
      n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, 
      n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, 
      n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, 
      n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, 
      n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, 
      n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, 
      n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, 
      n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, 
      n917, n918, n919, n920, n921, n922, n923, n939, n940, n941, n942, n943, 
      n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n955, n956, 
      n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, 
      n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, 
      n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, 
      n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, 
      n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, 
      n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, 
      n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, 
      n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, 
      n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, 
      n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, 
      n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, 
      n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, 
      n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, 
      n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, 
      n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, 
      n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, 
      n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, 
      n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, 
      n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, 
      n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, 
      n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, 
      n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, 
      n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, 
      n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, 
      n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, 
      n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, 
      n1224, n1225, n1226, n1375, n1376, n1377, n1378, n1379, n1380, n1381, 
      n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, 
      n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, 
      n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, 
      n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, 
      n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, 
      n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, 
      n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451 : 
      std_logic;

begin
   
   U125 : ADFULD1 port map( A => n203, B => n232, CI => n157, CO => n156, S => 
                           product(30));
   U126 : ADFULD1 port map( A => n233, B => n260, CI => n158, CO => n157, S => 
                           product(29));
   U127 : ADFULD1 port map( A => n261, B => n288, CI => n159, CO => n158, S => 
                           product(28));
   U128 : ADFULD1 port map( A => n289, B => n314, CI => n160, CO => n159, S => 
                           product(27));
   U129 : ADFULD1 port map( A => n315, B => n340, CI => n161, CO => n160, S => 
                           product(26));
   U130 : ADFULD1 port map( A => n341, B => n364, CI => n162, CO => n161, S => 
                           product(25));
   U131 : ADFULD1 port map( A => n365, B => n388, CI => n163, CO => n162, S => 
                           product(24));
   U132 : ADFULD1 port map( A => n389, B => n410, CI => n164, CO => n163, S => 
                           product(23));
   U133 : ADFULD1 port map( A => n411, B => n432, CI => n165, CO => n164, S => 
                           product(22));
   U134 : ADFULD1 port map( A => n433, B => n452, CI => n166, CO => n165, S => 
                           product(21));
   U135 : ADFULD1 port map( A => n453, B => n472, CI => n167, CO => n166, S => 
                           product(20));
   U136 : ADFULD1 port map( A => n473, B => n490, CI => n168, CO => n167, S => 
                           product(19));
   U137 : ADFULD1 port map( A => n491, B => n508, CI => n169, CO => n168, S => 
                           product(18));
   U138 : ADFULD1 port map( A => n509, B => n524, CI => n170, CO => n169, S => 
                           product(17));
   U139 : ADFULD1 port map( A => n525, B => n540, CI => n171, CO => n170, S => 
                           product(16));
   U140 : ADFULD1 port map( A => n541, B => n554, CI => n172, CO => n171, S => 
                           product(15));
   U141 : ADFULD1 port map( A => n555, B => n568, CI => n173, CO => n172, S => 
                           product(14));
   U142 : ADFULD1 port map( A => n569, B => n580, CI => n174, CO => n173, S => 
                           product(13));
   U143 : ADFULD1 port map( A => n581, B => n592, CI => n175, CO => n174, S => 
                           product(12));
   U144 : ADFULD1 port map( A => n593, B => n602, CI => n176, CO => n175, S => 
                           product(11));
   U145 : ADFULD1 port map( A => n603, B => n612, CI => n177, CO => n176, S => 
                           product(10));
   U146 : ADFULD1 port map( A => n613, B => n620, CI => n178, CO => n177, S => 
                           product(9));
   U147 : ADFULD1 port map( A => n621, B => n628, CI => n179, CO => n178, S => 
                           product(8));
   U148 : ADFULD1 port map( A => n629, B => n634, CI => n180, CO => n179, S => 
                           product(7));
   U149 : ADFULD1 port map( A => n635, B => n640, CI => n181, CO => n180, S => 
                           product(6));
   U150 : ADFULD1 port map( A => n641, B => n644, CI => n182, CO => n181, S => 
                           product(5));
   U151 : ADFULD1 port map( A => n645, B => n648, CI => n183, CO => n182, S => 
                           product(4));
   U152 : ADFULD1 port map( A => n649, B => n1193, CI => n184, CO => n183, S =>
                           product(3));
   U153 : ADFULD1 port map( A => n651, B => n1194, CI => n185, CO => n184, S =>
                           product(2));
   U154 : ADHALFDL port map( A => n186, B => n1225, CO => n185, S => product(1)
                           );
   U155 : ADHALFDL port map( A => n1226, B => a(1), CO => n186, S => product(0)
                           );
   U171 : ADFULD1 port map( A => n234, B => n207, CI => n205, CO => n202, S => 
                           n203);
   U172 : ADFULD1 port map( A => n209, B => n211, CI => n236, CO => n204, S => 
                           n205);
   U173 : ADFULD1 port map( A => n240, B => n213, CI => n238, CO => n206, S => 
                           n207);
   U174 : ADFULD1 port map( A => n217, B => n242, CI => n215, CO => n208, S => 
                           n209);
   U175 : ADFULD1 port map( A => n244, B => n246, CI => n219, CO => n210, S => 
                           n211);
   U176 : ADFULD1 port map( A => n225, B => n223, CI => n248, CO => n212, S => 
                           n213);
   U177 : ADFULD1 port map( A => n221, B => n229, CI => n227, CO => n214, S => 
                           n215);
   U178 : ADFULD1 port map( A => n256, B => n252, CI => n254, CO => n216, S => 
                           n217);
   U179 : ADFULD1 port map( A => n258, B => n1088, CI => n250, CO => n218, S =>
                           n219);
   U180 : ADFULD1 port map( A => n1046, B => n1112, CI => n1066, CO => n220, S 
                           => n221);
   U181 : ADFULD1 port map( A => n986, B => n976, CI => n998, CO => n222, S => 
                           n223);
   U182 : ADFULD1 port map( A => n962, B => n1138, CI => n968, CO => n224, S =>
                           n225);
   U183 : ADFULD1 port map( A => n1166, B => n1012, CI => n231, CO => n226, S 
                           => n227);
   U184 : ADFULD1 port map( A => n1028, B => n956, CI => n958, CO => n228, S =>
                           n229);
   U185 : ADHALFDL port map( A => n1196, B => n939, CO => n230, S => n231);
   U186 : ADFULD1 port map( A => n262, B => n237, CI => n235, CO => n232, S => 
                           n233);
   U187 : ADFULD1 port map( A => n239, B => n266, CI => n264, CO => n234, S => 
                           n235);
   U188 : ADFULD1 port map( A => n268, B => n243, CI => n241, CO => n236, S => 
                           n237);
   U189 : ADFULD1 port map( A => n270, B => n247, CI => n245, CO => n238, S => 
                           n239);
   U190 : ADFULD1 port map( A => n274, B => n249, CI => n272, CO => n240, S => 
                           n241);
   U191 : ADFULD1 port map( A => n253, B => n255, CI => n257, CO => n242, S => 
                           n243);
   U192 : ADFULD1 port map( A => n280, B => n276, CI => n251, CO => n244, S => 
                           n245);
   U193 : ADFULD1 port map( A => n278, B => n284, CI => n282, CO => n246, S => 
                           n247);
   U194 : ADFULD1 port map( A => n1047, B => n1013, CI => n259, CO => n248, S 
                           => n249);
   U195 : ADFULD1 port map( A => n977, B => n1067, CI => n999, CO => n250, S =>
                           n251);
   U196 : ADFULD1 port map( A => n959, B => n969, CI => n963, CO => n252, S => 
                           n253);
   U197 : ADFULD1 port map( A => n1113, B => n987, CI => n1089, CO => n254, S 
                           => n255);
   U198 : ADFULD1 port map( A => n1167, B => n1029, CI => n1139, CO => n256, S 
                           => n257);
   U199 : ADHALFDL port map( A => n286, B => n1197, CO => n258, S => n259);
   U200 : ADFULD1 port map( A => n290, B => n265, CI => n263, CO => n260, S => 
                           n261);
   U201 : ADFULD1 port map( A => n267, B => n294, CI => n292, CO => n262, S => 
                           n263);
   U202 : ADFULD1 port map( A => n296, B => n271, CI => n269, CO => n264, S => 
                           n265);
   U203 : ADFULD1 port map( A => n275, B => n298, CI => n273, CO => n266, S => 
                           n267);
   U204 : ADFULD1 port map( A => n302, B => n281, CI => n300, CO => n268, S => 
                           n269);
   U205 : ADFULD1 port map( A => n283, B => n277, CI => n279, CO => n270, S => 
                           n271);
   U206 : ADFULD1 port map( A => n310, B => n308, CI => n285, CO => n272, S => 
                           n273);
   U207 : ADFULD1 port map( A => n304, B => n312, CI => n306, CO => n274, S => 
                           n275);
   U208 : ADFULD1 port map( A => n1014, B => n1068, CI => n1048, CO => n276, S 
                           => n277);
   U209 : ADFULD1 port map( A => n978, B => n1090, CI => n988, CO => n278, S =>
                           n279);
   U210 : ADFULD1 port map( A => n964, B => n1114, CI => n970, CO => n280, S =>
                           n281);
   U211 : ADFULD1 port map( A => n1140, B => n1000, CI => n287, CO => n282, S 
                           => n283);
   U212 : ADFULD1 port map( A => n1030, B => n960, CI => n1168, CO => n284, S 
                           => n285);
   U213 : ADHALFDL port map( A => n1198, B => n940, CO => n286, S => n287);
   U214 : ADFULD1 port map( A => n316, B => n293, CI => n291, CO => n288, S => 
                           n289);
   U215 : ADFULD1 port map( A => n318, B => n297, CI => n295, CO => n290, S => 
                           n291);
   U216 : ADFULD1 port map( A => n299, B => n322, CI => n320, CO => n292, S => 
                           n293);
   U217 : ADFULD1 port map( A => n324, B => n303, CI => n301, CO => n294, S => 
                           n295);
   U218 : ADFULD1 port map( A => n307, B => n309, CI => n326, CO => n296, S => 
                           n297);
   U219 : ADFULD1 port map( A => n305, B => n328, CI => n311, CO => n298, S => 
                           n299);
   U220 : ADFULD1 port map( A => n332, B => n330, CI => n334, CO => n300, S => 
                           n301);
   U221 : ADFULD1 port map( A => n313, B => n1091, CI => n336, CO => n302, S =>
                           n303);
   U222 : ADFULD1 port map( A => n1015, B => n1115, CI => n1069, CO => n304, S 
                           => n305);
   U223 : ADFULD1 port map( A => n1141, B => n1001, CI => n989, CO => n306, S 
                           => n307);
   U224 : ADFULD1 port map( A => n979, B => n1049, CI => n1169, CO => n308, S 
                           => n309);
   U225 : ADFULD1 port map( A => n965, B => n1031, CI => n971, CO => n310, S =>
                           n311);
   U226 : ADHALFDL port map( A => n338, B => n1199, CO => n312, S => n313);
   U227 : ADFULD1 port map( A => n342, B => n319, CI => n317, CO => n314, S => 
                           n315);
   U228 : ADFULD1 port map( A => n344, B => n346, CI => n321, CO => n316, S => 
                           n317);
   U229 : ADFULD1 port map( A => n325, B => n327, CI => n323, CO => n318, S => 
                           n319);
   U230 : ADFULD1 port map( A => n350, B => n352, CI => n348, CO => n320, S => 
                           n321);
   U231 : ADFULD1 port map( A => n333, B => n335, CI => n329, CO => n322, S => 
                           n323);
   U232 : ADFULD1 port map( A => n337, B => n358, CI => n331, CO => n324, S => 
                           n325);
   U233 : ADFULD1 port map( A => n354, B => n360, CI => n356, CO => n326, S => 
                           n327);
   U234 : ADFULD1 port map( A => n1092, B => n1116, CI => n362, CO => n328, S 
                           => n329);
   U235 : ADFULD1 port map( A => n1016, B => n1142, CI => n1070, CO => n330, S 
                           => n331);
   U236 : ADFULD1 port map( A => n990, B => n1170, CI => n1002, CO => n332, S 
                           => n333);
   U237 : ADFULD1 port map( A => n980, B => n1032, CI => n339, CO => n334, S =>
                           n335);
   U238 : ADFULD1 port map( A => n1050, B => n966, CI => n972, CO => n336, S =>
                           n337);
   U239 : ADHALFDL port map( A => n1200, B => n941, CO => n338, S => n339);
   U240 : ADFULD1 port map( A => n366, B => n345, CI => n343, CO => n340, S => 
                           n341);
   U241 : ADFULD1 port map( A => n347, B => n370, CI => n368, CO => n342, S => 
                           n343);
   U242 : ADFULD1 port map( A => n351, B => n372, CI => n349, CO => n344, S => 
                           n345);
   U243 : ADFULD1 port map( A => n374, B => n376, CI => n353, CO => n346, S => 
                           n347);
   U244 : ADFULD1 port map( A => n361, B => n357, CI => n359, CO => n348, S => 
                           n349);
   U245 : ADFULD1 port map( A => n378, B => n380, CI => n355, CO => n350, S => 
                           n351);
   U246 : ADFULD1 port map( A => n384, B => n363, CI => n382, CO => n352, S => 
                           n353);
   U247 : ADFULD1 port map( A => n1033, B => n1093, CI => n1071, CO => n354, S 
                           => n355);
   U248 : ADFULD1 port map( A => n991, B => n1117, CI => n1017, CO => n356, S 
                           => n357);
   U249 : ADFULD1 port map( A => n973, B => n1003, CI => n981, CO => n358, S =>
                           n359);
   U250 : ADFULD1 port map( A => n1171, B => n1051, CI => n1143, CO => n360, S 
                           => n361);
   U251 : ADHALFDL port map( A => n386, B => n1201, CO => n362, S => n363);
   U252 : ADFULD1 port map( A => n390, B => n369, CI => n367, CO => n364, S => 
                           n365);
   U253 : ADFULD1 port map( A => n371, B => n394, CI => n392, CO => n366, S => 
                           n367);
   U254 : ADFULD1 port map( A => n375, B => n396, CI => n373, CO => n368, S => 
                           n369);
   U255 : ADFULD1 port map( A => n398, B => n400, CI => n377, CO => n370, S => 
                           n371);
   U256 : ADFULD1 port map( A => n383, B => n379, CI => n381, CO => n372, S => 
                           n373);
   U257 : ADFULD1 port map( A => n402, B => n404, CI => n385, CO => n374, S => 
                           n375);
   U258 : ADFULD1 port map( A => n408, B => n1072, CI => n406, CO => n376, S =>
                           n377);
   U259 : ADFULD1 port map( A => n1004, B => n1094, CI => n1034, CO => n378, S 
                           => n379);
   U260 : ADFULD1 port map( A => n992, B => n1144, CI => n1118, CO => n380, S 
                           => n381);
   U261 : ADFULD1 port map( A => n982, B => n1018, CI => n387, CO => n382, S =>
                           n383);
   U262 : ADFULD1 port map( A => n1052, B => n974, CI => n1172, CO => n384, S 
                           => n385);
   U263 : ADHALFDL port map( A => n1202, B => n942, CO => n386, S => n387);
   U264 : ADFULD1 port map( A => n412, B => n393, CI => n391, CO => n388, S => 
                           n389);
   U265 : ADFULD1 port map( A => n395, B => n397, CI => n414, CO => n390, S => 
                           n391);
   U266 : ADFULD1 port map( A => n399, B => n418, CI => n416, CO => n392, S => 
                           n393);
   U267 : ADFULD1 port map( A => n401, B => n407, CI => n420, CO => n394, S => 
                           n395);
   U268 : ADFULD1 port map( A => n403, B => n424, CI => n405, CO => n396, S => 
                           n397);
   U269 : ADFULD1 port map( A => n426, B => n428, CI => n422, CO => n398, S => 
                           n399);
   U270 : ADFULD1 port map( A => n1073, B => n1095, CI => n409, CO => n400, S 
                           => n401);
   U271 : ADFULD1 port map( A => n1005, B => n1119, CI => n1019, CO => n402, S 
                           => n403);
   U272 : ADFULD1 port map( A => n1173, B => n1035, CI => n1145, CO => n404, S 
                           => n405);
   U273 : ADFULD1 port map( A => n983, B => n1053, CI => n993, CO => n406, S =>
                           n407);
   U274 : ADHALFDL port map( A => n430, B => n1203, CO => n408, S => n409);
   U275 : ADFULD1 port map( A => n434, B => n415, CI => n413, CO => n410, S => 
                           n411);
   U276 : ADFULD1 port map( A => n417, B => n419, CI => n436, CO => n412, S => 
                           n413);
   U277 : ADFULD1 port map( A => n421, B => n440, CI => n438, CO => n414, S => 
                           n415);
   U278 : ADFULD1 port map( A => n427, B => n425, CI => n442, CO => n416, S => 
                           n417);
   U279 : ADFULD1 port map( A => n429, B => n444, CI => n423, CO => n418, S => 
                           n419);
   U280 : ADFULD1 port map( A => n448, B => n450, CI => n446, CO => n420, S => 
                           n421);
   U281 : ADFULD1 port map( A => n1074, B => n1120, CI => n1096, CO => n422, S 
                           => n423);
   U282 : ADFULD1 port map( A => n1006, B => n1146, CI => n1020, CO => n424, S 
                           => n425);
   U283 : ADFULD1 port map( A => n1174, B => n1036, CI => n431, CO => n426, S 
                           => n427);
   U284 : ADFULD1 port map( A => n1054, B => n984, CI => n994, CO => n428, S =>
                           n429);
   U285 : ADHALFDL port map( A => n1204, B => n943, CO => n430, S => n431);
   U286 : ADFULD1 port map( A => n454, B => n437, CI => n435, CO => n432, S => 
                           n433);
   U287 : ADFULD1 port map( A => n439, B => n441, CI => n456, CO => n434, S => 
                           n435);
   U288 : ADFULD1 port map( A => n443, B => n460, CI => n458, CO => n436, S => 
                           n437);
   U289 : ADFULD1 port map( A => n449, B => n445, CI => n447, CO => n438, S => 
                           n439);
   U290 : ADFULD1 port map( A => n464, B => n466, CI => n462, CO => n440, S => 
                           n441);
   U291 : ADFULD1 port map( A => n451, B => n1037, CI => n468, CO => n442, S =>
                           n443);
   U292 : ADFULD1 port map( A => n995, B => n1075, CI => n1007, CO => n444, S 
                           => n445);
   U293 : ADFULD1 port map( A => n1121, B => n1021, CI => n1097, CO => n446, S 
                           => n447);
   U294 : ADFULD1 port map( A => n1175, B => n1055, CI => n1147, CO => n448, S 
                           => n449);
   U295 : ADHALFDL port map( A => n470, B => n1205, CO => n450, S => n451);
   U296 : ADFULD1 port map( A => n474, B => n457, CI => n455, CO => n452, S => 
                           n453);
   U297 : ADFULD1 port map( A => n459, B => n461, CI => n476, CO => n454, S => 
                           n455);
   U298 : ADFULD1 port map( A => n480, B => n463, CI => n478, CO => n456, S => 
                           n457);
   U299 : ADFULD1 port map( A => n465, B => n469, CI => n467, CO => n458, S => 
                           n459);
   U300 : ADFULD1 port map( A => n482, B => n486, CI => n484, CO => n460, S => 
                           n461);
   U301 : ADFULD1 port map( A => n1098, B => n1122, CI => n488, CO => n462, S 
                           => n463);
   U302 : ADFULD1 port map( A => n1022, B => n1148, CI => n1056, CO => n464, S 
                           => n465);
   U303 : ADFULD1 port map( A => n1008, B => n1038, CI => n471, CO => n466, S 
                           => n467);
   U304 : ADFULD1 port map( A => n1076, B => n996, CI => n1176, CO => n468, S 
                           => n469);
   U305 : ADHALFDL port map( A => n1206, B => n944, CO => n470, S => n471);
   U306 : ADFULD1 port map( A => n492, B => n477, CI => n475, CO => n472, S => 
                           n473);
   U307 : ADFULD1 port map( A => n479, B => n481, CI => n494, CO => n474, S => 
                           n475);
   U308 : ADFULD1 port map( A => n498, B => n487, CI => n496, CO => n476, S => 
                           n477);
   U309 : ADFULD1 port map( A => n483, B => n500, CI => n485, CO => n478, S => 
                           n479);
   U310 : ADFULD1 port map( A => n504, B => n489, CI => n502, CO => n480, S => 
                           n481);
   U311 : ADFULD1 port map( A => n1057, B => n1149, CI => n1123, CO => n482, S 
                           => n483);
   U312 : ADFULD1 port map( A => n1177, B => n1099, CI => n1039, CO => n484, S 
                           => n485);
   U313 : ADFULD1 port map( A => n1009, B => n1077, CI => n1023, CO => n486, S 
                           => n487);
   U314 : ADHALFDL port map( A => n506, B => n1207, CO => n488, S => n489);
   U315 : ADFULD1 port map( A => n510, B => n495, CI => n493, CO => n490, S => 
                           n491);
   U316 : ADFULD1 port map( A => n497, B => n499, CI => n512, CO => n492, S => 
                           n493);
   U317 : ADFULD1 port map( A => n516, B => n503, CI => n514, CO => n494, S => 
                           n495);
   U318 : ADFULD1 port map( A => n505, B => n518, CI => n501, CO => n496, S => 
                           n497);
   U319 : ADFULD1 port map( A => n522, B => n1124, CI => n520, CO => n498, S =>
                           n499);
   U320 : ADFULD1 port map( A => n1040, B => n1150, CI => n1058, CO => n500, S 
                           => n501);
   U321 : ADFULD1 port map( A => n1178, B => n1100, CI => n507, CO => n502, S 
                           => n503);
   U322 : ADFULD1 port map( A => n1078, B => n1010, CI => n1024, CO => n504, S 
                           => n505);
   U323 : ADHALFDL port map( A => n1208, B => n945, CO => n506, S => n507);
   U324 : ADFULD1 port map( A => n526, B => n513, CI => n511, CO => n508, S => 
                           n509);
   U325 : ADFULD1 port map( A => n528, B => n530, CI => n515, CO => n510, S => 
                           n511);
   U326 : ADFULD1 port map( A => n521, B => n519, CI => n517, CO => n512, S => 
                           n513);
   U327 : ADFULD1 port map( A => n534, B => n536, CI => n532, CO => n514, S => 
                           n515);
   U328 : ADFULD1 port map( A => n1101, B => n1125, CI => n523, CO => n516, S 
                           => n517);
   U329 : ADFULD1 port map( A => n1025, B => n1041, CI => n1059, CO => n518, S 
                           => n519);
   U330 : ADFULD1 port map( A => n1179, B => n1079, CI => n1151, CO => n520, S 
                           => n521);
   U331 : ADHALFDL port map( A => n538, B => n1209, CO => n522, S => n523);
   U332 : ADFULD1 port map( A => n542, B => n529, CI => n527, CO => n524, S => 
                           n525);
   U333 : ADFULD1 port map( A => n544, B => n546, CI => n531, CO => n526, S => 
                           n527);
   U334 : ADFULD1 port map( A => n533, B => n537, CI => n535, CO => n528, S => 
                           n529);
   U335 : ADFULD1 port map( A => n550, B => n552, CI => n548, CO => n530, S => 
                           n531);
   U336 : ADFULD1 port map( A => n1080, B => n1152, CI => n1126, CO => n532, S 
                           => n533);
   U337 : ADFULD1 port map( A => n1042, B => n1060, CI => n539, CO => n534, S 
                           => n535);
   U338 : ADFULD1 port map( A => n1102, B => n1026, CI => n1180, CO => n536, S 
                           => n537);
   U339 : ADHALFDL port map( A => n1210, B => n946, CO => n538, S => n539);
   U340 : ADFULD1 port map( A => n556, B => n545, CI => n543, CO => n540, S => 
                           n541);
   U341 : ADFULD1 port map( A => n547, B => n551, CI => n558, CO => n542, S => 
                           n543);
   U342 : ADFULD1 port map( A => n560, B => n562, CI => n549, CO => n544, S => 
                           n545);
   U343 : ADFULD1 port map( A => n553, B => n1153, CI => n564, CO => n546, S =>
                           n547);
   U344 : ADFULD1 port map( A => n1181, B => n1081, CI => n1127, CO => n548, S 
                           => n549);
   U345 : ADFULD1 port map( A => n1043, B => n1103, CI => n1061, CO => n550, S 
                           => n551);
   U346 : ADHALFDL port map( A => n566, B => n1211, CO => n552, S => n553);
   U347 : ADFULD1 port map( A => n570, B => n559, CI => n557, CO => n554, S => 
                           n555);
   U348 : ADFULD1 port map( A => n561, B => n563, CI => n572, CO => n556, S => 
                           n557);
   U349 : ADFULD1 port map( A => n574, B => n576, CI => n565, CO => n558, S => 
                           n559);
   U350 : ADFULD1 port map( A => n1062, B => n1128, CI => n578, CO => n560, S 
                           => n561);
   U351 : ADFULD1 port map( A => n1154, B => n1082, CI => n567, CO => n562, S 
                           => n563);
   U352 : ADFULD1 port map( A => n1104, B => n1044, CI => n1182, CO => n564, S 
                           => n565);
   U353 : ADHALFDL port map( A => n1212, B => n947, CO => n566, S => n567);
   U354 : ADFULD1 port map( A => n582, B => n573, CI => n571, CO => n568, S => 
                           n569);
   U355 : ADFULD1 port map( A => n577, B => n575, CI => n584, CO => n570, S => 
                           n571);
   U356 : ADFULD1 port map( A => n588, B => n579, CI => n586, CO => n572, S => 
                           n573);
   U357 : ADFULD1 port map( A => n1063, B => n1129, CI => n1083, CO => n574, S 
                           => n575);
   U358 : ADFULD1 port map( A => n1183, B => n1105, CI => n1155, CO => n576, S 
                           => n577);
   U359 : ADHALFDL port map( A => n590, B => n1213, CO => n578, S => n579);
   U360 : ADFULD1 port map( A => n585, B => n594, CI => n583, CO => n580, S => 
                           n581);
   U361 : ADFULD1 port map( A => n587, B => n589, CI => n596, CO => n582, S => 
                           n583);
   U362 : ADFULD1 port map( A => n600, B => n1106, CI => n598, CO => n584, S =>
                           n585);
   U363 : ADFULD1 port map( A => n1084, B => n1156, CI => n591, CO => n586, S 
                           => n587);
   U364 : ADFULD1 port map( A => n1130, B => n1064, CI => n1184, CO => n588, S 
                           => n589);
   U365 : ADHALFDL port map( A => n1214, B => n948, CO => n590, S => n591);
   U366 : ADFULD1 port map( A => n604, B => n597, CI => n595, CO => n592, S => 
                           n593);
   U367 : ADFULD1 port map( A => n606, B => n608, CI => n599, CO => n594, S => 
                           n595);
   U368 : ADFULD1 port map( A => n1107, B => n1157, CI => n601, CO => n596, S 
                           => n597);
   U369 : ADFULD1 port map( A => n1085, B => n1131, CI => n1185, CO => n598, S 
                           => n599);
   U370 : ADHALFDL port map( A => n610, B => n1215, CO => n600, S => n601);
   U371 : ADFULD1 port map( A => n614, B => n607, CI => n605, CO => n602, S => 
                           n603);
   U372 : ADFULD1 port map( A => n616, B => n618, CI => n609, CO => n604, S => 
                           n605);
   U373 : ADFULD1 port map( A => n1108, B => n1158, CI => n611, CO => n606, S 
                           => n607);
   U374 : ADFULD1 port map( A => n1132, B => n1086, CI => n1186, CO => n608, S 
                           => n609);
   U375 : ADHALFDL port map( A => n1216, B => n949, CO => n610, S => n611);
   U376 : ADFULD1 port map( A => n617, B => n622, CI => n615, CO => n612, S => 
                           n613);
   U377 : ADFULD1 port map( A => n619, B => n1187, CI => n624, CO => n614, S =>
                           n615);
   U378 : ADFULD1 port map( A => n1109, B => n1133, CI => n1159, CO => n616, S 
                           => n617);
   U379 : ADHALFDL port map( A => n626, B => n1217, CO => n618, S => n619);
   U380 : ADFULD1 port map( A => n625, B => n630, CI => n623, CO => n620, S => 
                           n621);
   U381 : ADFULD1 port map( A => n627, B => n1160, CI => n632, CO => n622, S =>
                           n623);
   U382 : ADFULD1 port map( A => n1188, B => n1110, CI => n1134, CO => n624, S 
                           => n625);
   U383 : ADHALFDL port map( A => n1218, B => n950, CO => n626, S => n627);
   U384 : ADFULD1 port map( A => n636, B => n633, CI => n631, CO => n628, S => 
                           n629);
   U385 : ADFULD1 port map( A => n1135, B => n1189, CI => n1161, CO => n630, S 
                           => n631);
   U386 : ADHALFDL port map( A => n638, B => n1219, CO => n632, S => n633);
   U387 : ADFULD1 port map( A => n642, B => n639, CI => n637, CO => n634, S => 
                           n635);
   U388 : ADFULD1 port map( A => n1190, B => n1136, CI => n1162, CO => n636, S 
                           => n637);
   U389 : ADHALFDL port map( A => n1220, B => n951, CO => n638, S => n639);
   U390 : ADFULD1 port map( A => n1163, B => n1191, CI => n643, CO => n640, S 
                           => n641);
   U391 : ADHALFDL port map( A => n646, B => n1221, CO => n642, S => n643);
   U392 : ADFULD1 port map( A => n1192, B => n1164, CI => n647, CO => n644, S 
                           => n645);
   U393 : ADHALFDL port map( A => n1222, B => n952, CO => n646, S => n647);
   U394 : ADHALFDL port map( A => n650, B => n1223, CO => n648, S => n649);
   U395 : ADHALFDL port map( A => n1224, B => n953, CO => n650, S => n651);
   U397 : MUXB2DL port map( A0 => n104, A1 => n1420, SL => n652, Z => n955);
   U399 : MUXB2DL port map( A0 => n104, A1 => n1420, SL => n653, Z => n956);
   U402 : MUXB2DL port map( A0 => n99, A1 => n1419, SL => n654, Z => n957);
   U404 : MUXB2DL port map( A0 => n99, A1 => n1419, SL => n655, Z => n958);
   U406 : MUXB2DL port map( A0 => n99, A1 => n1419, SL => n656, Z => n959);
   U408 : MUXB2DL port map( A0 => n99, A1 => n1419, SL => n657, Z => n960);
   U411 : MUXB2DL port map( A0 => n94, A1 => n1416, SL => n658, Z => n961);
   U413 : MUXB2DL port map( A0 => n94, A1 => n1416, SL => n659, Z => n962);
   U415 : MUXB2DL port map( A0 => n94, A1 => n1416, SL => n660, Z => n963);
   U417 : MUXB2DL port map( A0 => n94, A1 => n1416, SL => n661, Z => n964);
   U419 : MUXB2DL port map( A0 => n94, A1 => n1416, SL => n662, Z => n965);
   U421 : MUXB2DL port map( A0 => n94, A1 => n1416, SL => n663, Z => n966);
   U424 : MUXB2DL port map( A0 => n89, A1 => n1414, SL => n664, Z => n967);
   U426 : MUXB2DL port map( A0 => n89, A1 => n1414, SL => n665, Z => n968);
   U428 : MUXB2DL port map( A0 => n89, A1 => n1414, SL => n666, Z => n969);
   U430 : MUXB2DL port map( A0 => n89, A1 => n1414, SL => n667, Z => n970);
   U432 : MUXB2DL port map( A0 => n89, A1 => n1414, SL => n668, Z => n971);
   U434 : MUXB2DL port map( A0 => n89, A1 => n1414, SL => n669, Z => n972);
   U436 : MUXB2DL port map( A0 => n89, A1 => n1414, SL => n670, Z => n973);
   U438 : MUXB2DL port map( A0 => n89, A1 => n1414, SL => n671, Z => n974);
   U441 : MUXB2DL port map( A0 => n84, A1 => n1412, SL => n672, Z => n975);
   U443 : MUXB2DL port map( A0 => n84, A1 => n1412, SL => n673, Z => n976);
   U445 : MUXB2DL port map( A0 => n84, A1 => n1412, SL => n674, Z => n977);
   U447 : MUXB2DL port map( A0 => n84, A1 => n1412, SL => n675, Z => n978);
   U449 : MUXB2DL port map( A0 => n84, A1 => n1412, SL => n676, Z => n979);
   U451 : MUXB2DL port map( A0 => n84, A1 => n1412, SL => n677, Z => n980);
   U453 : MUXB2DL port map( A0 => n84, A1 => n1412, SL => n678, Z => n981);
   U455 : MUXB2DL port map( A0 => n84, A1 => n1412, SL => n679, Z => n982);
   U457 : MUXB2DL port map( A0 => n84, A1 => n1412, SL => n680, Z => n983);
   U459 : MUXB2DL port map( A0 => n84, A1 => n1412, SL => n681, Z => n984);
   U462 : MUXB2DL port map( A0 => n80, A1 => n1410, SL => n682, Z => n985);
   U464 : MUXB2DL port map( A0 => n80, A1 => n1410, SL => n683, Z => n986);
   U466 : MUXB2DL port map( A0 => n80, A1 => n1410, SL => n684, Z => n987);
   U468 : MUXB2DL port map( A0 => n80, A1 => n1410, SL => n685, Z => n988);
   U470 : MUXB2DL port map( A0 => n80, A1 => n1410, SL => n686, Z => n989);
   U472 : MUXB2DL port map( A0 => n80, A1 => n1410, SL => n687, Z => n990);
   U474 : MUXB2DL port map( A0 => n80, A1 => n1410, SL => n688, Z => n991);
   U476 : MUXB2DL port map( A0 => n80, A1 => n1410, SL => n689, Z => n992);
   U478 : MUXB2DL port map( A0 => n80, A1 => n1410, SL => n690, Z => n993);
   U480 : MUXB2DL port map( A0 => n80, A1 => n1410, SL => n691, Z => n994);
   U482 : MUXB2DL port map( A0 => n80, A1 => n1410, SL => n692, Z => n995);
   U484 : MUXB2DL port map( A0 => n80, A1 => n1410, SL => n693, Z => n996);
   U487 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n694, Z => n997);
   U489 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n695, Z => n998);
   U491 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n696, Z => n999);
   U493 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n697, Z => n1000);
   U495 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n698, Z => n1001);
   U497 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n699, Z => n1002);
   U499 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n700, Z => n1003);
   U501 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n701, Z => n1004);
   U503 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n702, Z => n1005);
   U505 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n703, Z => n1006);
   U507 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n704, Z => n1007);
   U509 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n705, Z => n1008);
   U511 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n706, Z => n1009);
   U513 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n707, Z => n1010);
   U516 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n708, Z => n1011);
   U518 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n709, Z => n1012);
   U520 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n710, Z => n1013);
   U522 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n711, Z => n1014);
   U524 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n712, Z => n1015);
   U526 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n713, Z => n1016);
   U528 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n714, Z => n1017);
   U530 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n715, Z => n1018);
   U532 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n716, Z => n1019);
   U534 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n717, Z => n1020);
   U536 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n718, Z => n1021);
   U538 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n719, Z => n1022);
   U540 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n720, Z => n1023);
   U542 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n721, Z => n1024);
   U544 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n722, Z => n1025);
   U546 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n723, Z => n1026);
   U549 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n724, Z => n1027);
   U551 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n725, Z => n1028);
   U553 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n726, Z => n1029);
   U555 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n727, Z => n1030);
   U557 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n728, Z => n1031);
   U559 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n729, Z => n1032);
   U561 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n730, Z => n1033);
   U563 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n731, Z => n1034);
   U565 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n732, Z => n1035);
   U567 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n733, Z => n1036);
   U569 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n734, Z => n1037);
   U571 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n735, Z => n1038);
   U573 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n736, Z => n1039);
   U575 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n737, Z => n1040);
   U577 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n738, Z => n1041);
   U579 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n739, Z => n1042);
   U581 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n740, Z => n1043);
   U583 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n741, Z => n1044);
   U586 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n742, Z => n1045);
   U588 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n743, Z => n1046);
   U590 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n744, Z => n1047);
   U592 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n745, Z => n1048);
   U594 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n746, Z => n1049);
   U596 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n747, Z => n1050);
   U598 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n748, Z => n1051);
   U600 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n749, Z => n1052);
   U602 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n750, Z => n1053);
   U604 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n751, Z => n1054);
   U606 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n752, Z => n1055);
   U608 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n753, Z => n1056);
   U610 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n754, Z => n1057);
   U612 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n755, Z => n1058);
   U614 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n756, Z => n1059);
   U616 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n757, Z => n1060);
   U618 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n758, Z => n1061);
   U620 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n759, Z => n1062);
   U622 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n760, Z => n1063);
   U624 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n761, Z => n1064);
   U627 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n762, Z => n1065);
   U629 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n763, Z => n1066);
   U631 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n764, Z => n1067);
   U633 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n765, Z => n1068);
   U635 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n766, Z => n1069);
   U637 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n767, Z => n1070);
   U639 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n768, Z => n1071);
   U641 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n769, Z => n1072);
   U643 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n770, Z => n1073);
   U645 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n771, Z => n1074);
   U647 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n772, Z => n1075);
   U649 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n773, Z => n1076);
   U651 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n774, Z => n1077);
   U653 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n775, Z => n1078);
   U655 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n776, Z => n1079);
   U657 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n777, Z => n1080);
   U659 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n778, Z => n1081);
   U661 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n779, Z => n1082);
   U663 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n780, Z => n1083);
   U665 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n781, Z => n1084);
   U667 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n782, Z => n1085);
   U669 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n783, Z => n1086);
   U672 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n784, Z => n1087);
   U674 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n785, Z => n1088);
   U676 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n786, Z => n1089);
   U678 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n787, Z => n1090);
   U680 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n788, Z => n1091);
   U682 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n789, Z => n1092);
   U684 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n790, Z => n1093);
   U686 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n791, Z => n1094);
   U688 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n792, Z => n1095);
   U690 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n793, Z => n1096);
   U692 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n794, Z => n1097);
   U694 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n795, Z => n1098);
   U696 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n796, Z => n1099);
   U698 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n797, Z => n1100);
   U700 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n798, Z => n1101);
   U702 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n799, Z => n1102);
   U704 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n800, Z => n1103);
   U706 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n801, Z => n1104);
   U708 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n802, Z => n1105);
   U710 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n803, Z => n1106);
   U712 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n804, Z => n1107);
   U714 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n805, Z => n1108);
   U716 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n806, Z => n1109);
   U718 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n807, Z => n1110);
   U721 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n808, Z => n1111);
   U723 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n809, Z => n1112);
   U725 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n810, Z => n1113);
   U727 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n811, Z => n1114);
   U729 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n812, Z => n1115);
   U731 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n813, Z => n1116);
   U733 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n814, Z => n1117);
   U735 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n815, Z => n1118);
   U737 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n816, Z => n1119);
   U739 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n817, Z => n1120);
   U741 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n818, Z => n1121);
   U743 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n819, Z => n1122);
   U745 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n820, Z => n1123);
   U747 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n821, Z => n1124);
   U749 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n822, Z => n1125);
   U751 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n823, Z => n1126);
   U753 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n824, Z => n1127);
   U755 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n825, Z => n1128);
   U757 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n826, Z => n1129);
   U759 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n827, Z => n1130);
   U761 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n828, Z => n1131);
   U763 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n829, Z => n1132);
   U765 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n830, Z => n1133);
   U767 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n831, Z => n1134);
   U769 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n832, Z => n1135);
   U771 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n833, Z => n1136);
   U774 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n834, Z => n1137);
   U776 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n835, Z => n1138);
   U778 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n836, Z => n1139);
   U780 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n837, Z => n1140);
   U782 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n838, Z => n1141);
   U784 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n839, Z => n1142);
   U786 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n840, Z => n1143);
   U788 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n841, Z => n1144);
   U790 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n842, Z => n1145);
   U792 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n843, Z => n1146);
   U794 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n844, Z => n1147);
   U796 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n845, Z => n1148);
   U798 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n846, Z => n1149);
   U800 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n847, Z => n1150);
   U802 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n848, Z => n1151);
   U804 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n849, Z => n1152);
   U806 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n850, Z => n1153);
   U808 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n851, Z => n1154);
   U810 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n852, Z => n1155);
   U812 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n853, Z => n1156);
   U814 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n854, Z => n1157);
   U816 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n855, Z => n1158);
   U818 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n856, Z => n1159);
   U820 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n857, Z => n1160);
   U822 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n858, Z => n1161);
   U824 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n859, Z => n1162);
   U826 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n860, Z => n1163);
   U828 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n861, Z => n1164);
   U831 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n862, Z => n1165);
   U833 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n863, Z => n1166);
   U835 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n864, Z => n1167);
   U837 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n865, Z => n1168);
   U839 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n866, Z => n1169);
   U841 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n867, Z => n1170);
   U843 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n868, Z => n1171);
   U845 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n869, Z => n1172);
   U847 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n870, Z => n1173);
   U849 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n871, Z => n1174);
   U851 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n872, Z => n1175);
   U853 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n873, Z => n1176);
   U855 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n874, Z => n1177);
   U857 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n875, Z => n1178);
   U859 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n876, Z => n1179);
   U861 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n877, Z => n1180);
   U863 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n878, Z => n1181);
   U865 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n879, Z => n1182);
   U867 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n880, Z => n1183);
   U869 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n881, Z => n1184);
   U871 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n882, Z => n1185);
   U873 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n883, Z => n1186);
   U875 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n884, Z => n1187);
   U877 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n885, Z => n1188);
   U879 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n886, Z => n1189);
   U881 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n887, Z => n1190);
   U883 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n888, Z => n1191);
   U885 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n889, Z => n1192);
   U887 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n890, Z => n1193);
   U889 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n891, Z => n1194);
   U892 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n892, Z => n1195);
   U894 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n893, Z => n1196);
   U896 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n894, Z => n1197);
   U898 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n895, Z => n1198);
   U900 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n896, Z => n1199);
   U902 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n897, Z => n1200);
   U904 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n898, Z => n1201);
   U906 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n899, Z => n1202);
   U908 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n900, Z => n1203);
   U910 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n901, Z => n1204);
   U912 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n902, Z => n1205);
   U914 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n903, Z => n1206);
   U916 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n904, Z => n1207);
   U918 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n905, Z => n1208);
   U920 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n906, Z => n1209);
   U922 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n907, Z => n1210);
   U924 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n908, Z => n1211);
   U926 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n909, Z => n1212);
   U928 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n910, Z => n1213);
   U930 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n911, Z => n1214);
   U932 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n912, Z => n1215);
   U934 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n913, Z => n1216);
   U936 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n914, Z => n1217);
   U938 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n915, Z => n1218);
   U940 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n916, Z => n1219);
   U942 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n917, Z => n1220);
   U944 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n918, Z => n1221);
   U946 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n919, Z => n1222);
   U948 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n920, Z => n1223);
   U950 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n921, Z => n1224);
   U952 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n922, Z => n1225);
   U954 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n923, Z => n1226);
   U1021 : NAN2D1 port map( A1 => n1390, A2 => n1392, Z => n1375);
   U1022 : OAI21D1 port map( A1 => a(2), A2 => a(1), B => n1395, Z => n1376);
   U1023 : OAI21D1 port map( A1 => a(4), A2 => a(3), B => n1397, Z => n1377);
   U1024 : EXOR2D1 port map( A1 => a(6), A2 => a(5), Z => n1378);
   U1025 : EXOR2D1 port map( A1 => a(8), A2 => a(7), Z => n1379);
   U1026 : OAI21D1 port map( A1 => a(6), A2 => a(5), B => n1399, Z => n1380);
   U1027 : OAI21D1 port map( A1 => a(8), A2 => a(7), B => n1401, Z => n1381);
   U1028 : INVD1 port map( A => n1382, Z => n1384);
   U1029 : INVD1 port map( A => n1383, Z => n1385);
   U1030 : INVD1 port map( A => n953, Z => n1393);
   U1031 : INVD1 port map( A => n952, Z => n1394);
   U1032 : INVD1 port map( A => n951, Z => n1396);
   U1033 : INVD1 port map( A => n950, Z => n1398);
   U1034 : INVD1 port map( A => n949, Z => n1400);
   U1035 : INVD1 port map( A => n948, Z => n1402);
   U1036 : INVD1 port map( A => n947, Z => n1404);
   U1037 : INVD1 port map( A => n946, Z => n1406);
   U1038 : INVD1 port map( A => n945, Z => n1408);
   U1039 : INVD1 port map( A => n944, Z => n1410);
   U1040 : INVD1 port map( A => n943, Z => n1412);
   U1041 : INVD1 port map( A => n942, Z => n1414);
   U1042 : INVD1 port map( A => n941, Z => n1416);
   U1043 : INVD1 port map( A => n940, Z => n1419);
   U1044 : INVD1 port map( A => n939, Z => n1420);
   U1045 : INVD1 port map( A => n1391, Z => n1390);
   U1046 : INVD1 port map( A => a(1), Z => n1392);
   U1047 : EXNOR2D1 port map( A1 => a(2), A2 => a(1), Z => n1382);
   U1048 : INVD1 port map( A => n1389, Z => n1388);
   U1049 : EXNOR2D1 port map( A1 => a(4), A2 => a(3), Z => n1383);
   U1050 : INVD1 port map( A => n1387, Z => n1386);
   U1051 : INVD1 port map( A => a(3), Z => n1395);
   U1052 : INVD1 port map( A => a(5), Z => n1397);
   U1053 : INVD1 port map( A => a(7), Z => n1399);
   U1054 : INVD1 port map( A => a(9), Z => n1401);
   U1055 : EXOR2D1 port map( A1 => a(10), A2 => a(9), Z => n1441);
   U1056 : INVD1 port map( A => a(11), Z => n1403);
   U1057 : OAI21D1 port map( A1 => a(9), A2 => a(10), B => n1403, Z => n42);
   U1058 : EXOR2D1 port map( A1 => a(12), A2 => a(11), Z => n1442);
   U1059 : INVD1 port map( A => a(13), Z => n1405);
   U1060 : OAI21D1 port map( A1 => a(12), A2 => a(11), B => n1405, Z => n50);
   U1061 : EXOR2D1 port map( A1 => a(14), A2 => a(13), Z => n1443);
   U1062 : INVD1 port map( A => a(15), Z => n1407);
   U1063 : OAI21D1 port map( A1 => a(14), A2 => a(13), B => n1407, Z => n58);
   U1064 : EXOR2D1 port map( A1 => a(16), A2 => a(15), Z => n1444);
   U1065 : INVD1 port map( A => a(17), Z => n1409);
   U1066 : OAI21D1 port map( A1 => a(16), A2 => a(15), B => n1409, Z => n66);
   U1067 : EXOR2D1 port map( A1 => a(18), A2 => a(17), Z => n1445);
   U1068 : INVD1 port map( A => a(19), Z => n1411);
   U1069 : OAI21D1 port map( A1 => a(18), A2 => a(17), B => n1411, Z => n73);
   U1070 : EXOR2D1 port map( A1 => a(20), A2 => a(19), Z => n1446);
   U1071 : INVD1 port map( A => a(21), Z => n1413);
   U1072 : OAI21D1 port map( A1 => a(20), A2 => a(19), B => n1413, Z => n80);
   U1073 : EXOR2D1 port map( A1 => a(22), A2 => a(21), Z => n1447);
   U1074 : INVD1 port map( A => a(23), Z => n1415);
   U1075 : OAI21D1 port map( A1 => a(22), A2 => a(21), B => n1415, Z => n84);
   U1076 : INVD1 port map( A => a(25), Z => n1417);
   U1077 : INVD1 port map( A => a(27), Z => n1418);
   U1078 : INVD1 port map( A => a(29), Z => n1421);
   U1079 : MUXB2DL port map( A0 => b(29), A1 => b(28), SL => n1382, Z => n862);
   U1080 : INVD1 port map( A => a(0), Z => n1391);
   U1081 : INVD1 port map( A => b(1), Z => n1389);
   U1082 : INVD1 port map( A => b(3), Z => n1387);
   U1083 : INVD1 port map( A => a(31), Z => n1422);
   U1084 : EXOR3D1 port map( A1 => n1423, A2 => n1424, A3 => n1425, Z => 
                           product(31));
   U1085 : EXOR3D1 port map( A1 => n208, A2 => n206, A3 => n1426, Z => n1425);
   U1086 : EXOR2D1 port map( A1 => n214, A2 => n212, Z => n1426);
   U1087 : EXOR2D1 port map( A1 => n202, A2 => n156, Z => n1424);
   U1088 : EXOR3D1 port map( A1 => n1427, A2 => n1428, A3 => n1429, Z => n1423)
                           ;
   U1089 : EXOR3D1 port map( A1 => n957, A2 => n955, A3 => n1430, Z => n1429);
   U1090 : EXNOR2D1 port map( A1 => n997, A2 => n975, Z => n1430);
   U1091 : EXOR3D1 port map( A1 => n1431, A2 => n204, A3 => n1432, Z => n1428);
   U1092 : EXOR3D1 port map( A1 => n1087, A2 => n1065, A3 => n1433, Z => n1432)
                           ;
   U1093 : EXNOR2D1 port map( A1 => n210, A2 => n1111, Z => n1433);
   U1094 : EXOR3D1 port map( A1 => n961, A2 => n218, A3 => n1434, Z => n1431);
   U1095 : EXOR2D1 port map( A1 => n985, A2 => n967, Z => n1434);
   U1096 : EXOR3D1 port map( A1 => n1435, A2 => n1436, A3 => n1437, Z => n1427)
                           ;
   U1097 : EXOR3D1 port map( A1 => n1027, A2 => n1011, A3 => n1438, Z => n1437)
                           ;
   U1098 : EXOR3D1 port map( A1 => n1165, A2 => n1137, A3 => n1045, Z => n1438)
                           ;
   U1099 : EXOR3D1 port map( A1 => n216, A2 => n1195, A3 => n1439, Z => n1436);
   U1100 : EXOR2D1 port map( A1 => n222, A2 => n220, Z => n1439);
   U1101 : EXOR3D1 port map( A1 => n226, A2 => n224, A3 => n1440, Z => n1435);
   U1102 : EXOR2D1 port map( A1 => n230, A2 => n228, Z => n1440);
   U1103 : OAI21D1 port map( A1 => a(28), A2 => a(27), B => n1421, Z => n99);
   U1104 : AOI21D1 port map( A1 => a(25), A2 => a(26), B => n1418, Z => n941);
   U1105 : OAI21D1 port map( A1 => a(26), A2 => a(25), B => n1418, Z => n94);
   U1106 : NAN2D1 port map( A1 => b(0), A2 => n1390, Z => n923);
   U1107 : MUXB2DL port map( A0 => b(0), A1 => n1388, SL => n1390, Z => n922);
   U1108 : MUXB2DL port map( A0 => n1388, A1 => b(2), SL => n1390, Z => n921);
   U1109 : MUXB2DL port map( A0 => b(2), A1 => n1386, SL => n1390, Z => n920);
   U1110 : MUXB2DL port map( A0 => n1386, A1 => b(4), SL => n1390, Z => n919);
   U1111 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1390, Z => n918);
   U1112 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1390, Z => n917);
   U1113 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1390, Z => n916);
   U1114 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1390, Z => n915);
   U1115 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1390, Z => n914);
   U1116 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1390, Z => n913);
   U1117 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1390, Z => n912);
   U1118 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1390, Z => n911);
   U1119 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1390, Z => n910);
   U1120 : AOI21D1 port map( A1 => a(23), A2 => a(24), B => n1417, Z => n942);
   U1121 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => a(0), Z => n909);
   U1122 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => a(0), Z => n908);
   U1123 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => a(0), Z => n907);
   U1124 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => a(0), Z => n906);
   U1125 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => a(0), Z => n905);
   U1126 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => a(0), Z => n904);
   U1127 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => a(0), Z => n903);
   U1128 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => a(0), Z => n902);
   U1129 : MUXB2DL port map( A0 => b(21), A1 => b(22), SL => a(0), Z => n901);
   U1130 : MUXB2DL port map( A0 => b(22), A1 => b(23), SL => a(0), Z => n900);
   U1131 : MUXB2DL port map( A0 => b(23), A1 => b(24), SL => a(0), Z => n899);
   U1132 : MUXB2DL port map( A0 => b(24), A1 => b(25), SL => a(0), Z => n898);
   U1133 : MUXB2DL port map( A0 => b(25), A1 => b(26), SL => a(0), Z => n897);
   U1134 : MUXB2DL port map( A0 => b(26), A1 => b(27), SL => a(0), Z => n896);
   U1135 : MUXB2DL port map( A0 => b(27), A1 => b(28), SL => a(0), Z => n895);
   U1136 : MUXB2DL port map( A0 => b(28), A1 => b(29), SL => a(0), Z => n894);
   U1137 : MUXB2DL port map( A0 => b(29), A1 => b(30), SL => a(0), Z => n893);
   U1138 : MUXB2DL port map( A0 => b(30), A1 => b(31), SL => n1390, Z => n892);
   U1139 : NAN2D1 port map( A1 => b(0), A2 => n1384, Z => n891);
   U1140 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1384, Z => n890);
   U1141 : OAI21D1 port map( A1 => a(24), A2 => a(23), B => n1417, Z => n89);
   U1142 : MUXB2DL port map( A0 => n1388, A1 => b(2), SL => n1384, Z => n889);
   U1143 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1384, Z => n888);
   U1144 : MUXB2DL port map( A0 => n1386, A1 => b(4), SL => n1384, Z => n887);
   U1145 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1384, Z => n886);
   U1146 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1384, Z => n885);
   U1147 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1384, Z => n884);
   U1148 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1384, Z => n883);
   U1149 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1384, Z => n882);
   U1150 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1384, Z => n881);
   U1151 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1384, Z => n880);
   U1152 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1384, Z => n879);
   U1153 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1384, Z => n878);
   U1154 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1384, Z => n877);
   U1155 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1384, Z => n876);
   U1156 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1384, Z => n875);
   U1157 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1384, Z => n874);
   U1158 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1384, Z => n873);
   U1159 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1384, Z => n872);
   U1160 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => n1384, Z => n871);
   U1161 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => n1384, Z => n870);
   U1162 : MUXB2DL port map( A0 => b(21), A1 => b(22), SL => n1384, Z => n869);
   U1163 : MUXB2DL port map( A0 => b(22), A1 => b(23), SL => n1384, Z => n868);
   U1164 : MUXB2DL port map( A0 => b(23), A1 => b(24), SL => n1384, Z => n867);
   U1165 : MUXB2DL port map( A0 => b(24), A1 => b(25), SL => n1384, Z => n866);
   U1166 : MUXB2DL port map( A0 => b(25), A1 => b(26), SL => n1384, Z => n865);
   U1167 : MUXB2DL port map( A0 => b(26), A1 => b(27), SL => n1384, Z => n864);
   U1168 : MUXB2DL port map( A0 => b(27), A1 => b(28), SL => n1384, Z => n863);
   U1169 : NAN2D1 port map( A1 => b(0), A2 => n1385, Z => n861);
   U1170 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1385, Z => n860);
   U1171 : AOI21D1 port map( A1 => a(21), A2 => a(22), B => n1415, Z => n943);
   U1172 : MUXB2DL port map( A0 => n1388, A1 => b(2), SL => n1385, Z => n859);
   U1173 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1385, Z => n858);
   U1174 : MUXB2DL port map( A0 => n1386, A1 => b(4), SL => n1385, Z => n857);
   U1175 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1385, Z => n856);
   U1176 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1385, Z => n855);
   U1177 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1385, Z => n854);
   U1178 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1385, Z => n853);
   U1179 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1385, Z => n852);
   U1180 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1385, Z => n851);
   U1181 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1385, Z => n850);
   U1182 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1385, Z => n849);
   U1183 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1385, Z => n848);
   U1184 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1385, Z => n847);
   U1185 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1385, Z => n846);
   U1186 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1385, Z => n845);
   U1187 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1385, Z => n844);
   U1188 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1385, Z => n843);
   U1189 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1385, Z => n842);
   U1190 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => n1385, Z => n841);
   U1191 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => n1385, Z => n840);
   U1192 : MUXB2DL port map( A0 => b(21), A1 => b(22), SL => n1385, Z => n839);
   U1193 : MUXB2DL port map( A0 => b(22), A1 => b(23), SL => n1385, Z => n838);
   U1194 : MUXB2DL port map( A0 => b(23), A1 => b(24), SL => n1385, Z => n837);
   U1195 : MUXB2DL port map( A0 => b(24), A1 => b(25), SL => n1385, Z => n836);
   U1196 : MUXB2DL port map( A0 => b(25), A1 => b(26), SL => n1385, Z => n835);
   U1197 : MUXB2DL port map( A0 => b(26), A1 => b(27), SL => n1385, Z => n834);
   U1198 : NAN2D1 port map( A1 => b(0), A2 => n1378, Z => n833);
   U1199 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1378, Z => n832);
   U1200 : MUXB2DL port map( A0 => n1388, A1 => b(2), SL => n1378, Z => n831);
   U1201 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1378, Z => n830);
   U1202 : MUXB2DL port map( A0 => n1386, A1 => b(4), SL => n1378, Z => n829);
   U1203 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1378, Z => n828);
   U1204 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1378, Z => n827);
   U1205 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1378, Z => n826);
   U1206 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1378, Z => n825);
   U1207 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1378, Z => n824);
   U1208 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1378, Z => n823);
   U1209 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1378, Z => n822);
   U1210 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1378, Z => n821);
   U1211 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1378, Z => n820);
   U1212 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1378, Z => n819);
   U1213 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1378, Z => n818);
   U1214 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1378, Z => n817);
   U1215 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1378, Z => n816);
   U1216 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1378, Z => n815);
   U1217 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1378, Z => n814);
   U1218 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => n1378, Z => n813);
   U1219 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => n1378, Z => n812);
   U1220 : MUXB2DL port map( A0 => b(21), A1 => b(22), SL => n1378, Z => n811);
   U1221 : MUXB2DL port map( A0 => b(22), A1 => b(23), SL => n1378, Z => n810);
   U1222 : AOI21D1 port map( A1 => a(19), A2 => a(20), B => n1413, Z => n944);
   U1223 : MUXB2DL port map( A0 => b(23), A1 => b(24), SL => n1378, Z => n809);
   U1224 : MUXB2DL port map( A0 => b(24), A1 => b(25), SL => n1378, Z => n808);
   U1225 : NAN2D1 port map( A1 => b(0), A2 => n1379, Z => n807);
   U1226 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1379, Z => n806);
   U1227 : MUXB2DL port map( A0 => b(1), A1 => b(2), SL => n1379, Z => n805);
   U1228 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1379, Z => n804);
   U1229 : MUXB2DL port map( A0 => n1386, A1 => b(4), SL => n1379, Z => n803);
   U1230 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1379, Z => n802);
   U1231 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1379, Z => n801);
   U1232 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1379, Z => n800);
   U1233 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1379, Z => n799);
   U1234 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1379, Z => n798);
   U1235 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1379, Z => n797);
   U1236 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1379, Z => n796);
   U1237 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1379, Z => n795);
   U1238 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1379, Z => n794);
   U1239 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1379, Z => n793);
   U1240 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1379, Z => n792);
   U1241 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1379, Z => n791);
   U1242 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1379, Z => n790);
   U1243 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1379, Z => n789);
   U1244 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1379, Z => n788);
   U1245 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => n1379, Z => n787);
   U1246 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => n1379, Z => n786);
   U1247 : MUXB2DL port map( A0 => b(21), A1 => b(22), SL => n1379, Z => n785);
   U1248 : MUXB2DL port map( A0 => b(22), A1 => b(23), SL => n1379, Z => n784);
   U1249 : NAN2D1 port map( A1 => b(0), A2 => n1441, Z => n783);
   U1250 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1441, Z => n782);
   U1251 : MUXB2DL port map( A0 => n1388, A1 => b(2), SL => n1441, Z => n781);
   U1252 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1441, Z => n780);
   U1253 : MUXB2DL port map( A0 => b(3), A1 => b(4), SL => n1441, Z => n779);
   U1254 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1441, Z => n778);
   U1255 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1441, Z => n777);
   U1256 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1441, Z => n776);
   U1257 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1441, Z => n775);
   U1258 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1441, Z => n774);
   U1259 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1441, Z => n773);
   U1260 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1441, Z => n772);
   U1261 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1441, Z => n771);
   U1262 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1441, Z => n770);
   U1263 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1441, Z => n769);
   U1264 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1441, Z => n768);
   U1265 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1441, Z => n767);
   U1266 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1441, Z => n766);
   U1267 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1441, Z => n765);
   U1268 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1441, Z => n764);
   U1269 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => n1441, Z => n763);
   U1270 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => n1441, Z => n762);
   U1271 : NAN2D1 port map( A1 => b(0), A2 => n1442, Z => n761);
   U1272 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1442, Z => n760);
   U1273 : MUXB2DL port map( A0 => b(1), A1 => b(2), SL => n1442, Z => n759);
   U1274 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1442, Z => n758);
   U1275 : MUXB2DL port map( A0 => n1386, A1 => b(4), SL => n1442, Z => n757);
   U1276 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1442, Z => n756);
   U1277 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1442, Z => n755);
   U1278 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1442, Z => n754);
   U1279 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1442, Z => n753);
   U1280 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1442, Z => n752);
   U1281 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1442, Z => n751);
   U1282 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1442, Z => n750);
   U1283 : AOI21D1 port map( A1 => a(17), A2 => a(18), B => n1411, Z => n945);
   U1284 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1442, Z => n749);
   U1285 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1442, Z => n748);
   U1286 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1442, Z => n747);
   U1287 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1442, Z => n746);
   U1288 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1442, Z => n745);
   U1289 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1442, Z => n744);
   U1290 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1442, Z => n743);
   U1291 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1442, Z => n742);
   U1292 : NAN2D1 port map( A1 => b(0), A2 => n1443, Z => n741);
   U1293 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1443, Z => n740);
   U1294 : MUXB2DL port map( A0 => n1388, A1 => b(2), SL => n1443, Z => n739);
   U1295 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1443, Z => n738);
   U1296 : MUXB2DL port map( A0 => n1386, A1 => b(4), SL => n1443, Z => n737);
   U1297 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1443, Z => n736);
   U1298 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1443, Z => n735);
   U1299 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1443, Z => n734);
   U1300 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1443, Z => n733);
   U1301 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1443, Z => n732);
   U1302 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1443, Z => n731);
   U1303 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1443, Z => n730);
   U1304 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1443, Z => n729);
   U1305 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1443, Z => n728);
   U1306 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1443, Z => n727);
   U1307 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1443, Z => n726);
   U1308 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1443, Z => n725);
   U1309 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1443, Z => n724);
   U1310 : NAN2D1 port map( A1 => b(0), A2 => n1444, Z => n723);
   U1311 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1444, Z => n722);
   U1312 : MUXB2DL port map( A0 => n1388, A1 => b(2), SL => n1444, Z => n721);
   U1313 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1444, Z => n720);
   U1314 : MUXB2DL port map( A0 => n1386, A1 => b(4), SL => n1444, Z => n719);
   U1315 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1444, Z => n718);
   U1316 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1444, Z => n717);
   U1317 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1444, Z => n716);
   U1318 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1444, Z => n715);
   U1319 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1444, Z => n714);
   U1320 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1444, Z => n713);
   U1321 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1444, Z => n712);
   U1322 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1444, Z => n711);
   U1323 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1444, Z => n710);
   U1324 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1444, Z => n709);
   U1325 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1444, Z => n708);
   U1326 : NAN2D1 port map( A1 => b(0), A2 => n1445, Z => n707);
   U1327 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1445, Z => n706);
   U1328 : MUXB2DL port map( A0 => n1388, A1 => b(2), SL => n1445, Z => n705);
   U1329 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1445, Z => n704);
   U1330 : MUXB2DL port map( A0 => n1386, A1 => b(4), SL => n1445, Z => n703);
   U1331 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1445, Z => n702);
   U1332 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1445, Z => n701);
   U1333 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1445, Z => n700);
   U1334 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1445, Z => n699);
   U1335 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1445, Z => n698);
   U1336 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1445, Z => n697);
   U1337 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1445, Z => n696);
   U1338 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1445, Z => n695);
   U1339 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1445, Z => n694);
   U1340 : NAN2D1 port map( A1 => b(0), A2 => n1446, Z => n693);
   U1341 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1446, Z => n692);
   U1342 : MUXB2DL port map( A0 => n1388, A1 => b(2), SL => n1446, Z => n691);
   U1343 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1446, Z => n690);
   U1344 : MUXB2DL port map( A0 => n1386, A1 => b(4), SL => n1446, Z => n689);
   U1345 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1446, Z => n688);
   U1346 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1446, Z => n687);
   U1347 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1446, Z => n686);
   U1348 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1446, Z => n685);
   U1349 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1446, Z => n684);
   U1350 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1446, Z => n683);
   U1351 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1446, Z => n682);
   U1352 : NAN2D1 port map( A1 => b(0), A2 => n1447, Z => n681);
   U1353 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1447, Z => n680);
   U1354 : AOI21D1 port map( A1 => a(15), A2 => a(16), B => n1409, Z => n946);
   U1355 : MUXB2DL port map( A0 => n1388, A1 => b(2), SL => n1447, Z => n679);
   U1356 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1447, Z => n678);
   U1357 : MUXB2DL port map( A0 => n1386, A1 => b(4), SL => n1447, Z => n677);
   U1358 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1447, Z => n676);
   U1359 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1447, Z => n675);
   U1360 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1447, Z => n674);
   U1361 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1447, Z => n673);
   U1362 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1447, Z => n672);
   U1363 : NAN2D1 port map( A1 => b(0), A2 => n1448, Z => n671);
   U1364 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1448, Z => n670);
   U1365 : MUXB2DL port map( A0 => n1388, A1 => b(2), SL => n1448, Z => n669);
   U1366 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1448, Z => n668);
   U1367 : MUXB2DL port map( A0 => n1386, A1 => b(4), SL => n1448, Z => n667);
   U1368 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1448, Z => n666);
   U1369 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1448, Z => n665);
   U1370 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1448, Z => n664);
   U1371 : EXOR2D1 port map( A1 => a(24), A2 => a(23), Z => n1448);
   U1372 : NAN2D1 port map( A1 => b(0), A2 => n1449, Z => n663);
   U1373 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1449, Z => n662);
   U1374 : MUXB2DL port map( A0 => n1388, A1 => b(2), SL => n1449, Z => n661);
   U1375 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1449, Z => n660);
   U1376 : MUXB2DL port map( A0 => n1386, A1 => b(4), SL => n1449, Z => n659);
   U1377 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1449, Z => n658);
   U1378 : EXOR2D1 port map( A1 => a(26), A2 => a(25), Z => n1449);
   U1379 : NAN2D1 port map( A1 => b(0), A2 => n1450, Z => n657);
   U1380 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1450, Z => n656);
   U1381 : MUXB2DL port map( A0 => n1388, A1 => b(2), SL => n1450, Z => n655);
   U1382 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1450, Z => n654);
   U1383 : EXOR2D1 port map( A1 => a(28), A2 => a(27), Z => n1450);
   U1384 : NAN2D1 port map( A1 => b(0), A2 => n1451, Z => n653);
   U1385 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1451, Z => n652);
   U1386 : EXOR2D1 port map( A1 => a(30), A2 => a(29), Z => n1451);
   U1387 : AOI21D1 port map( A1 => a(13), A2 => a(14), B => n1407, Z => n947);
   U1388 : AOI21D1 port map( A1 => a(11), A2 => a(12), B => n1405, Z => n948);
   U1389 : AOI21D1 port map( A1 => a(9), A2 => a(10), B => n1403, Z => n949);
   U1390 : AOI21D1 port map( A1 => a(7), A2 => a(8), B => n1401, Z => n950);
   U1391 : AOI21D1 port map( A1 => a(5), A2 => a(6), B => n1399, Z => n951);
   U1392 : AOI21D1 port map( A1 => a(3), A2 => a(4), B => n1397, Z => n952);
   U1393 : AOI21D1 port map( A1 => a(1), A2 => a(2), B => n1395, Z => n953);
   U1394 : AOI21D1 port map( A1 => a(29), A2 => a(30), B => n1422, Z => n939);
   U1395 : OAI21D1 port map( A1 => a(30), A2 => a(29), B => n1422, Z => n104);
   U1396 : AOI21D1 port map( A1 => a(27), A2 => a(28), B => n1421, Z => n940);

end hier_filter_none_20;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_gp_custom.all;

architecture hier_filter_none_20 of gp_custom_DW_mult_tc_2 is

   component AOI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component MUXB2DL
      port( A0, A1, SL : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal n42, n50, n58, n66, n73, n80, n84, n89, n94, n99, n104, n156, n157, 
      n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, 
      n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, 
      n182, n183, n184, n185, n186, n202, n203, n204, n205, n206, n207, n208, 
      n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, 
      n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, 
      n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, 
      n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, 
      n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, 
      n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, 
      n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
      n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, 
      n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, 
      n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, 
      n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, 
      n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, 
      n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, 
      n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, 
      n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, 
      n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, 
      n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, 
      n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, 
      n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, 
      n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, 
      n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, 
      n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, 
      n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, 
      n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, 
      n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, 
      n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, 
      n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
      n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, 
      n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, 
      n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, 
      n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
      n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, 
      n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, 
      n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, 
      n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, 
      n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, 
      n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, 
      n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, 
      n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, 
      n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, 
      n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, 
      n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, 
      n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, 
      n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, 
      n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, 
      n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, 
      n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, 
      n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, 
      n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, 
      n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, 
      n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, 
      n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, 
      n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, 
      n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, 
      n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, 
      n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, 
      n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, 
      n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, 
      n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, 
      n917, n918, n919, n920, n921, n922, n923, n939, n940, n941, n942, n943, 
      n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n955, n956, 
      n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, 
      n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, 
      n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, 
      n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, 
      n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, 
      n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, 
      n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, 
      n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, 
      n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, 
      n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, 
      n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, 
      n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, 
      n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, 
      n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, 
      n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, 
      n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, 
      n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, 
      n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, 
      n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, 
      n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, 
      n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, 
      n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, 
      n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, 
      n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, 
      n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, 
      n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, 
      n1224, n1225, n1226, n1375, n1376, n1377, n1378, n1379, n1380, n1381, 
      n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, 
      n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, 
      n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, 
      n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, 
      n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, 
      n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, 
      n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451 : 
      std_logic;

begin
   
   U125 : ADFULD1 port map( A => n203, B => n232, CI => n157, CO => n156, S => 
                           product(30));
   U126 : ADFULD1 port map( A => n233, B => n260, CI => n158, CO => n157, S => 
                           product(29));
   U127 : ADFULD1 port map( A => n261, B => n288, CI => n159, CO => n158, S => 
                           product(28));
   U128 : ADFULD1 port map( A => n289, B => n314, CI => n160, CO => n159, S => 
                           product(27));
   U129 : ADFULD1 port map( A => n315, B => n340, CI => n161, CO => n160, S => 
                           product(26));
   U130 : ADFULD1 port map( A => n341, B => n364, CI => n162, CO => n161, S => 
                           product(25));
   U131 : ADFULD1 port map( A => n365, B => n388, CI => n163, CO => n162, S => 
                           product(24));
   U132 : ADFULD1 port map( A => n389, B => n410, CI => n164, CO => n163, S => 
                           product(23));
   U133 : ADFULD1 port map( A => n411, B => n432, CI => n165, CO => n164, S => 
                           product(22));
   U134 : ADFULD1 port map( A => n433, B => n452, CI => n166, CO => n165, S => 
                           product(21));
   U135 : ADFULD1 port map( A => n453, B => n472, CI => n167, CO => n166, S => 
                           product(20));
   U136 : ADFULD1 port map( A => n473, B => n490, CI => n168, CO => n167, S => 
                           product(19));
   U137 : ADFULD1 port map( A => n491, B => n508, CI => n169, CO => n168, S => 
                           product(18));
   U138 : ADFULD1 port map( A => n509, B => n524, CI => n170, CO => n169, S => 
                           product(17));
   U139 : ADFULD1 port map( A => n525, B => n540, CI => n171, CO => n170, S => 
                           product(16));
   U140 : ADFULD1 port map( A => n541, B => n554, CI => n172, CO => n171, S => 
                           product(15));
   U141 : ADFULD1 port map( A => n555, B => n568, CI => n173, CO => n172, S => 
                           product(14));
   U142 : ADFULD1 port map( A => n569, B => n580, CI => n174, CO => n173, S => 
                           product(13));
   U143 : ADFULD1 port map( A => n581, B => n592, CI => n175, CO => n174, S => 
                           product(12));
   U144 : ADFULD1 port map( A => n593, B => n602, CI => n176, CO => n175, S => 
                           product(11));
   U145 : ADFULD1 port map( A => n603, B => n612, CI => n177, CO => n176, S => 
                           product(10));
   U146 : ADFULD1 port map( A => n613, B => n620, CI => n178, CO => n177, S => 
                           product(9));
   U147 : ADFULD1 port map( A => n621, B => n628, CI => n179, CO => n178, S => 
                           product(8));
   U148 : ADFULD1 port map( A => n629, B => n634, CI => n180, CO => n179, S => 
                           product(7));
   U149 : ADFULD1 port map( A => n635, B => n640, CI => n181, CO => n180, S => 
                           product(6));
   U150 : ADFULD1 port map( A => n641, B => n644, CI => n182, CO => n181, S => 
                           product(5));
   U151 : ADFULD1 port map( A => n645, B => n648, CI => n183, CO => n182, S => 
                           product(4));
   U152 : ADFULD1 port map( A => n649, B => n1193, CI => n184, CO => n183, S =>
                           product(3));
   U153 : ADFULD1 port map( A => n651, B => n1194, CI => n185, CO => n184, S =>
                           product(2));
   U154 : ADHALFDL port map( A => n186, B => n1225, CO => n185, S => product(1)
                           );
   U155 : ADHALFDL port map( A => n1226, B => a(1), CO => n186, S => product(0)
                           );
   U171 : ADFULD1 port map( A => n234, B => n207, CI => n205, CO => n202, S => 
                           n203);
   U172 : ADFULD1 port map( A => n209, B => n211, CI => n236, CO => n204, S => 
                           n205);
   U173 : ADFULD1 port map( A => n240, B => n213, CI => n238, CO => n206, S => 
                           n207);
   U174 : ADFULD1 port map( A => n217, B => n242, CI => n215, CO => n208, S => 
                           n209);
   U175 : ADFULD1 port map( A => n244, B => n246, CI => n219, CO => n210, S => 
                           n211);
   U176 : ADFULD1 port map( A => n225, B => n223, CI => n248, CO => n212, S => 
                           n213);
   U177 : ADFULD1 port map( A => n221, B => n229, CI => n227, CO => n214, S => 
                           n215);
   U178 : ADFULD1 port map( A => n256, B => n252, CI => n254, CO => n216, S => 
                           n217);
   U179 : ADFULD1 port map( A => n258, B => n1088, CI => n250, CO => n218, S =>
                           n219);
   U180 : ADFULD1 port map( A => n1046, B => n1112, CI => n1066, CO => n220, S 
                           => n221);
   U181 : ADFULD1 port map( A => n986, B => n976, CI => n998, CO => n222, S => 
                           n223);
   U182 : ADFULD1 port map( A => n962, B => n1138, CI => n968, CO => n224, S =>
                           n225);
   U183 : ADFULD1 port map( A => n1166, B => n1012, CI => n231, CO => n226, S 
                           => n227);
   U184 : ADFULD1 port map( A => n1028, B => n956, CI => n958, CO => n228, S =>
                           n229);
   U185 : ADHALFDL port map( A => n1196, B => n939, CO => n230, S => n231);
   U186 : ADFULD1 port map( A => n262, B => n237, CI => n235, CO => n232, S => 
                           n233);
   U187 : ADFULD1 port map( A => n239, B => n266, CI => n264, CO => n234, S => 
                           n235);
   U188 : ADFULD1 port map( A => n268, B => n243, CI => n241, CO => n236, S => 
                           n237);
   U189 : ADFULD1 port map( A => n270, B => n247, CI => n245, CO => n238, S => 
                           n239);
   U190 : ADFULD1 port map( A => n274, B => n249, CI => n272, CO => n240, S => 
                           n241);
   U191 : ADFULD1 port map( A => n253, B => n255, CI => n257, CO => n242, S => 
                           n243);
   U192 : ADFULD1 port map( A => n280, B => n276, CI => n251, CO => n244, S => 
                           n245);
   U193 : ADFULD1 port map( A => n278, B => n284, CI => n282, CO => n246, S => 
                           n247);
   U194 : ADFULD1 port map( A => n1047, B => n1013, CI => n259, CO => n248, S 
                           => n249);
   U195 : ADFULD1 port map( A => n977, B => n1067, CI => n999, CO => n250, S =>
                           n251);
   U196 : ADFULD1 port map( A => n959, B => n969, CI => n963, CO => n252, S => 
                           n253);
   U197 : ADFULD1 port map( A => n1113, B => n987, CI => n1089, CO => n254, S 
                           => n255);
   U198 : ADFULD1 port map( A => n1167, B => n1029, CI => n1139, CO => n256, S 
                           => n257);
   U199 : ADHALFDL port map( A => n286, B => n1197, CO => n258, S => n259);
   U200 : ADFULD1 port map( A => n290, B => n265, CI => n263, CO => n260, S => 
                           n261);
   U201 : ADFULD1 port map( A => n267, B => n294, CI => n292, CO => n262, S => 
                           n263);
   U202 : ADFULD1 port map( A => n296, B => n271, CI => n269, CO => n264, S => 
                           n265);
   U203 : ADFULD1 port map( A => n275, B => n298, CI => n273, CO => n266, S => 
                           n267);
   U204 : ADFULD1 port map( A => n302, B => n281, CI => n300, CO => n268, S => 
                           n269);
   U205 : ADFULD1 port map( A => n283, B => n277, CI => n279, CO => n270, S => 
                           n271);
   U206 : ADFULD1 port map( A => n310, B => n308, CI => n285, CO => n272, S => 
                           n273);
   U207 : ADFULD1 port map( A => n304, B => n312, CI => n306, CO => n274, S => 
                           n275);
   U208 : ADFULD1 port map( A => n1014, B => n1068, CI => n1048, CO => n276, S 
                           => n277);
   U209 : ADFULD1 port map( A => n978, B => n1090, CI => n988, CO => n278, S =>
                           n279);
   U210 : ADFULD1 port map( A => n964, B => n1114, CI => n970, CO => n280, S =>
                           n281);
   U211 : ADFULD1 port map( A => n1140, B => n1000, CI => n287, CO => n282, S 
                           => n283);
   U212 : ADFULD1 port map( A => n1030, B => n960, CI => n1168, CO => n284, S 
                           => n285);
   U213 : ADHALFDL port map( A => n1198, B => n940, CO => n286, S => n287);
   U214 : ADFULD1 port map( A => n316, B => n293, CI => n291, CO => n288, S => 
                           n289);
   U215 : ADFULD1 port map( A => n318, B => n297, CI => n295, CO => n290, S => 
                           n291);
   U216 : ADFULD1 port map( A => n299, B => n322, CI => n320, CO => n292, S => 
                           n293);
   U217 : ADFULD1 port map( A => n324, B => n303, CI => n301, CO => n294, S => 
                           n295);
   U218 : ADFULD1 port map( A => n307, B => n309, CI => n326, CO => n296, S => 
                           n297);
   U219 : ADFULD1 port map( A => n305, B => n328, CI => n311, CO => n298, S => 
                           n299);
   U220 : ADFULD1 port map( A => n332, B => n330, CI => n334, CO => n300, S => 
                           n301);
   U221 : ADFULD1 port map( A => n313, B => n1091, CI => n336, CO => n302, S =>
                           n303);
   U222 : ADFULD1 port map( A => n1015, B => n1115, CI => n1069, CO => n304, S 
                           => n305);
   U223 : ADFULD1 port map( A => n1141, B => n1001, CI => n989, CO => n306, S 
                           => n307);
   U224 : ADFULD1 port map( A => n979, B => n1049, CI => n1169, CO => n308, S 
                           => n309);
   U225 : ADFULD1 port map( A => n965, B => n1031, CI => n971, CO => n310, S =>
                           n311);
   U226 : ADHALFDL port map( A => n338, B => n1199, CO => n312, S => n313);
   U227 : ADFULD1 port map( A => n342, B => n319, CI => n317, CO => n314, S => 
                           n315);
   U228 : ADFULD1 port map( A => n344, B => n346, CI => n321, CO => n316, S => 
                           n317);
   U229 : ADFULD1 port map( A => n325, B => n327, CI => n323, CO => n318, S => 
                           n319);
   U230 : ADFULD1 port map( A => n350, B => n352, CI => n348, CO => n320, S => 
                           n321);
   U231 : ADFULD1 port map( A => n333, B => n335, CI => n329, CO => n322, S => 
                           n323);
   U232 : ADFULD1 port map( A => n337, B => n358, CI => n331, CO => n324, S => 
                           n325);
   U233 : ADFULD1 port map( A => n354, B => n360, CI => n356, CO => n326, S => 
                           n327);
   U234 : ADFULD1 port map( A => n1092, B => n1116, CI => n362, CO => n328, S 
                           => n329);
   U235 : ADFULD1 port map( A => n1016, B => n1142, CI => n1070, CO => n330, S 
                           => n331);
   U236 : ADFULD1 port map( A => n990, B => n1170, CI => n1002, CO => n332, S 
                           => n333);
   U237 : ADFULD1 port map( A => n980, B => n1032, CI => n339, CO => n334, S =>
                           n335);
   U238 : ADFULD1 port map( A => n1050, B => n966, CI => n972, CO => n336, S =>
                           n337);
   U239 : ADHALFDL port map( A => n1200, B => n941, CO => n338, S => n339);
   U240 : ADFULD1 port map( A => n366, B => n345, CI => n343, CO => n340, S => 
                           n341);
   U241 : ADFULD1 port map( A => n347, B => n370, CI => n368, CO => n342, S => 
                           n343);
   U242 : ADFULD1 port map( A => n351, B => n372, CI => n349, CO => n344, S => 
                           n345);
   U243 : ADFULD1 port map( A => n374, B => n376, CI => n353, CO => n346, S => 
                           n347);
   U244 : ADFULD1 port map( A => n361, B => n357, CI => n359, CO => n348, S => 
                           n349);
   U245 : ADFULD1 port map( A => n378, B => n380, CI => n355, CO => n350, S => 
                           n351);
   U246 : ADFULD1 port map( A => n384, B => n363, CI => n382, CO => n352, S => 
                           n353);
   U247 : ADFULD1 port map( A => n1033, B => n1093, CI => n1071, CO => n354, S 
                           => n355);
   U248 : ADFULD1 port map( A => n991, B => n1117, CI => n1017, CO => n356, S 
                           => n357);
   U249 : ADFULD1 port map( A => n973, B => n1003, CI => n981, CO => n358, S =>
                           n359);
   U250 : ADFULD1 port map( A => n1171, B => n1051, CI => n1143, CO => n360, S 
                           => n361);
   U251 : ADHALFDL port map( A => n386, B => n1201, CO => n362, S => n363);
   U252 : ADFULD1 port map( A => n390, B => n369, CI => n367, CO => n364, S => 
                           n365);
   U253 : ADFULD1 port map( A => n371, B => n394, CI => n392, CO => n366, S => 
                           n367);
   U254 : ADFULD1 port map( A => n375, B => n396, CI => n373, CO => n368, S => 
                           n369);
   U255 : ADFULD1 port map( A => n398, B => n400, CI => n377, CO => n370, S => 
                           n371);
   U256 : ADFULD1 port map( A => n383, B => n379, CI => n381, CO => n372, S => 
                           n373);
   U257 : ADFULD1 port map( A => n402, B => n404, CI => n385, CO => n374, S => 
                           n375);
   U258 : ADFULD1 port map( A => n408, B => n1072, CI => n406, CO => n376, S =>
                           n377);
   U259 : ADFULD1 port map( A => n1004, B => n1094, CI => n1034, CO => n378, S 
                           => n379);
   U260 : ADFULD1 port map( A => n992, B => n1144, CI => n1118, CO => n380, S 
                           => n381);
   U261 : ADFULD1 port map( A => n982, B => n1018, CI => n387, CO => n382, S =>
                           n383);
   U262 : ADFULD1 port map( A => n1052, B => n974, CI => n1172, CO => n384, S 
                           => n385);
   U263 : ADHALFDL port map( A => n1202, B => n942, CO => n386, S => n387);
   U264 : ADFULD1 port map( A => n412, B => n393, CI => n391, CO => n388, S => 
                           n389);
   U265 : ADFULD1 port map( A => n395, B => n397, CI => n414, CO => n390, S => 
                           n391);
   U266 : ADFULD1 port map( A => n399, B => n418, CI => n416, CO => n392, S => 
                           n393);
   U267 : ADFULD1 port map( A => n401, B => n407, CI => n420, CO => n394, S => 
                           n395);
   U268 : ADFULD1 port map( A => n403, B => n424, CI => n405, CO => n396, S => 
                           n397);
   U269 : ADFULD1 port map( A => n426, B => n428, CI => n422, CO => n398, S => 
                           n399);
   U270 : ADFULD1 port map( A => n1073, B => n1095, CI => n409, CO => n400, S 
                           => n401);
   U271 : ADFULD1 port map( A => n1005, B => n1119, CI => n1019, CO => n402, S 
                           => n403);
   U272 : ADFULD1 port map( A => n1173, B => n1035, CI => n1145, CO => n404, S 
                           => n405);
   U273 : ADFULD1 port map( A => n983, B => n1053, CI => n993, CO => n406, S =>
                           n407);
   U274 : ADHALFDL port map( A => n430, B => n1203, CO => n408, S => n409);
   U275 : ADFULD1 port map( A => n434, B => n415, CI => n413, CO => n410, S => 
                           n411);
   U276 : ADFULD1 port map( A => n417, B => n419, CI => n436, CO => n412, S => 
                           n413);
   U277 : ADFULD1 port map( A => n421, B => n440, CI => n438, CO => n414, S => 
                           n415);
   U278 : ADFULD1 port map( A => n427, B => n425, CI => n442, CO => n416, S => 
                           n417);
   U279 : ADFULD1 port map( A => n429, B => n444, CI => n423, CO => n418, S => 
                           n419);
   U280 : ADFULD1 port map( A => n448, B => n450, CI => n446, CO => n420, S => 
                           n421);
   U281 : ADFULD1 port map( A => n1074, B => n1120, CI => n1096, CO => n422, S 
                           => n423);
   U282 : ADFULD1 port map( A => n1006, B => n1146, CI => n1020, CO => n424, S 
                           => n425);
   U283 : ADFULD1 port map( A => n1174, B => n1036, CI => n431, CO => n426, S 
                           => n427);
   U284 : ADFULD1 port map( A => n1054, B => n984, CI => n994, CO => n428, S =>
                           n429);
   U285 : ADHALFDL port map( A => n1204, B => n943, CO => n430, S => n431);
   U286 : ADFULD1 port map( A => n454, B => n437, CI => n435, CO => n432, S => 
                           n433);
   U287 : ADFULD1 port map( A => n439, B => n441, CI => n456, CO => n434, S => 
                           n435);
   U288 : ADFULD1 port map( A => n443, B => n460, CI => n458, CO => n436, S => 
                           n437);
   U289 : ADFULD1 port map( A => n449, B => n445, CI => n447, CO => n438, S => 
                           n439);
   U290 : ADFULD1 port map( A => n464, B => n466, CI => n462, CO => n440, S => 
                           n441);
   U291 : ADFULD1 port map( A => n451, B => n1037, CI => n468, CO => n442, S =>
                           n443);
   U292 : ADFULD1 port map( A => n995, B => n1075, CI => n1007, CO => n444, S 
                           => n445);
   U293 : ADFULD1 port map( A => n1121, B => n1021, CI => n1097, CO => n446, S 
                           => n447);
   U294 : ADFULD1 port map( A => n1175, B => n1055, CI => n1147, CO => n448, S 
                           => n449);
   U295 : ADHALFDL port map( A => n470, B => n1205, CO => n450, S => n451);
   U296 : ADFULD1 port map( A => n474, B => n457, CI => n455, CO => n452, S => 
                           n453);
   U297 : ADFULD1 port map( A => n459, B => n461, CI => n476, CO => n454, S => 
                           n455);
   U298 : ADFULD1 port map( A => n480, B => n463, CI => n478, CO => n456, S => 
                           n457);
   U299 : ADFULD1 port map( A => n465, B => n469, CI => n467, CO => n458, S => 
                           n459);
   U300 : ADFULD1 port map( A => n482, B => n486, CI => n484, CO => n460, S => 
                           n461);
   U301 : ADFULD1 port map( A => n1098, B => n1122, CI => n488, CO => n462, S 
                           => n463);
   U302 : ADFULD1 port map( A => n1022, B => n1148, CI => n1056, CO => n464, S 
                           => n465);
   U303 : ADFULD1 port map( A => n1008, B => n1038, CI => n471, CO => n466, S 
                           => n467);
   U304 : ADFULD1 port map( A => n1076, B => n996, CI => n1176, CO => n468, S 
                           => n469);
   U305 : ADHALFDL port map( A => n1206, B => n944, CO => n470, S => n471);
   U306 : ADFULD1 port map( A => n492, B => n477, CI => n475, CO => n472, S => 
                           n473);
   U307 : ADFULD1 port map( A => n479, B => n481, CI => n494, CO => n474, S => 
                           n475);
   U308 : ADFULD1 port map( A => n498, B => n487, CI => n496, CO => n476, S => 
                           n477);
   U309 : ADFULD1 port map( A => n483, B => n500, CI => n485, CO => n478, S => 
                           n479);
   U310 : ADFULD1 port map( A => n504, B => n489, CI => n502, CO => n480, S => 
                           n481);
   U311 : ADFULD1 port map( A => n1057, B => n1149, CI => n1123, CO => n482, S 
                           => n483);
   U312 : ADFULD1 port map( A => n1177, B => n1099, CI => n1039, CO => n484, S 
                           => n485);
   U313 : ADFULD1 port map( A => n1009, B => n1077, CI => n1023, CO => n486, S 
                           => n487);
   U314 : ADHALFDL port map( A => n506, B => n1207, CO => n488, S => n489);
   U315 : ADFULD1 port map( A => n510, B => n495, CI => n493, CO => n490, S => 
                           n491);
   U316 : ADFULD1 port map( A => n497, B => n499, CI => n512, CO => n492, S => 
                           n493);
   U317 : ADFULD1 port map( A => n516, B => n503, CI => n514, CO => n494, S => 
                           n495);
   U318 : ADFULD1 port map( A => n505, B => n518, CI => n501, CO => n496, S => 
                           n497);
   U319 : ADFULD1 port map( A => n522, B => n1124, CI => n520, CO => n498, S =>
                           n499);
   U320 : ADFULD1 port map( A => n1040, B => n1150, CI => n1058, CO => n500, S 
                           => n501);
   U321 : ADFULD1 port map( A => n1178, B => n1100, CI => n507, CO => n502, S 
                           => n503);
   U322 : ADFULD1 port map( A => n1078, B => n1010, CI => n1024, CO => n504, S 
                           => n505);
   U323 : ADHALFDL port map( A => n1208, B => n945, CO => n506, S => n507);
   U324 : ADFULD1 port map( A => n526, B => n513, CI => n511, CO => n508, S => 
                           n509);
   U325 : ADFULD1 port map( A => n528, B => n530, CI => n515, CO => n510, S => 
                           n511);
   U326 : ADFULD1 port map( A => n521, B => n519, CI => n517, CO => n512, S => 
                           n513);
   U327 : ADFULD1 port map( A => n534, B => n536, CI => n532, CO => n514, S => 
                           n515);
   U328 : ADFULD1 port map( A => n1101, B => n1125, CI => n523, CO => n516, S 
                           => n517);
   U329 : ADFULD1 port map( A => n1025, B => n1041, CI => n1059, CO => n518, S 
                           => n519);
   U330 : ADFULD1 port map( A => n1179, B => n1079, CI => n1151, CO => n520, S 
                           => n521);
   U331 : ADHALFDL port map( A => n538, B => n1209, CO => n522, S => n523);
   U332 : ADFULD1 port map( A => n542, B => n529, CI => n527, CO => n524, S => 
                           n525);
   U333 : ADFULD1 port map( A => n544, B => n546, CI => n531, CO => n526, S => 
                           n527);
   U334 : ADFULD1 port map( A => n533, B => n537, CI => n535, CO => n528, S => 
                           n529);
   U335 : ADFULD1 port map( A => n550, B => n552, CI => n548, CO => n530, S => 
                           n531);
   U336 : ADFULD1 port map( A => n1080, B => n1152, CI => n1126, CO => n532, S 
                           => n533);
   U337 : ADFULD1 port map( A => n1042, B => n1060, CI => n539, CO => n534, S 
                           => n535);
   U338 : ADFULD1 port map( A => n1102, B => n1026, CI => n1180, CO => n536, S 
                           => n537);
   U339 : ADHALFDL port map( A => n1210, B => n946, CO => n538, S => n539);
   U340 : ADFULD1 port map( A => n556, B => n545, CI => n543, CO => n540, S => 
                           n541);
   U341 : ADFULD1 port map( A => n547, B => n551, CI => n558, CO => n542, S => 
                           n543);
   U342 : ADFULD1 port map( A => n560, B => n562, CI => n549, CO => n544, S => 
                           n545);
   U343 : ADFULD1 port map( A => n553, B => n1153, CI => n564, CO => n546, S =>
                           n547);
   U344 : ADFULD1 port map( A => n1181, B => n1081, CI => n1127, CO => n548, S 
                           => n549);
   U345 : ADFULD1 port map( A => n1043, B => n1103, CI => n1061, CO => n550, S 
                           => n551);
   U346 : ADHALFDL port map( A => n566, B => n1211, CO => n552, S => n553);
   U347 : ADFULD1 port map( A => n570, B => n559, CI => n557, CO => n554, S => 
                           n555);
   U348 : ADFULD1 port map( A => n561, B => n563, CI => n572, CO => n556, S => 
                           n557);
   U349 : ADFULD1 port map( A => n574, B => n576, CI => n565, CO => n558, S => 
                           n559);
   U350 : ADFULD1 port map( A => n1062, B => n1128, CI => n578, CO => n560, S 
                           => n561);
   U351 : ADFULD1 port map( A => n1154, B => n1082, CI => n567, CO => n562, S 
                           => n563);
   U352 : ADFULD1 port map( A => n1104, B => n1044, CI => n1182, CO => n564, S 
                           => n565);
   U353 : ADHALFDL port map( A => n1212, B => n947, CO => n566, S => n567);
   U354 : ADFULD1 port map( A => n582, B => n573, CI => n571, CO => n568, S => 
                           n569);
   U355 : ADFULD1 port map( A => n577, B => n575, CI => n584, CO => n570, S => 
                           n571);
   U356 : ADFULD1 port map( A => n588, B => n579, CI => n586, CO => n572, S => 
                           n573);
   U357 : ADFULD1 port map( A => n1063, B => n1129, CI => n1083, CO => n574, S 
                           => n575);
   U358 : ADFULD1 port map( A => n1183, B => n1105, CI => n1155, CO => n576, S 
                           => n577);
   U359 : ADHALFDL port map( A => n590, B => n1213, CO => n578, S => n579);
   U360 : ADFULD1 port map( A => n585, B => n594, CI => n583, CO => n580, S => 
                           n581);
   U361 : ADFULD1 port map( A => n587, B => n589, CI => n596, CO => n582, S => 
                           n583);
   U362 : ADFULD1 port map( A => n600, B => n1106, CI => n598, CO => n584, S =>
                           n585);
   U363 : ADFULD1 port map( A => n1084, B => n1156, CI => n591, CO => n586, S 
                           => n587);
   U364 : ADFULD1 port map( A => n1130, B => n1064, CI => n1184, CO => n588, S 
                           => n589);
   U365 : ADHALFDL port map( A => n1214, B => n948, CO => n590, S => n591);
   U366 : ADFULD1 port map( A => n604, B => n597, CI => n595, CO => n592, S => 
                           n593);
   U367 : ADFULD1 port map( A => n606, B => n608, CI => n599, CO => n594, S => 
                           n595);
   U368 : ADFULD1 port map( A => n1107, B => n1157, CI => n601, CO => n596, S 
                           => n597);
   U369 : ADFULD1 port map( A => n1085, B => n1131, CI => n1185, CO => n598, S 
                           => n599);
   U370 : ADHALFDL port map( A => n610, B => n1215, CO => n600, S => n601);
   U371 : ADFULD1 port map( A => n614, B => n607, CI => n605, CO => n602, S => 
                           n603);
   U372 : ADFULD1 port map( A => n616, B => n618, CI => n609, CO => n604, S => 
                           n605);
   U373 : ADFULD1 port map( A => n1108, B => n1158, CI => n611, CO => n606, S 
                           => n607);
   U374 : ADFULD1 port map( A => n1132, B => n1086, CI => n1186, CO => n608, S 
                           => n609);
   U375 : ADHALFDL port map( A => n1216, B => n949, CO => n610, S => n611);
   U376 : ADFULD1 port map( A => n617, B => n622, CI => n615, CO => n612, S => 
                           n613);
   U377 : ADFULD1 port map( A => n619, B => n1187, CI => n624, CO => n614, S =>
                           n615);
   U378 : ADFULD1 port map( A => n1109, B => n1133, CI => n1159, CO => n616, S 
                           => n617);
   U379 : ADHALFDL port map( A => n626, B => n1217, CO => n618, S => n619);
   U380 : ADFULD1 port map( A => n625, B => n630, CI => n623, CO => n620, S => 
                           n621);
   U381 : ADFULD1 port map( A => n627, B => n1160, CI => n632, CO => n622, S =>
                           n623);
   U382 : ADFULD1 port map( A => n1188, B => n1110, CI => n1134, CO => n624, S 
                           => n625);
   U383 : ADHALFDL port map( A => n1218, B => n950, CO => n626, S => n627);
   U384 : ADFULD1 port map( A => n636, B => n633, CI => n631, CO => n628, S => 
                           n629);
   U385 : ADFULD1 port map( A => n1135, B => n1189, CI => n1161, CO => n630, S 
                           => n631);
   U386 : ADHALFDL port map( A => n638, B => n1219, CO => n632, S => n633);
   U387 : ADFULD1 port map( A => n642, B => n639, CI => n637, CO => n634, S => 
                           n635);
   U388 : ADFULD1 port map( A => n1190, B => n1136, CI => n1162, CO => n636, S 
                           => n637);
   U389 : ADHALFDL port map( A => n1220, B => n951, CO => n638, S => n639);
   U390 : ADFULD1 port map( A => n1163, B => n1191, CI => n643, CO => n640, S 
                           => n641);
   U391 : ADHALFDL port map( A => n646, B => n1221, CO => n642, S => n643);
   U392 : ADFULD1 port map( A => n1192, B => n1164, CI => n647, CO => n644, S 
                           => n645);
   U393 : ADHALFDL port map( A => n1222, B => n952, CO => n646, S => n647);
   U394 : ADHALFDL port map( A => n650, B => n1223, CO => n648, S => n649);
   U395 : ADHALFDL port map( A => n1224, B => n953, CO => n650, S => n651);
   U397 : MUXB2DL port map( A0 => n104, A1 => n1420, SL => n652, Z => n955);
   U399 : MUXB2DL port map( A0 => n104, A1 => n1420, SL => n653, Z => n956);
   U402 : MUXB2DL port map( A0 => n99, A1 => n1419, SL => n654, Z => n957);
   U404 : MUXB2DL port map( A0 => n99, A1 => n1419, SL => n655, Z => n958);
   U406 : MUXB2DL port map( A0 => n99, A1 => n1419, SL => n656, Z => n959);
   U408 : MUXB2DL port map( A0 => n99, A1 => n1419, SL => n657, Z => n960);
   U411 : MUXB2DL port map( A0 => n94, A1 => n1416, SL => n658, Z => n961);
   U413 : MUXB2DL port map( A0 => n94, A1 => n1416, SL => n659, Z => n962);
   U415 : MUXB2DL port map( A0 => n94, A1 => n1416, SL => n660, Z => n963);
   U417 : MUXB2DL port map( A0 => n94, A1 => n1416, SL => n661, Z => n964);
   U419 : MUXB2DL port map( A0 => n94, A1 => n1416, SL => n662, Z => n965);
   U421 : MUXB2DL port map( A0 => n94, A1 => n1416, SL => n663, Z => n966);
   U424 : MUXB2DL port map( A0 => n89, A1 => n1414, SL => n664, Z => n967);
   U426 : MUXB2DL port map( A0 => n89, A1 => n1414, SL => n665, Z => n968);
   U428 : MUXB2DL port map( A0 => n89, A1 => n1414, SL => n666, Z => n969);
   U430 : MUXB2DL port map( A0 => n89, A1 => n1414, SL => n667, Z => n970);
   U432 : MUXB2DL port map( A0 => n89, A1 => n1414, SL => n668, Z => n971);
   U434 : MUXB2DL port map( A0 => n89, A1 => n1414, SL => n669, Z => n972);
   U436 : MUXB2DL port map( A0 => n89, A1 => n1414, SL => n670, Z => n973);
   U438 : MUXB2DL port map( A0 => n89, A1 => n1414, SL => n671, Z => n974);
   U441 : MUXB2DL port map( A0 => n84, A1 => n1412, SL => n672, Z => n975);
   U443 : MUXB2DL port map( A0 => n84, A1 => n1412, SL => n673, Z => n976);
   U445 : MUXB2DL port map( A0 => n84, A1 => n1412, SL => n674, Z => n977);
   U447 : MUXB2DL port map( A0 => n84, A1 => n1412, SL => n675, Z => n978);
   U449 : MUXB2DL port map( A0 => n84, A1 => n1412, SL => n676, Z => n979);
   U451 : MUXB2DL port map( A0 => n84, A1 => n1412, SL => n677, Z => n980);
   U453 : MUXB2DL port map( A0 => n84, A1 => n1412, SL => n678, Z => n981);
   U455 : MUXB2DL port map( A0 => n84, A1 => n1412, SL => n679, Z => n982);
   U457 : MUXB2DL port map( A0 => n84, A1 => n1412, SL => n680, Z => n983);
   U459 : MUXB2DL port map( A0 => n84, A1 => n1412, SL => n681, Z => n984);
   U462 : MUXB2DL port map( A0 => n80, A1 => n1410, SL => n682, Z => n985);
   U464 : MUXB2DL port map( A0 => n80, A1 => n1410, SL => n683, Z => n986);
   U466 : MUXB2DL port map( A0 => n80, A1 => n1410, SL => n684, Z => n987);
   U468 : MUXB2DL port map( A0 => n80, A1 => n1410, SL => n685, Z => n988);
   U470 : MUXB2DL port map( A0 => n80, A1 => n1410, SL => n686, Z => n989);
   U472 : MUXB2DL port map( A0 => n80, A1 => n1410, SL => n687, Z => n990);
   U474 : MUXB2DL port map( A0 => n80, A1 => n1410, SL => n688, Z => n991);
   U476 : MUXB2DL port map( A0 => n80, A1 => n1410, SL => n689, Z => n992);
   U478 : MUXB2DL port map( A0 => n80, A1 => n1410, SL => n690, Z => n993);
   U480 : MUXB2DL port map( A0 => n80, A1 => n1410, SL => n691, Z => n994);
   U482 : MUXB2DL port map( A0 => n80, A1 => n1410, SL => n692, Z => n995);
   U484 : MUXB2DL port map( A0 => n80, A1 => n1410, SL => n693, Z => n996);
   U487 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n694, Z => n997);
   U489 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n695, Z => n998);
   U491 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n696, Z => n999);
   U493 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n697, Z => n1000);
   U495 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n698, Z => n1001);
   U497 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n699, Z => n1002);
   U499 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n700, Z => n1003);
   U501 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n701, Z => n1004);
   U503 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n702, Z => n1005);
   U505 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n703, Z => n1006);
   U507 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n704, Z => n1007);
   U509 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n705, Z => n1008);
   U511 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n706, Z => n1009);
   U513 : MUXB2DL port map( A0 => n73, A1 => n1408, SL => n707, Z => n1010);
   U516 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n708, Z => n1011);
   U518 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n709, Z => n1012);
   U520 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n710, Z => n1013);
   U522 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n711, Z => n1014);
   U524 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n712, Z => n1015);
   U526 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n713, Z => n1016);
   U528 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n714, Z => n1017);
   U530 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n715, Z => n1018);
   U532 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n716, Z => n1019);
   U534 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n717, Z => n1020);
   U536 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n718, Z => n1021);
   U538 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n719, Z => n1022);
   U540 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n720, Z => n1023);
   U542 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n721, Z => n1024);
   U544 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n722, Z => n1025);
   U546 : MUXB2DL port map( A0 => n66, A1 => n1406, SL => n723, Z => n1026);
   U549 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n724, Z => n1027);
   U551 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n725, Z => n1028);
   U553 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n726, Z => n1029);
   U555 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n727, Z => n1030);
   U557 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n728, Z => n1031);
   U559 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n729, Z => n1032);
   U561 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n730, Z => n1033);
   U563 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n731, Z => n1034);
   U565 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n732, Z => n1035);
   U567 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n733, Z => n1036);
   U569 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n734, Z => n1037);
   U571 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n735, Z => n1038);
   U573 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n736, Z => n1039);
   U575 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n737, Z => n1040);
   U577 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n738, Z => n1041);
   U579 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n739, Z => n1042);
   U581 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n740, Z => n1043);
   U583 : MUXB2DL port map( A0 => n58, A1 => n1404, SL => n741, Z => n1044);
   U586 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n742, Z => n1045);
   U588 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n743, Z => n1046);
   U590 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n744, Z => n1047);
   U592 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n745, Z => n1048);
   U594 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n746, Z => n1049);
   U596 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n747, Z => n1050);
   U598 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n748, Z => n1051);
   U600 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n749, Z => n1052);
   U602 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n750, Z => n1053);
   U604 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n751, Z => n1054);
   U606 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n752, Z => n1055);
   U608 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n753, Z => n1056);
   U610 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n754, Z => n1057);
   U612 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n755, Z => n1058);
   U614 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n756, Z => n1059);
   U616 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n757, Z => n1060);
   U618 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n758, Z => n1061);
   U620 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n759, Z => n1062);
   U622 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n760, Z => n1063);
   U624 : MUXB2DL port map( A0 => n50, A1 => n1402, SL => n761, Z => n1064);
   U627 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n762, Z => n1065);
   U629 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n763, Z => n1066);
   U631 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n764, Z => n1067);
   U633 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n765, Z => n1068);
   U635 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n766, Z => n1069);
   U637 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n767, Z => n1070);
   U639 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n768, Z => n1071);
   U641 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n769, Z => n1072);
   U643 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n770, Z => n1073);
   U645 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n771, Z => n1074);
   U647 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n772, Z => n1075);
   U649 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n773, Z => n1076);
   U651 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n774, Z => n1077);
   U653 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n775, Z => n1078);
   U655 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n776, Z => n1079);
   U657 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n777, Z => n1080);
   U659 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n778, Z => n1081);
   U661 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n779, Z => n1082);
   U663 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n780, Z => n1083);
   U665 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n781, Z => n1084);
   U667 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n782, Z => n1085);
   U669 : MUXB2DL port map( A0 => n42, A1 => n1400, SL => n783, Z => n1086);
   U672 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n784, Z => n1087);
   U674 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n785, Z => n1088);
   U676 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n786, Z => n1089);
   U678 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n787, Z => n1090);
   U680 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n788, Z => n1091);
   U682 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n789, Z => n1092);
   U684 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n790, Z => n1093);
   U686 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n791, Z => n1094);
   U688 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n792, Z => n1095);
   U690 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n793, Z => n1096);
   U692 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n794, Z => n1097);
   U694 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n795, Z => n1098);
   U696 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n796, Z => n1099);
   U698 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n797, Z => n1100);
   U700 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n798, Z => n1101);
   U702 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n799, Z => n1102);
   U704 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n800, Z => n1103);
   U706 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n801, Z => n1104);
   U708 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n802, Z => n1105);
   U710 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n803, Z => n1106);
   U712 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n804, Z => n1107);
   U714 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n805, Z => n1108);
   U716 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n806, Z => n1109);
   U718 : MUXB2DL port map( A0 => n1381, A1 => n1398, SL => n807, Z => n1110);
   U721 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n808, Z => n1111);
   U723 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n809, Z => n1112);
   U725 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n810, Z => n1113);
   U727 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n811, Z => n1114);
   U729 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n812, Z => n1115);
   U731 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n813, Z => n1116);
   U733 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n814, Z => n1117);
   U735 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n815, Z => n1118);
   U737 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n816, Z => n1119);
   U739 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n817, Z => n1120);
   U741 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n818, Z => n1121);
   U743 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n819, Z => n1122);
   U745 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n820, Z => n1123);
   U747 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n821, Z => n1124);
   U749 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n822, Z => n1125);
   U751 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n823, Z => n1126);
   U753 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n824, Z => n1127);
   U755 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n825, Z => n1128);
   U757 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n826, Z => n1129);
   U759 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n827, Z => n1130);
   U761 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n828, Z => n1131);
   U763 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n829, Z => n1132);
   U765 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n830, Z => n1133);
   U767 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n831, Z => n1134);
   U769 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n832, Z => n1135);
   U771 : MUXB2DL port map( A0 => n1380, A1 => n1396, SL => n833, Z => n1136);
   U774 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n834, Z => n1137);
   U776 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n835, Z => n1138);
   U778 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n836, Z => n1139);
   U780 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n837, Z => n1140);
   U782 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n838, Z => n1141);
   U784 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n839, Z => n1142);
   U786 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n840, Z => n1143);
   U788 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n841, Z => n1144);
   U790 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n842, Z => n1145);
   U792 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n843, Z => n1146);
   U794 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n844, Z => n1147);
   U796 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n845, Z => n1148);
   U798 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n846, Z => n1149);
   U800 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n847, Z => n1150);
   U802 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n848, Z => n1151);
   U804 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n849, Z => n1152);
   U806 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n850, Z => n1153);
   U808 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n851, Z => n1154);
   U810 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n852, Z => n1155);
   U812 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n853, Z => n1156);
   U814 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n854, Z => n1157);
   U816 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n855, Z => n1158);
   U818 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n856, Z => n1159);
   U820 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n857, Z => n1160);
   U822 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n858, Z => n1161);
   U824 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n859, Z => n1162);
   U826 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n860, Z => n1163);
   U828 : MUXB2DL port map( A0 => n1377, A1 => n1394, SL => n861, Z => n1164);
   U831 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n862, Z => n1165);
   U833 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n863, Z => n1166);
   U835 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n864, Z => n1167);
   U837 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n865, Z => n1168);
   U839 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n866, Z => n1169);
   U841 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n867, Z => n1170);
   U843 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n868, Z => n1171);
   U845 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n869, Z => n1172);
   U847 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n870, Z => n1173);
   U849 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n871, Z => n1174);
   U851 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n872, Z => n1175);
   U853 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n873, Z => n1176);
   U855 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n874, Z => n1177);
   U857 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n875, Z => n1178);
   U859 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n876, Z => n1179);
   U861 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n877, Z => n1180);
   U863 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n878, Z => n1181);
   U865 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n879, Z => n1182);
   U867 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n880, Z => n1183);
   U869 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n881, Z => n1184);
   U871 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n882, Z => n1185);
   U873 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n883, Z => n1186);
   U875 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n884, Z => n1187);
   U877 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n885, Z => n1188);
   U879 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n886, Z => n1189);
   U881 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n887, Z => n1190);
   U883 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n888, Z => n1191);
   U885 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n889, Z => n1192);
   U887 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n890, Z => n1193);
   U889 : MUXB2DL port map( A0 => n1376, A1 => n1393, SL => n891, Z => n1194);
   U892 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n892, Z => n1195);
   U894 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n893, Z => n1196);
   U896 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n894, Z => n1197);
   U898 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n895, Z => n1198);
   U900 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n896, Z => n1199);
   U902 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n897, Z => n1200);
   U904 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n898, Z => n1201);
   U906 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n899, Z => n1202);
   U908 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n900, Z => n1203);
   U910 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n901, Z => n1204);
   U912 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n902, Z => n1205);
   U914 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n903, Z => n1206);
   U916 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n904, Z => n1207);
   U918 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n905, Z => n1208);
   U920 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n906, Z => n1209);
   U922 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n907, Z => n1210);
   U924 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n908, Z => n1211);
   U926 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n909, Z => n1212);
   U928 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n910, Z => n1213);
   U930 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n911, Z => n1214);
   U932 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n912, Z => n1215);
   U934 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n913, Z => n1216);
   U936 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n914, Z => n1217);
   U938 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n915, Z => n1218);
   U940 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n916, Z => n1219);
   U942 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n917, Z => n1220);
   U944 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n918, Z => n1221);
   U946 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n919, Z => n1222);
   U948 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n920, Z => n1223);
   U950 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n921, Z => n1224);
   U952 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n922, Z => n1225);
   U954 : MUXB2DL port map( A0 => n1375, A1 => n1392, SL => n923, Z => n1226);
   U1021 : NAN2D1 port map( A1 => n1390, A2 => n1392, Z => n1375);
   U1022 : OAI21D1 port map( A1 => a(2), A2 => a(1), B => n1395, Z => n1376);
   U1023 : OAI21D1 port map( A1 => a(4), A2 => a(3), B => n1397, Z => n1377);
   U1024 : EXOR2D1 port map( A1 => a(6), A2 => a(5), Z => n1378);
   U1025 : EXOR2D1 port map( A1 => a(8), A2 => a(7), Z => n1379);
   U1026 : OAI21D1 port map( A1 => a(6), A2 => a(5), B => n1399, Z => n1380);
   U1027 : OAI21D1 port map( A1 => a(8), A2 => a(7), B => n1401, Z => n1381);
   U1028 : INVD1 port map( A => n1382, Z => n1384);
   U1029 : INVD1 port map( A => n1383, Z => n1385);
   U1030 : INVD1 port map( A => n953, Z => n1393);
   U1031 : INVD1 port map( A => n952, Z => n1394);
   U1032 : INVD1 port map( A => n951, Z => n1396);
   U1033 : INVD1 port map( A => n950, Z => n1398);
   U1034 : INVD1 port map( A => n949, Z => n1400);
   U1035 : INVD1 port map( A => n948, Z => n1402);
   U1036 : INVD1 port map( A => n947, Z => n1404);
   U1037 : INVD1 port map( A => n946, Z => n1406);
   U1038 : INVD1 port map( A => n945, Z => n1408);
   U1039 : INVD1 port map( A => n944, Z => n1410);
   U1040 : INVD1 port map( A => n943, Z => n1412);
   U1041 : INVD1 port map( A => n942, Z => n1414);
   U1042 : INVD1 port map( A => n941, Z => n1416);
   U1043 : INVD1 port map( A => n940, Z => n1419);
   U1044 : INVD1 port map( A => n939, Z => n1420);
   U1045 : INVD1 port map( A => n1391, Z => n1390);
   U1046 : INVD1 port map( A => a(1), Z => n1392);
   U1047 : EXNOR2D1 port map( A1 => a(2), A2 => a(1), Z => n1382);
   U1048 : INVD1 port map( A => n1389, Z => n1388);
   U1049 : EXNOR2D1 port map( A1 => a(4), A2 => a(3), Z => n1383);
   U1050 : INVD1 port map( A => n1387, Z => n1386);
   U1051 : INVD1 port map( A => a(3), Z => n1395);
   U1052 : INVD1 port map( A => a(5), Z => n1397);
   U1053 : INVD1 port map( A => a(7), Z => n1399);
   U1054 : INVD1 port map( A => a(9), Z => n1401);
   U1055 : EXOR2D1 port map( A1 => a(10), A2 => a(9), Z => n1441);
   U1056 : INVD1 port map( A => a(11), Z => n1403);
   U1057 : OAI21D1 port map( A1 => a(9), A2 => a(10), B => n1403, Z => n42);
   U1058 : EXOR2D1 port map( A1 => a(12), A2 => a(11), Z => n1442);
   U1059 : INVD1 port map( A => a(13), Z => n1405);
   U1060 : OAI21D1 port map( A1 => a(12), A2 => a(11), B => n1405, Z => n50);
   U1061 : EXOR2D1 port map( A1 => a(14), A2 => a(13), Z => n1443);
   U1062 : INVD1 port map( A => a(15), Z => n1407);
   U1063 : OAI21D1 port map( A1 => a(14), A2 => a(13), B => n1407, Z => n58);
   U1064 : EXOR2D1 port map( A1 => a(16), A2 => a(15), Z => n1444);
   U1065 : INVD1 port map( A => a(17), Z => n1409);
   U1066 : OAI21D1 port map( A1 => a(16), A2 => a(15), B => n1409, Z => n66);
   U1067 : EXOR2D1 port map( A1 => a(18), A2 => a(17), Z => n1445);
   U1068 : INVD1 port map( A => a(19), Z => n1411);
   U1069 : OAI21D1 port map( A1 => a(18), A2 => a(17), B => n1411, Z => n73);
   U1070 : EXOR2D1 port map( A1 => a(20), A2 => a(19), Z => n1446);
   U1071 : INVD1 port map( A => a(21), Z => n1413);
   U1072 : OAI21D1 port map( A1 => a(20), A2 => a(19), B => n1413, Z => n80);
   U1073 : EXOR2D1 port map( A1 => a(22), A2 => a(21), Z => n1447);
   U1074 : INVD1 port map( A => a(23), Z => n1415);
   U1075 : OAI21D1 port map( A1 => a(22), A2 => a(21), B => n1415, Z => n84);
   U1076 : INVD1 port map( A => a(25), Z => n1417);
   U1077 : INVD1 port map( A => a(27), Z => n1418);
   U1078 : INVD1 port map( A => a(29), Z => n1421);
   U1079 : MUXB2DL port map( A0 => b(29), A1 => b(28), SL => n1382, Z => n862);
   U1080 : INVD1 port map( A => a(0), Z => n1391);
   U1081 : INVD1 port map( A => b(1), Z => n1389);
   U1082 : INVD1 port map( A => b(3), Z => n1387);
   U1083 : INVD1 port map( A => a(31), Z => n1422);
   U1084 : EXOR3D1 port map( A1 => n1423, A2 => n1424, A3 => n1425, Z => 
                           product(31));
   U1085 : EXOR3D1 port map( A1 => n208, A2 => n206, A3 => n1426, Z => n1425);
   U1086 : EXOR2D1 port map( A1 => n214, A2 => n212, Z => n1426);
   U1087 : EXOR2D1 port map( A1 => n202, A2 => n156, Z => n1424);
   U1088 : EXOR3D1 port map( A1 => n1427, A2 => n1428, A3 => n1429, Z => n1423)
                           ;
   U1089 : EXOR3D1 port map( A1 => n957, A2 => n955, A3 => n1430, Z => n1429);
   U1090 : EXNOR2D1 port map( A1 => n997, A2 => n975, Z => n1430);
   U1091 : EXOR3D1 port map( A1 => n1431, A2 => n204, A3 => n1432, Z => n1428);
   U1092 : EXOR3D1 port map( A1 => n1087, A2 => n1065, A3 => n1433, Z => n1432)
                           ;
   U1093 : EXNOR2D1 port map( A1 => n210, A2 => n1111, Z => n1433);
   U1094 : EXOR3D1 port map( A1 => n961, A2 => n218, A3 => n1434, Z => n1431);
   U1095 : EXOR2D1 port map( A1 => n985, A2 => n967, Z => n1434);
   U1096 : EXOR3D1 port map( A1 => n1435, A2 => n1436, A3 => n1437, Z => n1427)
                           ;
   U1097 : EXOR3D1 port map( A1 => n1027, A2 => n1011, A3 => n1438, Z => n1437)
                           ;
   U1098 : EXOR3D1 port map( A1 => n1165, A2 => n1137, A3 => n1045, Z => n1438)
                           ;
   U1099 : EXOR3D1 port map( A1 => n216, A2 => n1195, A3 => n1439, Z => n1436);
   U1100 : EXOR2D1 port map( A1 => n222, A2 => n220, Z => n1439);
   U1101 : EXOR3D1 port map( A1 => n226, A2 => n224, A3 => n1440, Z => n1435);
   U1102 : EXOR2D1 port map( A1 => n230, A2 => n228, Z => n1440);
   U1103 : OAI21D1 port map( A1 => a(28), A2 => a(27), B => n1421, Z => n99);
   U1104 : AOI21D1 port map( A1 => a(25), A2 => a(26), B => n1418, Z => n941);
   U1105 : OAI21D1 port map( A1 => a(26), A2 => a(25), B => n1418, Z => n94);
   U1106 : NAN2D1 port map( A1 => b(0), A2 => n1390, Z => n923);
   U1107 : MUXB2DL port map( A0 => b(0), A1 => n1388, SL => n1390, Z => n922);
   U1108 : MUXB2DL port map( A0 => n1388, A1 => b(2), SL => n1390, Z => n921);
   U1109 : MUXB2DL port map( A0 => b(2), A1 => n1386, SL => n1390, Z => n920);
   U1110 : MUXB2DL port map( A0 => n1386, A1 => b(4), SL => n1390, Z => n919);
   U1111 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1390, Z => n918);
   U1112 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1390, Z => n917);
   U1113 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1390, Z => n916);
   U1114 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1390, Z => n915);
   U1115 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1390, Z => n914);
   U1116 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1390, Z => n913);
   U1117 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1390, Z => n912);
   U1118 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1390, Z => n911);
   U1119 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1390, Z => n910);
   U1120 : AOI21D1 port map( A1 => a(23), A2 => a(24), B => n1417, Z => n942);
   U1121 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => a(0), Z => n909);
   U1122 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => a(0), Z => n908);
   U1123 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => a(0), Z => n907);
   U1124 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => a(0), Z => n906);
   U1125 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => a(0), Z => n905);
   U1126 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => a(0), Z => n904);
   U1127 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => a(0), Z => n903);
   U1128 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => a(0), Z => n902);
   U1129 : MUXB2DL port map( A0 => b(21), A1 => b(22), SL => a(0), Z => n901);
   U1130 : MUXB2DL port map( A0 => b(22), A1 => b(23), SL => a(0), Z => n900);
   U1131 : MUXB2DL port map( A0 => b(23), A1 => b(24), SL => a(0), Z => n899);
   U1132 : MUXB2DL port map( A0 => b(24), A1 => b(25), SL => a(0), Z => n898);
   U1133 : MUXB2DL port map( A0 => b(25), A1 => b(26), SL => a(0), Z => n897);
   U1134 : MUXB2DL port map( A0 => b(26), A1 => b(27), SL => a(0), Z => n896);
   U1135 : MUXB2DL port map( A0 => b(27), A1 => b(28), SL => a(0), Z => n895);
   U1136 : MUXB2DL port map( A0 => b(28), A1 => b(29), SL => a(0), Z => n894);
   U1137 : MUXB2DL port map( A0 => b(29), A1 => b(30), SL => a(0), Z => n893);
   U1138 : MUXB2DL port map( A0 => b(30), A1 => b(31), SL => n1390, Z => n892);
   U1139 : NAN2D1 port map( A1 => b(0), A2 => n1384, Z => n891);
   U1140 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1384, Z => n890);
   U1141 : OAI21D1 port map( A1 => a(24), A2 => a(23), B => n1417, Z => n89);
   U1142 : MUXB2DL port map( A0 => n1388, A1 => b(2), SL => n1384, Z => n889);
   U1143 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1384, Z => n888);
   U1144 : MUXB2DL port map( A0 => n1386, A1 => b(4), SL => n1384, Z => n887);
   U1145 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1384, Z => n886);
   U1146 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1384, Z => n885);
   U1147 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1384, Z => n884);
   U1148 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1384, Z => n883);
   U1149 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1384, Z => n882);
   U1150 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1384, Z => n881);
   U1151 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1384, Z => n880);
   U1152 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1384, Z => n879);
   U1153 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1384, Z => n878);
   U1154 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1384, Z => n877);
   U1155 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1384, Z => n876);
   U1156 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1384, Z => n875);
   U1157 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1384, Z => n874);
   U1158 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1384, Z => n873);
   U1159 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1384, Z => n872);
   U1160 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => n1384, Z => n871);
   U1161 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => n1384, Z => n870);
   U1162 : MUXB2DL port map( A0 => b(21), A1 => b(22), SL => n1384, Z => n869);
   U1163 : MUXB2DL port map( A0 => b(22), A1 => b(23), SL => n1384, Z => n868);
   U1164 : MUXB2DL port map( A0 => b(23), A1 => b(24), SL => n1384, Z => n867);
   U1165 : MUXB2DL port map( A0 => b(24), A1 => b(25), SL => n1384, Z => n866);
   U1166 : MUXB2DL port map( A0 => b(25), A1 => b(26), SL => n1384, Z => n865);
   U1167 : MUXB2DL port map( A0 => b(26), A1 => b(27), SL => n1384, Z => n864);
   U1168 : MUXB2DL port map( A0 => b(27), A1 => b(28), SL => n1384, Z => n863);
   U1169 : NAN2D1 port map( A1 => b(0), A2 => n1385, Z => n861);
   U1170 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1385, Z => n860);
   U1171 : AOI21D1 port map( A1 => a(21), A2 => a(22), B => n1415, Z => n943);
   U1172 : MUXB2DL port map( A0 => n1388, A1 => b(2), SL => n1385, Z => n859);
   U1173 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1385, Z => n858);
   U1174 : MUXB2DL port map( A0 => n1386, A1 => b(4), SL => n1385, Z => n857);
   U1175 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1385, Z => n856);
   U1176 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1385, Z => n855);
   U1177 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1385, Z => n854);
   U1178 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1385, Z => n853);
   U1179 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1385, Z => n852);
   U1180 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1385, Z => n851);
   U1181 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1385, Z => n850);
   U1182 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1385, Z => n849);
   U1183 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1385, Z => n848);
   U1184 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1385, Z => n847);
   U1185 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1385, Z => n846);
   U1186 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1385, Z => n845);
   U1187 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1385, Z => n844);
   U1188 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1385, Z => n843);
   U1189 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1385, Z => n842);
   U1190 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => n1385, Z => n841);
   U1191 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => n1385, Z => n840);
   U1192 : MUXB2DL port map( A0 => b(21), A1 => b(22), SL => n1385, Z => n839);
   U1193 : MUXB2DL port map( A0 => b(22), A1 => b(23), SL => n1385, Z => n838);
   U1194 : MUXB2DL port map( A0 => b(23), A1 => b(24), SL => n1385, Z => n837);
   U1195 : MUXB2DL port map( A0 => b(24), A1 => b(25), SL => n1385, Z => n836);
   U1196 : MUXB2DL port map( A0 => b(25), A1 => b(26), SL => n1385, Z => n835);
   U1197 : MUXB2DL port map( A0 => b(26), A1 => b(27), SL => n1385, Z => n834);
   U1198 : NAN2D1 port map( A1 => b(0), A2 => n1378, Z => n833);
   U1199 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1378, Z => n832);
   U1200 : MUXB2DL port map( A0 => n1388, A1 => b(2), SL => n1378, Z => n831);
   U1201 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1378, Z => n830);
   U1202 : MUXB2DL port map( A0 => n1386, A1 => b(4), SL => n1378, Z => n829);
   U1203 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1378, Z => n828);
   U1204 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1378, Z => n827);
   U1205 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1378, Z => n826);
   U1206 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1378, Z => n825);
   U1207 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1378, Z => n824);
   U1208 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1378, Z => n823);
   U1209 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1378, Z => n822);
   U1210 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1378, Z => n821);
   U1211 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1378, Z => n820);
   U1212 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1378, Z => n819);
   U1213 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1378, Z => n818);
   U1214 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1378, Z => n817);
   U1215 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1378, Z => n816);
   U1216 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1378, Z => n815);
   U1217 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1378, Z => n814);
   U1218 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => n1378, Z => n813);
   U1219 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => n1378, Z => n812);
   U1220 : MUXB2DL port map( A0 => b(21), A1 => b(22), SL => n1378, Z => n811);
   U1221 : MUXB2DL port map( A0 => b(22), A1 => b(23), SL => n1378, Z => n810);
   U1222 : AOI21D1 port map( A1 => a(19), A2 => a(20), B => n1413, Z => n944);
   U1223 : MUXB2DL port map( A0 => b(23), A1 => b(24), SL => n1378, Z => n809);
   U1224 : MUXB2DL port map( A0 => b(24), A1 => b(25), SL => n1378, Z => n808);
   U1225 : NAN2D1 port map( A1 => b(0), A2 => n1379, Z => n807);
   U1226 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1379, Z => n806);
   U1227 : MUXB2DL port map( A0 => b(1), A1 => b(2), SL => n1379, Z => n805);
   U1228 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1379, Z => n804);
   U1229 : MUXB2DL port map( A0 => n1386, A1 => b(4), SL => n1379, Z => n803);
   U1230 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1379, Z => n802);
   U1231 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1379, Z => n801);
   U1232 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1379, Z => n800);
   U1233 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1379, Z => n799);
   U1234 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1379, Z => n798);
   U1235 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1379, Z => n797);
   U1236 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1379, Z => n796);
   U1237 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1379, Z => n795);
   U1238 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1379, Z => n794);
   U1239 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1379, Z => n793);
   U1240 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1379, Z => n792);
   U1241 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1379, Z => n791);
   U1242 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1379, Z => n790);
   U1243 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1379, Z => n789);
   U1244 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1379, Z => n788);
   U1245 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => n1379, Z => n787);
   U1246 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => n1379, Z => n786);
   U1247 : MUXB2DL port map( A0 => b(21), A1 => b(22), SL => n1379, Z => n785);
   U1248 : MUXB2DL port map( A0 => b(22), A1 => b(23), SL => n1379, Z => n784);
   U1249 : NAN2D1 port map( A1 => b(0), A2 => n1441, Z => n783);
   U1250 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1441, Z => n782);
   U1251 : MUXB2DL port map( A0 => n1388, A1 => b(2), SL => n1441, Z => n781);
   U1252 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1441, Z => n780);
   U1253 : MUXB2DL port map( A0 => b(3), A1 => b(4), SL => n1441, Z => n779);
   U1254 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1441, Z => n778);
   U1255 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1441, Z => n777);
   U1256 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1441, Z => n776);
   U1257 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1441, Z => n775);
   U1258 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1441, Z => n774);
   U1259 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1441, Z => n773);
   U1260 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1441, Z => n772);
   U1261 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1441, Z => n771);
   U1262 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1441, Z => n770);
   U1263 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1441, Z => n769);
   U1264 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1441, Z => n768);
   U1265 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1441, Z => n767);
   U1266 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1441, Z => n766);
   U1267 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1441, Z => n765);
   U1268 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1441, Z => n764);
   U1269 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => n1441, Z => n763);
   U1270 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => n1441, Z => n762);
   U1271 : NAN2D1 port map( A1 => b(0), A2 => n1442, Z => n761);
   U1272 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1442, Z => n760);
   U1273 : MUXB2DL port map( A0 => b(1), A1 => b(2), SL => n1442, Z => n759);
   U1274 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1442, Z => n758);
   U1275 : MUXB2DL port map( A0 => n1386, A1 => b(4), SL => n1442, Z => n757);
   U1276 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1442, Z => n756);
   U1277 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1442, Z => n755);
   U1278 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1442, Z => n754);
   U1279 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1442, Z => n753);
   U1280 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1442, Z => n752);
   U1281 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1442, Z => n751);
   U1282 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1442, Z => n750);
   U1283 : AOI21D1 port map( A1 => a(17), A2 => a(18), B => n1411, Z => n945);
   U1284 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1442, Z => n749);
   U1285 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1442, Z => n748);
   U1286 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1442, Z => n747);
   U1287 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1442, Z => n746);
   U1288 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1442, Z => n745);
   U1289 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1442, Z => n744);
   U1290 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1442, Z => n743);
   U1291 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1442, Z => n742);
   U1292 : NAN2D1 port map( A1 => b(0), A2 => n1443, Z => n741);
   U1293 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1443, Z => n740);
   U1294 : MUXB2DL port map( A0 => n1388, A1 => b(2), SL => n1443, Z => n739);
   U1295 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1443, Z => n738);
   U1296 : MUXB2DL port map( A0 => n1386, A1 => b(4), SL => n1443, Z => n737);
   U1297 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1443, Z => n736);
   U1298 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1443, Z => n735);
   U1299 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1443, Z => n734);
   U1300 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1443, Z => n733);
   U1301 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1443, Z => n732);
   U1302 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1443, Z => n731);
   U1303 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1443, Z => n730);
   U1304 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1443, Z => n729);
   U1305 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1443, Z => n728);
   U1306 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1443, Z => n727);
   U1307 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1443, Z => n726);
   U1308 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1443, Z => n725);
   U1309 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1443, Z => n724);
   U1310 : NAN2D1 port map( A1 => b(0), A2 => n1444, Z => n723);
   U1311 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1444, Z => n722);
   U1312 : MUXB2DL port map( A0 => n1388, A1 => b(2), SL => n1444, Z => n721);
   U1313 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1444, Z => n720);
   U1314 : MUXB2DL port map( A0 => n1386, A1 => b(4), SL => n1444, Z => n719);
   U1315 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1444, Z => n718);
   U1316 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1444, Z => n717);
   U1317 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1444, Z => n716);
   U1318 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1444, Z => n715);
   U1319 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1444, Z => n714);
   U1320 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1444, Z => n713);
   U1321 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1444, Z => n712);
   U1322 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1444, Z => n711);
   U1323 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1444, Z => n710);
   U1324 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1444, Z => n709);
   U1325 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1444, Z => n708);
   U1326 : NAN2D1 port map( A1 => b(0), A2 => n1445, Z => n707);
   U1327 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1445, Z => n706);
   U1328 : MUXB2DL port map( A0 => n1388, A1 => b(2), SL => n1445, Z => n705);
   U1329 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1445, Z => n704);
   U1330 : MUXB2DL port map( A0 => n1386, A1 => b(4), SL => n1445, Z => n703);
   U1331 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1445, Z => n702);
   U1332 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1445, Z => n701);
   U1333 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1445, Z => n700);
   U1334 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1445, Z => n699);
   U1335 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1445, Z => n698);
   U1336 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1445, Z => n697);
   U1337 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1445, Z => n696);
   U1338 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1445, Z => n695);
   U1339 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1445, Z => n694);
   U1340 : NAN2D1 port map( A1 => b(0), A2 => n1446, Z => n693);
   U1341 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1446, Z => n692);
   U1342 : MUXB2DL port map( A0 => n1388, A1 => b(2), SL => n1446, Z => n691);
   U1343 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1446, Z => n690);
   U1344 : MUXB2DL port map( A0 => n1386, A1 => b(4), SL => n1446, Z => n689);
   U1345 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1446, Z => n688);
   U1346 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1446, Z => n687);
   U1347 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1446, Z => n686);
   U1348 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1446, Z => n685);
   U1349 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1446, Z => n684);
   U1350 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1446, Z => n683);
   U1351 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1446, Z => n682);
   U1352 : NAN2D1 port map( A1 => b(0), A2 => n1447, Z => n681);
   U1353 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1447, Z => n680);
   U1354 : AOI21D1 port map( A1 => a(15), A2 => a(16), B => n1409, Z => n946);
   U1355 : MUXB2DL port map( A0 => n1388, A1 => b(2), SL => n1447, Z => n679);
   U1356 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1447, Z => n678);
   U1357 : MUXB2DL port map( A0 => n1386, A1 => b(4), SL => n1447, Z => n677);
   U1358 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1447, Z => n676);
   U1359 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1447, Z => n675);
   U1360 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1447, Z => n674);
   U1361 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1447, Z => n673);
   U1362 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1447, Z => n672);
   U1363 : NAN2D1 port map( A1 => b(0), A2 => n1448, Z => n671);
   U1364 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1448, Z => n670);
   U1365 : MUXB2DL port map( A0 => n1388, A1 => b(2), SL => n1448, Z => n669);
   U1366 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1448, Z => n668);
   U1367 : MUXB2DL port map( A0 => n1386, A1 => b(4), SL => n1448, Z => n667);
   U1368 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1448, Z => n666);
   U1369 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1448, Z => n665);
   U1370 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1448, Z => n664);
   U1371 : EXOR2D1 port map( A1 => a(24), A2 => a(23), Z => n1448);
   U1372 : NAN2D1 port map( A1 => b(0), A2 => n1449, Z => n663);
   U1373 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1449, Z => n662);
   U1374 : MUXB2DL port map( A0 => n1388, A1 => b(2), SL => n1449, Z => n661);
   U1375 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1449, Z => n660);
   U1376 : MUXB2DL port map( A0 => n1386, A1 => b(4), SL => n1449, Z => n659);
   U1377 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1449, Z => n658);
   U1378 : EXOR2D1 port map( A1 => a(26), A2 => a(25), Z => n1449);
   U1379 : NAN2D1 port map( A1 => b(0), A2 => n1450, Z => n657);
   U1380 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1450, Z => n656);
   U1381 : MUXB2DL port map( A0 => n1388, A1 => b(2), SL => n1450, Z => n655);
   U1382 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1450, Z => n654);
   U1383 : EXOR2D1 port map( A1 => a(28), A2 => a(27), Z => n1450);
   U1384 : NAN2D1 port map( A1 => b(0), A2 => n1451, Z => n653);
   U1385 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1451, Z => n652);
   U1386 : EXOR2D1 port map( A1 => a(30), A2 => a(29), Z => n1451);
   U1387 : AOI21D1 port map( A1 => a(13), A2 => a(14), B => n1407, Z => n947);
   U1388 : AOI21D1 port map( A1 => a(11), A2 => a(12), B => n1405, Z => n948);
   U1389 : AOI21D1 port map( A1 => a(9), A2 => a(10), B => n1403, Z => n949);
   U1390 : AOI21D1 port map( A1 => a(7), A2 => a(8), B => n1401, Z => n950);
   U1391 : AOI21D1 port map( A1 => a(5), A2 => a(6), B => n1399, Z => n951);
   U1392 : AOI21D1 port map( A1 => a(3), A2 => a(4), B => n1397, Z => n952);
   U1393 : AOI21D1 port map( A1 => a(1), A2 => a(2), B => n1395, Z => n953);
   U1394 : AOI21D1 port map( A1 => a(29), A2 => a(30), B => n1422, Z => n939);
   U1395 : OAI21D1 port map( A1 => a(30), A2 => a(29), B => n1422, Z => n104);
   U1396 : AOI21D1 port map( A1 => a(27), A2 => a(28), B => n1421, Z => n940);

end hier_filter_none_20;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_gp_custom.all;

architecture hier_filter_none_20 of gp_custom_DW_mult_tc_1 is

   component AOI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component MUXB2DL
      port( A0, A1, SL : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal n42, n50, n58, n66, n73, n80, n84, n89, n94, n99, n104, n156, n157, 
      n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, 
      n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, 
      n182, n183, n184, n185, n186, n202, n203, n204, n205, n206, n207, n208, 
      n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, 
      n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, 
      n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, 
      n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, 
      n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, 
      n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, 
      n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
      n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, 
      n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, 
      n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, 
      n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, 
      n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, 
      n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, 
      n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, 
      n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, 
      n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, 
      n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, 
      n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, 
      n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, 
      n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, 
      n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, 
      n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, 
      n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, 
      n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, 
      n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, 
      n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, 
      n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
      n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, 
      n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, 
      n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, 
      n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
      n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, 
      n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, 
      n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, 
      n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, 
      n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, 
      n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, 
      n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, 
      n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, 
      n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, 
      n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, 
      n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, 
      n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, 
      n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, 
      n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, 
      n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, 
      n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, 
      n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, 
      n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, 
      n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, 
      n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, 
      n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, 
      n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, 
      n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, 
      n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, 
      n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, 
      n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, 
      n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, 
      n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, 
      n917, n918, n919, n920, n921, n922, n923, n939, n940, n941, n942, n943, 
      n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n955, n956, 
      n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, 
      n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, 
      n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, 
      n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, 
      n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, 
      n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, 
      n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, 
      n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, 
      n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, 
      n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, 
      n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, 
      n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, 
      n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, 
      n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, 
      n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, 
      n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, 
      n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, 
      n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, 
      n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, 
      n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, 
      n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, 
      n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, 
      n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, 
      n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, 
      n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, 
      n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, 
      n1224, n1225, n1226, n1375, n1376, n1377, n1378, n1379, n1380, n1381, 
      n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, 
      n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, 
      n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, 
      n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, 
      n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, 
      n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, 
      n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, 
      n1452, n1453, n1454, n1455, n1456, n1457 : std_logic;

begin
   
   U125 : ADFULD1 port map( A => n203, B => n232, CI => n157, CO => n156, S => 
                           product(30));
   U126 : ADFULD1 port map( A => n233, B => n260, CI => n158, CO => n157, S => 
                           product(29));
   U127 : ADFULD1 port map( A => n261, B => n288, CI => n159, CO => n158, S => 
                           product(28));
   U128 : ADFULD1 port map( A => n289, B => n314, CI => n160, CO => n159, S => 
                           product(27));
   U129 : ADFULD1 port map( A => n315, B => n340, CI => n161, CO => n160, S => 
                           product(26));
   U130 : ADFULD1 port map( A => n341, B => n364, CI => n162, CO => n161, S => 
                           product(25));
   U131 : ADFULD1 port map( A => n365, B => n388, CI => n163, CO => n162, S => 
                           product(24));
   U132 : ADFULD1 port map( A => n389, B => n410, CI => n164, CO => n163, S => 
                           product(23));
   U133 : ADFULD1 port map( A => n411, B => n432, CI => n165, CO => n164, S => 
                           product(22));
   U134 : ADFULD1 port map( A => n433, B => n452, CI => n166, CO => n165, S => 
                           product(21));
   U135 : ADFULD1 port map( A => n453, B => n472, CI => n167, CO => n166, S => 
                           product(20));
   U136 : ADFULD1 port map( A => n473, B => n490, CI => n168, CO => n167, S => 
                           product(19));
   U137 : ADFULD1 port map( A => n491, B => n508, CI => n169, CO => n168, S => 
                           product(18));
   U138 : ADFULD1 port map( A => n509, B => n524, CI => n170, CO => n169, S => 
                           product(17));
   U139 : ADFULD1 port map( A => n525, B => n540, CI => n171, CO => n170, S => 
                           product(16));
   U140 : ADFULD1 port map( A => n541, B => n554, CI => n172, CO => n171, S => 
                           product(15));
   U141 : ADFULD1 port map( A => n555, B => n568, CI => n173, CO => n172, S => 
                           product(14));
   U142 : ADFULD1 port map( A => n569, B => n580, CI => n174, CO => n173, S => 
                           product(13));
   U143 : ADFULD1 port map( A => n581, B => n592, CI => n175, CO => n174, S => 
                           product(12));
   U144 : ADFULD1 port map( A => n593, B => n602, CI => n176, CO => n175, S => 
                           product(11));
   U145 : ADFULD1 port map( A => n603, B => n612, CI => n177, CO => n176, S => 
                           product(10));
   U146 : ADFULD1 port map( A => n613, B => n620, CI => n178, CO => n177, S => 
                           product(9));
   U147 : ADFULD1 port map( A => n621, B => n628, CI => n179, CO => n178, S => 
                           product(8));
   U148 : ADFULD1 port map( A => n629, B => n634, CI => n180, CO => n179, S => 
                           product(7));
   U149 : ADFULD1 port map( A => n635, B => n640, CI => n181, CO => n180, S => 
                           product(6));
   U150 : ADFULD1 port map( A => n641, B => n644, CI => n182, CO => n181, S => 
                           product(5));
   U151 : ADFULD1 port map( A => n645, B => n648, CI => n183, CO => n182, S => 
                           product(4));
   U152 : ADFULD1 port map( A => n649, B => n1193, CI => n184, CO => n183, S =>
                           product(3));
   U153 : ADFULD1 port map( A => n651, B => n1194, CI => n185, CO => n184, S =>
                           product(2));
   U154 : ADHALFDL port map( A => n186, B => n1225, CO => n185, S => product(1)
                           );
   U155 : ADHALFDL port map( A => n1226, B => a(1), CO => n186, S => product(0)
                           );
   U171 : ADFULD1 port map( A => n234, B => n207, CI => n205, CO => n202, S => 
                           n203);
   U172 : ADFULD1 port map( A => n209, B => n211, CI => n236, CO => n204, S => 
                           n205);
   U173 : ADFULD1 port map( A => n240, B => n213, CI => n238, CO => n206, S => 
                           n207);
   U174 : ADFULD1 port map( A => n217, B => n242, CI => n215, CO => n208, S => 
                           n209);
   U175 : ADFULD1 port map( A => n244, B => n246, CI => n219, CO => n210, S => 
                           n211);
   U176 : ADFULD1 port map( A => n225, B => n223, CI => n248, CO => n212, S => 
                           n213);
   U177 : ADFULD1 port map( A => n221, B => n229, CI => n227, CO => n214, S => 
                           n215);
   U178 : ADFULD1 port map( A => n256, B => n252, CI => n254, CO => n216, S => 
                           n217);
   U179 : ADFULD1 port map( A => n258, B => n1088, CI => n250, CO => n218, S =>
                           n219);
   U180 : ADFULD1 port map( A => n1046, B => n1112, CI => n1066, CO => n220, S 
                           => n221);
   U181 : ADFULD1 port map( A => n986, B => n976, CI => n998, CO => n222, S => 
                           n223);
   U182 : ADFULD1 port map( A => n962, B => n1138, CI => n968, CO => n224, S =>
                           n225);
   U183 : ADFULD1 port map( A => n1166, B => n1012, CI => n231, CO => n226, S 
                           => n227);
   U184 : ADFULD1 port map( A => n1028, B => n956, CI => n958, CO => n228, S =>
                           n229);
   U185 : ADHALFDL port map( A => n1196, B => n939, CO => n230, S => n231);
   U186 : ADFULD1 port map( A => n262, B => n237, CI => n235, CO => n232, S => 
                           n233);
   U187 : ADFULD1 port map( A => n239, B => n266, CI => n264, CO => n234, S => 
                           n235);
   U188 : ADFULD1 port map( A => n268, B => n243, CI => n241, CO => n236, S => 
                           n237);
   U189 : ADFULD1 port map( A => n270, B => n247, CI => n245, CO => n238, S => 
                           n239);
   U190 : ADFULD1 port map( A => n274, B => n249, CI => n272, CO => n240, S => 
                           n241);
   U191 : ADFULD1 port map( A => n253, B => n255, CI => n257, CO => n242, S => 
                           n243);
   U192 : ADFULD1 port map( A => n280, B => n276, CI => n251, CO => n244, S => 
                           n245);
   U193 : ADFULD1 port map( A => n278, B => n284, CI => n282, CO => n246, S => 
                           n247);
   U194 : ADFULD1 port map( A => n1047, B => n1013, CI => n259, CO => n248, S 
                           => n249);
   U195 : ADFULD1 port map( A => n977, B => n1067, CI => n999, CO => n250, S =>
                           n251);
   U196 : ADFULD1 port map( A => n959, B => n969, CI => n963, CO => n252, S => 
                           n253);
   U197 : ADFULD1 port map( A => n1113, B => n987, CI => n1089, CO => n254, S 
                           => n255);
   U198 : ADFULD1 port map( A => n1167, B => n1029, CI => n1139, CO => n256, S 
                           => n257);
   U199 : ADHALFDL port map( A => n286, B => n1197, CO => n258, S => n259);
   U200 : ADFULD1 port map( A => n290, B => n265, CI => n263, CO => n260, S => 
                           n261);
   U201 : ADFULD1 port map( A => n267, B => n294, CI => n292, CO => n262, S => 
                           n263);
   U202 : ADFULD1 port map( A => n296, B => n271, CI => n269, CO => n264, S => 
                           n265);
   U203 : ADFULD1 port map( A => n275, B => n298, CI => n273, CO => n266, S => 
                           n267);
   U204 : ADFULD1 port map( A => n302, B => n281, CI => n300, CO => n268, S => 
                           n269);
   U205 : ADFULD1 port map( A => n283, B => n277, CI => n279, CO => n270, S => 
                           n271);
   U206 : ADFULD1 port map( A => n310, B => n308, CI => n285, CO => n272, S => 
                           n273);
   U207 : ADFULD1 port map( A => n304, B => n312, CI => n306, CO => n274, S => 
                           n275);
   U208 : ADFULD1 port map( A => n1014, B => n1068, CI => n1048, CO => n276, S 
                           => n277);
   U209 : ADFULD1 port map( A => n978, B => n1090, CI => n988, CO => n278, S =>
                           n279);
   U210 : ADFULD1 port map( A => n964, B => n1114, CI => n970, CO => n280, S =>
                           n281);
   U211 : ADFULD1 port map( A => n1140, B => n1000, CI => n287, CO => n282, S 
                           => n283);
   U212 : ADFULD1 port map( A => n1030, B => n960, CI => n1168, CO => n284, S 
                           => n285);
   U213 : ADHALFDL port map( A => n1198, B => n940, CO => n286, S => n287);
   U214 : ADFULD1 port map( A => n316, B => n293, CI => n291, CO => n288, S => 
                           n289);
   U215 : ADFULD1 port map( A => n318, B => n297, CI => n295, CO => n290, S => 
                           n291);
   U216 : ADFULD1 port map( A => n299, B => n322, CI => n320, CO => n292, S => 
                           n293);
   U217 : ADFULD1 port map( A => n324, B => n303, CI => n301, CO => n294, S => 
                           n295);
   U218 : ADFULD1 port map( A => n307, B => n309, CI => n326, CO => n296, S => 
                           n297);
   U219 : ADFULD1 port map( A => n305, B => n328, CI => n311, CO => n298, S => 
                           n299);
   U220 : ADFULD1 port map( A => n332, B => n330, CI => n334, CO => n300, S => 
                           n301);
   U221 : ADFULD1 port map( A => n313, B => n1091, CI => n336, CO => n302, S =>
                           n303);
   U222 : ADFULD1 port map( A => n1015, B => n1115, CI => n1069, CO => n304, S 
                           => n305);
   U223 : ADFULD1 port map( A => n1141, B => n1001, CI => n989, CO => n306, S 
                           => n307);
   U224 : ADFULD1 port map( A => n979, B => n1049, CI => n1169, CO => n308, S 
                           => n309);
   U225 : ADFULD1 port map( A => n965, B => n1031, CI => n971, CO => n310, S =>
                           n311);
   U226 : ADHALFDL port map( A => n338, B => n1199, CO => n312, S => n313);
   U227 : ADFULD1 port map( A => n342, B => n319, CI => n317, CO => n314, S => 
                           n315);
   U228 : ADFULD1 port map( A => n344, B => n346, CI => n321, CO => n316, S => 
                           n317);
   U229 : ADFULD1 port map( A => n325, B => n327, CI => n323, CO => n318, S => 
                           n319);
   U230 : ADFULD1 port map( A => n350, B => n352, CI => n348, CO => n320, S => 
                           n321);
   U231 : ADFULD1 port map( A => n333, B => n335, CI => n329, CO => n322, S => 
                           n323);
   U232 : ADFULD1 port map( A => n337, B => n358, CI => n331, CO => n324, S => 
                           n325);
   U233 : ADFULD1 port map( A => n354, B => n360, CI => n356, CO => n326, S => 
                           n327);
   U234 : ADFULD1 port map( A => n1092, B => n1116, CI => n362, CO => n328, S 
                           => n329);
   U235 : ADFULD1 port map( A => n1016, B => n1142, CI => n1070, CO => n330, S 
                           => n331);
   U236 : ADFULD1 port map( A => n990, B => n1170, CI => n1002, CO => n332, S 
                           => n333);
   U237 : ADFULD1 port map( A => n980, B => n1032, CI => n339, CO => n334, S =>
                           n335);
   U238 : ADFULD1 port map( A => n1050, B => n966, CI => n972, CO => n336, S =>
                           n337);
   U239 : ADHALFDL port map( A => n1200, B => n941, CO => n338, S => n339);
   U240 : ADFULD1 port map( A => n366, B => n345, CI => n343, CO => n340, S => 
                           n341);
   U241 : ADFULD1 port map( A => n347, B => n370, CI => n368, CO => n342, S => 
                           n343);
   U242 : ADFULD1 port map( A => n351, B => n372, CI => n349, CO => n344, S => 
                           n345);
   U243 : ADFULD1 port map( A => n374, B => n376, CI => n353, CO => n346, S => 
                           n347);
   U244 : ADFULD1 port map( A => n361, B => n357, CI => n359, CO => n348, S => 
                           n349);
   U245 : ADFULD1 port map( A => n378, B => n380, CI => n355, CO => n350, S => 
                           n351);
   U246 : ADFULD1 port map( A => n384, B => n363, CI => n382, CO => n352, S => 
                           n353);
   U247 : ADFULD1 port map( A => n1033, B => n1093, CI => n1071, CO => n354, S 
                           => n355);
   U248 : ADFULD1 port map( A => n991, B => n1117, CI => n1017, CO => n356, S 
                           => n357);
   U249 : ADFULD1 port map( A => n973, B => n1003, CI => n981, CO => n358, S =>
                           n359);
   U250 : ADFULD1 port map( A => n1171, B => n1051, CI => n1143, CO => n360, S 
                           => n361);
   U251 : ADHALFDL port map( A => n386, B => n1201, CO => n362, S => n363);
   U252 : ADFULD1 port map( A => n390, B => n369, CI => n367, CO => n364, S => 
                           n365);
   U253 : ADFULD1 port map( A => n371, B => n394, CI => n392, CO => n366, S => 
                           n367);
   U254 : ADFULD1 port map( A => n375, B => n396, CI => n373, CO => n368, S => 
                           n369);
   U255 : ADFULD1 port map( A => n398, B => n400, CI => n377, CO => n370, S => 
                           n371);
   U256 : ADFULD1 port map( A => n383, B => n379, CI => n381, CO => n372, S => 
                           n373);
   U257 : ADFULD1 port map( A => n402, B => n404, CI => n385, CO => n374, S => 
                           n375);
   U258 : ADFULD1 port map( A => n408, B => n1072, CI => n406, CO => n376, S =>
                           n377);
   U259 : ADFULD1 port map( A => n1004, B => n1094, CI => n1034, CO => n378, S 
                           => n379);
   U260 : ADFULD1 port map( A => n992, B => n1144, CI => n1118, CO => n380, S 
                           => n381);
   U261 : ADFULD1 port map( A => n982, B => n1018, CI => n387, CO => n382, S =>
                           n383);
   U262 : ADFULD1 port map( A => n1052, B => n974, CI => n1172, CO => n384, S 
                           => n385);
   U263 : ADHALFDL port map( A => n1202, B => n942, CO => n386, S => n387);
   U264 : ADFULD1 port map( A => n412, B => n393, CI => n391, CO => n388, S => 
                           n389);
   U265 : ADFULD1 port map( A => n395, B => n397, CI => n414, CO => n390, S => 
                           n391);
   U266 : ADFULD1 port map( A => n399, B => n418, CI => n416, CO => n392, S => 
                           n393);
   U267 : ADFULD1 port map( A => n401, B => n407, CI => n420, CO => n394, S => 
                           n395);
   U268 : ADFULD1 port map( A => n403, B => n424, CI => n405, CO => n396, S => 
                           n397);
   U269 : ADFULD1 port map( A => n426, B => n428, CI => n422, CO => n398, S => 
                           n399);
   U270 : ADFULD1 port map( A => n1073, B => n1095, CI => n409, CO => n400, S 
                           => n401);
   U271 : ADFULD1 port map( A => n1005, B => n1119, CI => n1019, CO => n402, S 
                           => n403);
   U272 : ADFULD1 port map( A => n1173, B => n1035, CI => n1145, CO => n404, S 
                           => n405);
   U273 : ADFULD1 port map( A => n983, B => n1053, CI => n993, CO => n406, S =>
                           n407);
   U274 : ADHALFDL port map( A => n430, B => n1203, CO => n408, S => n409);
   U275 : ADFULD1 port map( A => n434, B => n415, CI => n413, CO => n410, S => 
                           n411);
   U276 : ADFULD1 port map( A => n417, B => n419, CI => n436, CO => n412, S => 
                           n413);
   U277 : ADFULD1 port map( A => n421, B => n440, CI => n438, CO => n414, S => 
                           n415);
   U278 : ADFULD1 port map( A => n427, B => n425, CI => n442, CO => n416, S => 
                           n417);
   U279 : ADFULD1 port map( A => n429, B => n444, CI => n423, CO => n418, S => 
                           n419);
   U280 : ADFULD1 port map( A => n448, B => n450, CI => n446, CO => n420, S => 
                           n421);
   U281 : ADFULD1 port map( A => n1074, B => n1120, CI => n1096, CO => n422, S 
                           => n423);
   U282 : ADFULD1 port map( A => n1006, B => n1146, CI => n1020, CO => n424, S 
                           => n425);
   U283 : ADFULD1 port map( A => n1174, B => n1036, CI => n431, CO => n426, S 
                           => n427);
   U284 : ADFULD1 port map( A => n1054, B => n984, CI => n994, CO => n428, S =>
                           n429);
   U285 : ADHALFDL port map( A => n1204, B => n943, CO => n430, S => n431);
   U286 : ADFULD1 port map( A => n454, B => n437, CI => n435, CO => n432, S => 
                           n433);
   U287 : ADFULD1 port map( A => n439, B => n441, CI => n456, CO => n434, S => 
                           n435);
   U288 : ADFULD1 port map( A => n443, B => n460, CI => n458, CO => n436, S => 
                           n437);
   U289 : ADFULD1 port map( A => n449, B => n445, CI => n447, CO => n438, S => 
                           n439);
   U290 : ADFULD1 port map( A => n464, B => n466, CI => n462, CO => n440, S => 
                           n441);
   U291 : ADFULD1 port map( A => n451, B => n1037, CI => n468, CO => n442, S =>
                           n443);
   U292 : ADFULD1 port map( A => n995, B => n1075, CI => n1007, CO => n444, S 
                           => n445);
   U293 : ADFULD1 port map( A => n1121, B => n1021, CI => n1097, CO => n446, S 
                           => n447);
   U294 : ADFULD1 port map( A => n1175, B => n1055, CI => n1147, CO => n448, S 
                           => n449);
   U295 : ADHALFDL port map( A => n470, B => n1205, CO => n450, S => n451);
   U296 : ADFULD1 port map( A => n474, B => n457, CI => n455, CO => n452, S => 
                           n453);
   U297 : ADFULD1 port map( A => n459, B => n461, CI => n476, CO => n454, S => 
                           n455);
   U298 : ADFULD1 port map( A => n480, B => n463, CI => n478, CO => n456, S => 
                           n457);
   U299 : ADFULD1 port map( A => n465, B => n469, CI => n467, CO => n458, S => 
                           n459);
   U300 : ADFULD1 port map( A => n482, B => n486, CI => n484, CO => n460, S => 
                           n461);
   U301 : ADFULD1 port map( A => n1098, B => n1122, CI => n488, CO => n462, S 
                           => n463);
   U302 : ADFULD1 port map( A => n1022, B => n1148, CI => n1056, CO => n464, S 
                           => n465);
   U303 : ADFULD1 port map( A => n1008, B => n1038, CI => n471, CO => n466, S 
                           => n467);
   U304 : ADFULD1 port map( A => n1076, B => n996, CI => n1176, CO => n468, S 
                           => n469);
   U305 : ADHALFDL port map( A => n1206, B => n944, CO => n470, S => n471);
   U306 : ADFULD1 port map( A => n492, B => n477, CI => n475, CO => n472, S => 
                           n473);
   U307 : ADFULD1 port map( A => n479, B => n481, CI => n494, CO => n474, S => 
                           n475);
   U308 : ADFULD1 port map( A => n498, B => n487, CI => n496, CO => n476, S => 
                           n477);
   U309 : ADFULD1 port map( A => n483, B => n500, CI => n485, CO => n478, S => 
                           n479);
   U310 : ADFULD1 port map( A => n504, B => n489, CI => n502, CO => n480, S => 
                           n481);
   U311 : ADFULD1 port map( A => n1057, B => n1149, CI => n1123, CO => n482, S 
                           => n483);
   U312 : ADFULD1 port map( A => n1177, B => n1099, CI => n1039, CO => n484, S 
                           => n485);
   U313 : ADFULD1 port map( A => n1009, B => n1077, CI => n1023, CO => n486, S 
                           => n487);
   U314 : ADHALFDL port map( A => n506, B => n1207, CO => n488, S => n489);
   U315 : ADFULD1 port map( A => n510, B => n495, CI => n493, CO => n490, S => 
                           n491);
   U316 : ADFULD1 port map( A => n497, B => n499, CI => n512, CO => n492, S => 
                           n493);
   U317 : ADFULD1 port map( A => n516, B => n503, CI => n514, CO => n494, S => 
                           n495);
   U318 : ADFULD1 port map( A => n505, B => n518, CI => n501, CO => n496, S => 
                           n497);
   U319 : ADFULD1 port map( A => n522, B => n1124, CI => n520, CO => n498, S =>
                           n499);
   U320 : ADFULD1 port map( A => n1040, B => n1150, CI => n1058, CO => n500, S 
                           => n501);
   U321 : ADFULD1 port map( A => n1178, B => n1100, CI => n507, CO => n502, S 
                           => n503);
   U322 : ADFULD1 port map( A => n1078, B => n1010, CI => n1024, CO => n504, S 
                           => n505);
   U323 : ADHALFDL port map( A => n1208, B => n945, CO => n506, S => n507);
   U324 : ADFULD1 port map( A => n526, B => n513, CI => n511, CO => n508, S => 
                           n509);
   U325 : ADFULD1 port map( A => n528, B => n530, CI => n515, CO => n510, S => 
                           n511);
   U326 : ADFULD1 port map( A => n521, B => n519, CI => n517, CO => n512, S => 
                           n513);
   U327 : ADFULD1 port map( A => n534, B => n536, CI => n532, CO => n514, S => 
                           n515);
   U328 : ADFULD1 port map( A => n1101, B => n1125, CI => n523, CO => n516, S 
                           => n517);
   U329 : ADFULD1 port map( A => n1025, B => n1041, CI => n1059, CO => n518, S 
                           => n519);
   U330 : ADFULD1 port map( A => n1179, B => n1079, CI => n1151, CO => n520, S 
                           => n521);
   U331 : ADHALFDL port map( A => n538, B => n1209, CO => n522, S => n523);
   U332 : ADFULD1 port map( A => n542, B => n529, CI => n527, CO => n524, S => 
                           n525);
   U333 : ADFULD1 port map( A => n544, B => n546, CI => n531, CO => n526, S => 
                           n527);
   U334 : ADFULD1 port map( A => n533, B => n537, CI => n535, CO => n528, S => 
                           n529);
   U335 : ADFULD1 port map( A => n550, B => n552, CI => n548, CO => n530, S => 
                           n531);
   U336 : ADFULD1 port map( A => n1080, B => n1152, CI => n1126, CO => n532, S 
                           => n533);
   U337 : ADFULD1 port map( A => n1042, B => n1060, CI => n539, CO => n534, S 
                           => n535);
   U338 : ADFULD1 port map( A => n1102, B => n1026, CI => n1180, CO => n536, S 
                           => n537);
   U339 : ADHALFDL port map( A => n1210, B => n946, CO => n538, S => n539);
   U340 : ADFULD1 port map( A => n556, B => n545, CI => n543, CO => n540, S => 
                           n541);
   U341 : ADFULD1 port map( A => n547, B => n551, CI => n558, CO => n542, S => 
                           n543);
   U342 : ADFULD1 port map( A => n560, B => n562, CI => n549, CO => n544, S => 
                           n545);
   U343 : ADFULD1 port map( A => n553, B => n1153, CI => n564, CO => n546, S =>
                           n547);
   U344 : ADFULD1 port map( A => n1181, B => n1081, CI => n1127, CO => n548, S 
                           => n549);
   U345 : ADFULD1 port map( A => n1043, B => n1103, CI => n1061, CO => n550, S 
                           => n551);
   U346 : ADHALFDL port map( A => n566, B => n1211, CO => n552, S => n553);
   U347 : ADFULD1 port map( A => n570, B => n559, CI => n557, CO => n554, S => 
                           n555);
   U348 : ADFULD1 port map( A => n561, B => n563, CI => n572, CO => n556, S => 
                           n557);
   U349 : ADFULD1 port map( A => n574, B => n576, CI => n565, CO => n558, S => 
                           n559);
   U350 : ADFULD1 port map( A => n1062, B => n1128, CI => n578, CO => n560, S 
                           => n561);
   U351 : ADFULD1 port map( A => n1154, B => n1082, CI => n567, CO => n562, S 
                           => n563);
   U352 : ADFULD1 port map( A => n1104, B => n1044, CI => n1182, CO => n564, S 
                           => n565);
   U353 : ADHALFDL port map( A => n1212, B => n947, CO => n566, S => n567);
   U354 : ADFULD1 port map( A => n582, B => n573, CI => n571, CO => n568, S => 
                           n569);
   U355 : ADFULD1 port map( A => n577, B => n575, CI => n584, CO => n570, S => 
                           n571);
   U356 : ADFULD1 port map( A => n588, B => n579, CI => n586, CO => n572, S => 
                           n573);
   U357 : ADFULD1 port map( A => n1063, B => n1129, CI => n1083, CO => n574, S 
                           => n575);
   U358 : ADFULD1 port map( A => n1183, B => n1105, CI => n1155, CO => n576, S 
                           => n577);
   U359 : ADHALFDL port map( A => n590, B => n1213, CO => n578, S => n579);
   U360 : ADFULD1 port map( A => n585, B => n594, CI => n583, CO => n580, S => 
                           n581);
   U361 : ADFULD1 port map( A => n587, B => n589, CI => n596, CO => n582, S => 
                           n583);
   U362 : ADFULD1 port map( A => n600, B => n1106, CI => n598, CO => n584, S =>
                           n585);
   U363 : ADFULD1 port map( A => n1084, B => n1156, CI => n591, CO => n586, S 
                           => n587);
   U364 : ADFULD1 port map( A => n1130, B => n1064, CI => n1184, CO => n588, S 
                           => n589);
   U365 : ADHALFDL port map( A => n1214, B => n948, CO => n590, S => n591);
   U366 : ADFULD1 port map( A => n604, B => n597, CI => n595, CO => n592, S => 
                           n593);
   U367 : ADFULD1 port map( A => n606, B => n608, CI => n599, CO => n594, S => 
                           n595);
   U368 : ADFULD1 port map( A => n1107, B => n1157, CI => n601, CO => n596, S 
                           => n597);
   U369 : ADFULD1 port map( A => n1085, B => n1131, CI => n1185, CO => n598, S 
                           => n599);
   U370 : ADHALFDL port map( A => n610, B => n1215, CO => n600, S => n601);
   U371 : ADFULD1 port map( A => n614, B => n607, CI => n605, CO => n602, S => 
                           n603);
   U372 : ADFULD1 port map( A => n616, B => n618, CI => n609, CO => n604, S => 
                           n605);
   U373 : ADFULD1 port map( A => n1108, B => n1158, CI => n611, CO => n606, S 
                           => n607);
   U374 : ADFULD1 port map( A => n1132, B => n1086, CI => n1186, CO => n608, S 
                           => n609);
   U375 : ADHALFDL port map( A => n1216, B => n949, CO => n610, S => n611);
   U376 : ADFULD1 port map( A => n617, B => n622, CI => n615, CO => n612, S => 
                           n613);
   U377 : ADFULD1 port map( A => n619, B => n1187, CI => n624, CO => n614, S =>
                           n615);
   U378 : ADFULD1 port map( A => n1109, B => n1133, CI => n1159, CO => n616, S 
                           => n617);
   U379 : ADHALFDL port map( A => n626, B => n1217, CO => n618, S => n619);
   U380 : ADFULD1 port map( A => n625, B => n630, CI => n623, CO => n620, S => 
                           n621);
   U381 : ADFULD1 port map( A => n627, B => n1160, CI => n632, CO => n622, S =>
                           n623);
   U382 : ADFULD1 port map( A => n1188, B => n1110, CI => n1134, CO => n624, S 
                           => n625);
   U383 : ADHALFDL port map( A => n1218, B => n950, CO => n626, S => n627);
   U384 : ADFULD1 port map( A => n636, B => n633, CI => n631, CO => n628, S => 
                           n629);
   U385 : ADFULD1 port map( A => n1135, B => n1189, CI => n1161, CO => n630, S 
                           => n631);
   U386 : ADHALFDL port map( A => n638, B => n1219, CO => n632, S => n633);
   U387 : ADFULD1 port map( A => n642, B => n639, CI => n637, CO => n634, S => 
                           n635);
   U388 : ADFULD1 port map( A => n1190, B => n1136, CI => n1162, CO => n636, S 
                           => n637);
   U389 : ADHALFDL port map( A => n1220, B => n951, CO => n638, S => n639);
   U390 : ADFULD1 port map( A => n1163, B => n1191, CI => n643, CO => n640, S 
                           => n641);
   U391 : ADHALFDL port map( A => n646, B => n1221, CO => n642, S => n643);
   U392 : ADFULD1 port map( A => n1192, B => n1164, CI => n647, CO => n644, S 
                           => n645);
   U393 : ADHALFDL port map( A => n1222, B => n952, CO => n646, S => n647);
   U394 : ADHALFDL port map( A => n650, B => n1223, CO => n648, S => n649);
   U395 : ADHALFDL port map( A => n1224, B => n953, CO => n650, S => n651);
   U397 : MUXB2DL port map( A0 => n104, A1 => n1426, SL => n652, Z => n955);
   U399 : MUXB2DL port map( A0 => n104, A1 => n1426, SL => n653, Z => n956);
   U402 : MUXB2DL port map( A0 => n99, A1 => n1425, SL => n654, Z => n957);
   U404 : MUXB2DL port map( A0 => n99, A1 => n1425, SL => n655, Z => n958);
   U406 : MUXB2DL port map( A0 => n99, A1 => n1425, SL => n656, Z => n959);
   U408 : MUXB2DL port map( A0 => n99, A1 => n1425, SL => n657, Z => n960);
   U411 : MUXB2DL port map( A0 => n94, A1 => n1422, SL => n658, Z => n961);
   U413 : MUXB2DL port map( A0 => n94, A1 => n1422, SL => n659, Z => n962);
   U415 : MUXB2DL port map( A0 => n94, A1 => n1422, SL => n660, Z => n963);
   U417 : MUXB2DL port map( A0 => n94, A1 => n1422, SL => n661, Z => n964);
   U419 : MUXB2DL port map( A0 => n94, A1 => n1422, SL => n662, Z => n965);
   U421 : MUXB2DL port map( A0 => n94, A1 => n1422, SL => n663, Z => n966);
   U424 : MUXB2DL port map( A0 => n89, A1 => n1420, SL => n664, Z => n967);
   U426 : MUXB2DL port map( A0 => n89, A1 => n1420, SL => n665, Z => n968);
   U428 : MUXB2DL port map( A0 => n89, A1 => n1420, SL => n666, Z => n969);
   U430 : MUXB2DL port map( A0 => n89, A1 => n1420, SL => n667, Z => n970);
   U432 : MUXB2DL port map( A0 => n89, A1 => n1420, SL => n668, Z => n971);
   U434 : MUXB2DL port map( A0 => n89, A1 => n1420, SL => n669, Z => n972);
   U436 : MUXB2DL port map( A0 => n89, A1 => n1420, SL => n670, Z => n973);
   U438 : MUXB2DL port map( A0 => n89, A1 => n1420, SL => n671, Z => n974);
   U441 : MUXB2DL port map( A0 => n84, A1 => n1418, SL => n672, Z => n975);
   U443 : MUXB2DL port map( A0 => n84, A1 => n1418, SL => n673, Z => n976);
   U445 : MUXB2DL port map( A0 => n84, A1 => n1418, SL => n674, Z => n977);
   U447 : MUXB2DL port map( A0 => n84, A1 => n1418, SL => n675, Z => n978);
   U449 : MUXB2DL port map( A0 => n84, A1 => n1418, SL => n676, Z => n979);
   U451 : MUXB2DL port map( A0 => n84, A1 => n1418, SL => n677, Z => n980);
   U453 : MUXB2DL port map( A0 => n84, A1 => n1418, SL => n678, Z => n981);
   U455 : MUXB2DL port map( A0 => n84, A1 => n1418, SL => n679, Z => n982);
   U457 : MUXB2DL port map( A0 => n84, A1 => n1418, SL => n680, Z => n983);
   U459 : MUXB2DL port map( A0 => n84, A1 => n1418, SL => n681, Z => n984);
   U462 : MUXB2DL port map( A0 => n80, A1 => n1416, SL => n682, Z => n985);
   U464 : MUXB2DL port map( A0 => n80, A1 => n1416, SL => n683, Z => n986);
   U466 : MUXB2DL port map( A0 => n80, A1 => n1416, SL => n684, Z => n987);
   U468 : MUXB2DL port map( A0 => n80, A1 => n1416, SL => n685, Z => n988);
   U470 : MUXB2DL port map( A0 => n80, A1 => n1416, SL => n686, Z => n989);
   U472 : MUXB2DL port map( A0 => n80, A1 => n1416, SL => n687, Z => n990);
   U474 : MUXB2DL port map( A0 => n80, A1 => n1416, SL => n688, Z => n991);
   U476 : MUXB2DL port map( A0 => n80, A1 => n1416, SL => n689, Z => n992);
   U478 : MUXB2DL port map( A0 => n80, A1 => n1416, SL => n690, Z => n993);
   U480 : MUXB2DL port map( A0 => n80, A1 => n1416, SL => n691, Z => n994);
   U482 : MUXB2DL port map( A0 => n80, A1 => n1416, SL => n692, Z => n995);
   U484 : MUXB2DL port map( A0 => n80, A1 => n1416, SL => n693, Z => n996);
   U487 : MUXB2DL port map( A0 => n73, A1 => n1414, SL => n694, Z => n997);
   U489 : MUXB2DL port map( A0 => n73, A1 => n1414, SL => n695, Z => n998);
   U491 : MUXB2DL port map( A0 => n73, A1 => n1414, SL => n696, Z => n999);
   U493 : MUXB2DL port map( A0 => n73, A1 => n1414, SL => n697, Z => n1000);
   U495 : MUXB2DL port map( A0 => n73, A1 => n1414, SL => n698, Z => n1001);
   U497 : MUXB2DL port map( A0 => n73, A1 => n1414, SL => n699, Z => n1002);
   U499 : MUXB2DL port map( A0 => n73, A1 => n1414, SL => n700, Z => n1003);
   U501 : MUXB2DL port map( A0 => n73, A1 => n1414, SL => n701, Z => n1004);
   U503 : MUXB2DL port map( A0 => n73, A1 => n1414, SL => n702, Z => n1005);
   U505 : MUXB2DL port map( A0 => n73, A1 => n1414, SL => n703, Z => n1006);
   U507 : MUXB2DL port map( A0 => n73, A1 => n1414, SL => n704, Z => n1007);
   U509 : MUXB2DL port map( A0 => n73, A1 => n1414, SL => n705, Z => n1008);
   U511 : MUXB2DL port map( A0 => n73, A1 => n1414, SL => n706, Z => n1009);
   U513 : MUXB2DL port map( A0 => n73, A1 => n1414, SL => n707, Z => n1010);
   U516 : MUXB2DL port map( A0 => n66, A1 => n1412, SL => n708, Z => n1011);
   U518 : MUXB2DL port map( A0 => n66, A1 => n1412, SL => n709, Z => n1012);
   U520 : MUXB2DL port map( A0 => n66, A1 => n1412, SL => n710, Z => n1013);
   U522 : MUXB2DL port map( A0 => n66, A1 => n1412, SL => n711, Z => n1014);
   U524 : MUXB2DL port map( A0 => n66, A1 => n1412, SL => n712, Z => n1015);
   U526 : MUXB2DL port map( A0 => n66, A1 => n1412, SL => n713, Z => n1016);
   U528 : MUXB2DL port map( A0 => n66, A1 => n1412, SL => n714, Z => n1017);
   U530 : MUXB2DL port map( A0 => n66, A1 => n1412, SL => n715, Z => n1018);
   U532 : MUXB2DL port map( A0 => n66, A1 => n1412, SL => n716, Z => n1019);
   U534 : MUXB2DL port map( A0 => n66, A1 => n1412, SL => n717, Z => n1020);
   U536 : MUXB2DL port map( A0 => n66, A1 => n1412, SL => n718, Z => n1021);
   U538 : MUXB2DL port map( A0 => n66, A1 => n1412, SL => n719, Z => n1022);
   U540 : MUXB2DL port map( A0 => n66, A1 => n1412, SL => n720, Z => n1023);
   U542 : MUXB2DL port map( A0 => n66, A1 => n1412, SL => n721, Z => n1024);
   U544 : MUXB2DL port map( A0 => n66, A1 => n1412, SL => n722, Z => n1025);
   U546 : MUXB2DL port map( A0 => n66, A1 => n1412, SL => n723, Z => n1026);
   U549 : MUXB2DL port map( A0 => n58, A1 => n1410, SL => n724, Z => n1027);
   U551 : MUXB2DL port map( A0 => n58, A1 => n1410, SL => n725, Z => n1028);
   U553 : MUXB2DL port map( A0 => n58, A1 => n1410, SL => n726, Z => n1029);
   U555 : MUXB2DL port map( A0 => n58, A1 => n1410, SL => n727, Z => n1030);
   U557 : MUXB2DL port map( A0 => n58, A1 => n1410, SL => n728, Z => n1031);
   U559 : MUXB2DL port map( A0 => n58, A1 => n1410, SL => n729, Z => n1032);
   U561 : MUXB2DL port map( A0 => n58, A1 => n1410, SL => n730, Z => n1033);
   U563 : MUXB2DL port map( A0 => n58, A1 => n1410, SL => n731, Z => n1034);
   U565 : MUXB2DL port map( A0 => n58, A1 => n1410, SL => n732, Z => n1035);
   U567 : MUXB2DL port map( A0 => n58, A1 => n1410, SL => n733, Z => n1036);
   U569 : MUXB2DL port map( A0 => n58, A1 => n1410, SL => n734, Z => n1037);
   U571 : MUXB2DL port map( A0 => n58, A1 => n1410, SL => n735, Z => n1038);
   U573 : MUXB2DL port map( A0 => n58, A1 => n1410, SL => n736, Z => n1039);
   U575 : MUXB2DL port map( A0 => n58, A1 => n1410, SL => n737, Z => n1040);
   U577 : MUXB2DL port map( A0 => n58, A1 => n1410, SL => n738, Z => n1041);
   U579 : MUXB2DL port map( A0 => n58, A1 => n1410, SL => n739, Z => n1042);
   U581 : MUXB2DL port map( A0 => n58, A1 => n1410, SL => n740, Z => n1043);
   U583 : MUXB2DL port map( A0 => n58, A1 => n1410, SL => n741, Z => n1044);
   U586 : MUXB2DL port map( A0 => n50, A1 => n1408, SL => n742, Z => n1045);
   U588 : MUXB2DL port map( A0 => n50, A1 => n1408, SL => n743, Z => n1046);
   U590 : MUXB2DL port map( A0 => n50, A1 => n1408, SL => n744, Z => n1047);
   U592 : MUXB2DL port map( A0 => n50, A1 => n1408, SL => n745, Z => n1048);
   U594 : MUXB2DL port map( A0 => n50, A1 => n1408, SL => n746, Z => n1049);
   U596 : MUXB2DL port map( A0 => n50, A1 => n1408, SL => n747, Z => n1050);
   U598 : MUXB2DL port map( A0 => n50, A1 => n1408, SL => n748, Z => n1051);
   U600 : MUXB2DL port map( A0 => n50, A1 => n1408, SL => n749, Z => n1052);
   U602 : MUXB2DL port map( A0 => n50, A1 => n1408, SL => n750, Z => n1053);
   U604 : MUXB2DL port map( A0 => n50, A1 => n1408, SL => n751, Z => n1054);
   U606 : MUXB2DL port map( A0 => n50, A1 => n1408, SL => n752, Z => n1055);
   U608 : MUXB2DL port map( A0 => n50, A1 => n1408, SL => n753, Z => n1056);
   U610 : MUXB2DL port map( A0 => n50, A1 => n1408, SL => n754, Z => n1057);
   U612 : MUXB2DL port map( A0 => n50, A1 => n1408, SL => n755, Z => n1058);
   U614 : MUXB2DL port map( A0 => n50, A1 => n1408, SL => n756, Z => n1059);
   U616 : MUXB2DL port map( A0 => n50, A1 => n1408, SL => n757, Z => n1060);
   U618 : MUXB2DL port map( A0 => n50, A1 => n1408, SL => n758, Z => n1061);
   U620 : MUXB2DL port map( A0 => n50, A1 => n1408, SL => n759, Z => n1062);
   U622 : MUXB2DL port map( A0 => n50, A1 => n1408, SL => n760, Z => n1063);
   U624 : MUXB2DL port map( A0 => n50, A1 => n1408, SL => n761, Z => n1064);
   U627 : MUXB2DL port map( A0 => n42, A1 => n1406, SL => n762, Z => n1065);
   U629 : MUXB2DL port map( A0 => n42, A1 => n1406, SL => n763, Z => n1066);
   U631 : MUXB2DL port map( A0 => n42, A1 => n1406, SL => n764, Z => n1067);
   U633 : MUXB2DL port map( A0 => n42, A1 => n1406, SL => n765, Z => n1068);
   U635 : MUXB2DL port map( A0 => n42, A1 => n1406, SL => n766, Z => n1069);
   U637 : MUXB2DL port map( A0 => n42, A1 => n1406, SL => n767, Z => n1070);
   U639 : MUXB2DL port map( A0 => n42, A1 => n1406, SL => n768, Z => n1071);
   U641 : MUXB2DL port map( A0 => n42, A1 => n1406, SL => n769, Z => n1072);
   U643 : MUXB2DL port map( A0 => n42, A1 => n1406, SL => n770, Z => n1073);
   U645 : MUXB2DL port map( A0 => n42, A1 => n1406, SL => n771, Z => n1074);
   U647 : MUXB2DL port map( A0 => n42, A1 => n1406, SL => n772, Z => n1075);
   U649 : MUXB2DL port map( A0 => n42, A1 => n1406, SL => n773, Z => n1076);
   U651 : MUXB2DL port map( A0 => n42, A1 => n1406, SL => n774, Z => n1077);
   U653 : MUXB2DL port map( A0 => n42, A1 => n1406, SL => n775, Z => n1078);
   U655 : MUXB2DL port map( A0 => n42, A1 => n1406, SL => n776, Z => n1079);
   U657 : MUXB2DL port map( A0 => n42, A1 => n1406, SL => n777, Z => n1080);
   U659 : MUXB2DL port map( A0 => n42, A1 => n1406, SL => n778, Z => n1081);
   U661 : MUXB2DL port map( A0 => n42, A1 => n1406, SL => n779, Z => n1082);
   U663 : MUXB2DL port map( A0 => n42, A1 => n1406, SL => n780, Z => n1083);
   U665 : MUXB2DL port map( A0 => n42, A1 => n1406, SL => n781, Z => n1084);
   U667 : MUXB2DL port map( A0 => n42, A1 => n1406, SL => n782, Z => n1085);
   U669 : MUXB2DL port map( A0 => n42, A1 => n1406, SL => n783, Z => n1086);
   U672 : MUXB2DL port map( A0 => n1382, A1 => n1404, SL => n784, Z => n1087);
   U674 : MUXB2DL port map( A0 => n1382, A1 => n1404, SL => n785, Z => n1088);
   U676 : MUXB2DL port map( A0 => n1382, A1 => n1404, SL => n786, Z => n1089);
   U678 : MUXB2DL port map( A0 => n1382, A1 => n1404, SL => n787, Z => n1090);
   U680 : MUXB2DL port map( A0 => n1382, A1 => n1404, SL => n788, Z => n1091);
   U682 : MUXB2DL port map( A0 => n1382, A1 => n1404, SL => n789, Z => n1092);
   U684 : MUXB2DL port map( A0 => n1382, A1 => n1404, SL => n790, Z => n1093);
   U686 : MUXB2DL port map( A0 => n1382, A1 => n1404, SL => n791, Z => n1094);
   U688 : MUXB2DL port map( A0 => n1382, A1 => n1404, SL => n792, Z => n1095);
   U690 : MUXB2DL port map( A0 => n1382, A1 => n1404, SL => n793, Z => n1096);
   U692 : MUXB2DL port map( A0 => n1382, A1 => n1404, SL => n794, Z => n1097);
   U694 : MUXB2DL port map( A0 => n1382, A1 => n1404, SL => n795, Z => n1098);
   U696 : MUXB2DL port map( A0 => n1382, A1 => n1404, SL => n796, Z => n1099);
   U698 : MUXB2DL port map( A0 => n1382, A1 => n1404, SL => n797, Z => n1100);
   U700 : MUXB2DL port map( A0 => n1382, A1 => n1404, SL => n798, Z => n1101);
   U702 : MUXB2DL port map( A0 => n1382, A1 => n1404, SL => n799, Z => n1102);
   U704 : MUXB2DL port map( A0 => n1382, A1 => n1404, SL => n800, Z => n1103);
   U706 : MUXB2DL port map( A0 => n1382, A1 => n1404, SL => n801, Z => n1104);
   U708 : MUXB2DL port map( A0 => n1382, A1 => n1404, SL => n802, Z => n1105);
   U710 : MUXB2DL port map( A0 => n1382, A1 => n1404, SL => n803, Z => n1106);
   U712 : MUXB2DL port map( A0 => n1382, A1 => n1404, SL => n804, Z => n1107);
   U714 : MUXB2DL port map( A0 => n1382, A1 => n1404, SL => n805, Z => n1108);
   U716 : MUXB2DL port map( A0 => n1382, A1 => n1404, SL => n806, Z => n1109);
   U718 : MUXB2DL port map( A0 => n1382, A1 => n1404, SL => n807, Z => n1110);
   U721 : MUXB2DL port map( A0 => n1381, A1 => n1402, SL => n808, Z => n1111);
   U723 : MUXB2DL port map( A0 => n1381, A1 => n1402, SL => n809, Z => n1112);
   U725 : MUXB2DL port map( A0 => n1381, A1 => n1402, SL => n810, Z => n1113);
   U727 : MUXB2DL port map( A0 => n1381, A1 => n1402, SL => n811, Z => n1114);
   U729 : MUXB2DL port map( A0 => n1381, A1 => n1402, SL => n812, Z => n1115);
   U731 : MUXB2DL port map( A0 => n1381, A1 => n1402, SL => n813, Z => n1116);
   U733 : MUXB2DL port map( A0 => n1381, A1 => n1402, SL => n814, Z => n1117);
   U735 : MUXB2DL port map( A0 => n1381, A1 => n1402, SL => n815, Z => n1118);
   U737 : MUXB2DL port map( A0 => n1381, A1 => n1402, SL => n816, Z => n1119);
   U739 : MUXB2DL port map( A0 => n1381, A1 => n1402, SL => n817, Z => n1120);
   U741 : MUXB2DL port map( A0 => n1381, A1 => n1402, SL => n818, Z => n1121);
   U743 : MUXB2DL port map( A0 => n1381, A1 => n1402, SL => n819, Z => n1122);
   U745 : MUXB2DL port map( A0 => n1381, A1 => n1402, SL => n820, Z => n1123);
   U747 : MUXB2DL port map( A0 => n1381, A1 => n1402, SL => n821, Z => n1124);
   U749 : MUXB2DL port map( A0 => n1381, A1 => n1402, SL => n822, Z => n1125);
   U751 : MUXB2DL port map( A0 => n1381, A1 => n1402, SL => n823, Z => n1126);
   U753 : MUXB2DL port map( A0 => n1381, A1 => n1402, SL => n824, Z => n1127);
   U755 : MUXB2DL port map( A0 => n1381, A1 => n1402, SL => n825, Z => n1128);
   U757 : MUXB2DL port map( A0 => n1381, A1 => n1402, SL => n826, Z => n1129);
   U759 : MUXB2DL port map( A0 => n1381, A1 => n1402, SL => n827, Z => n1130);
   U761 : MUXB2DL port map( A0 => n1381, A1 => n1402, SL => n828, Z => n1131);
   U763 : MUXB2DL port map( A0 => n1381, A1 => n1402, SL => n829, Z => n1132);
   U765 : MUXB2DL port map( A0 => n1381, A1 => n1402, SL => n830, Z => n1133);
   U767 : MUXB2DL port map( A0 => n1381, A1 => n1402, SL => n831, Z => n1134);
   U769 : MUXB2DL port map( A0 => n1381, A1 => n1402, SL => n832, Z => n1135);
   U771 : MUXB2DL port map( A0 => n1381, A1 => n1402, SL => n833, Z => n1136);
   U774 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n834, Z => n1137);
   U776 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n835, Z => n1138);
   U778 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n836, Z => n1139);
   U780 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n837, Z => n1140);
   U782 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n838, Z => n1141);
   U784 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n839, Z => n1142);
   U786 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n840, Z => n1143);
   U788 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n841, Z => n1144);
   U790 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n842, Z => n1145);
   U792 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n843, Z => n1146);
   U794 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n844, Z => n1147);
   U796 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n845, Z => n1148);
   U798 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n846, Z => n1149);
   U800 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n847, Z => n1150);
   U802 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n848, Z => n1151);
   U804 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n849, Z => n1152);
   U806 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n850, Z => n1153);
   U808 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n851, Z => n1154);
   U810 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n852, Z => n1155);
   U812 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n853, Z => n1156);
   U814 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n854, Z => n1157);
   U816 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n855, Z => n1158);
   U818 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n856, Z => n1159);
   U820 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n857, Z => n1160);
   U822 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n858, Z => n1161);
   U824 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n859, Z => n1162);
   U826 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n860, Z => n1163);
   U828 : MUXB2DL port map( A0 => n1380, A1 => n1400, SL => n861, Z => n1164);
   U831 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n862, Z => n1165);
   U833 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n863, Z => n1166);
   U835 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n864, Z => n1167);
   U837 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n865, Z => n1168);
   U839 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n866, Z => n1169);
   U841 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n867, Z => n1170);
   U843 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n868, Z => n1171);
   U845 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n869, Z => n1172);
   U847 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n870, Z => n1173);
   U849 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n871, Z => n1174);
   U851 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n872, Z => n1175);
   U853 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n873, Z => n1176);
   U855 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n874, Z => n1177);
   U857 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n875, Z => n1178);
   U859 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n876, Z => n1179);
   U861 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n877, Z => n1180);
   U863 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n878, Z => n1181);
   U865 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n879, Z => n1182);
   U867 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n880, Z => n1183);
   U869 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n881, Z => n1184);
   U871 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n882, Z => n1185);
   U873 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n883, Z => n1186);
   U875 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n884, Z => n1187);
   U877 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n885, Z => n1188);
   U879 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n886, Z => n1189);
   U881 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n887, Z => n1190);
   U883 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n888, Z => n1191);
   U885 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n889, Z => n1192);
   U887 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n890, Z => n1193);
   U889 : MUXB2DL port map( A0 => n1379, A1 => n1399, SL => n891, Z => n1194);
   U892 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n892, Z => n1195);
   U894 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n893, Z => n1196);
   U896 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n894, Z => n1197);
   U898 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n895, Z => n1198);
   U900 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n896, Z => n1199);
   U902 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n897, Z => n1200);
   U904 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n898, Z => n1201);
   U906 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n899, Z => n1202);
   U908 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n900, Z => n1203);
   U910 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n901, Z => n1204);
   U912 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n902, Z => n1205);
   U914 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n903, Z => n1206);
   U916 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n904, Z => n1207);
   U918 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n905, Z => n1208);
   U920 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n906, Z => n1209);
   U922 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n907, Z => n1210);
   U924 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n908, Z => n1211);
   U926 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n909, Z => n1212);
   U928 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n910, Z => n1213);
   U930 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n911, Z => n1214);
   U932 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n912, Z => n1215);
   U934 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n913, Z => n1216);
   U936 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n914, Z => n1217);
   U938 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n915, Z => n1218);
   U940 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n916, Z => n1219);
   U942 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n917, Z => n1220);
   U944 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n918, Z => n1221);
   U946 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n919, Z => n1222);
   U948 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n920, Z => n1223);
   U950 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n921, Z => n1224);
   U952 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n922, Z => n1225);
   U954 : MUXB2DL port map( A0 => n1378, A1 => n1398, SL => n923, Z => n1226);
   U1021 : EXOR2D1 port map( A1 => a(4), A2 => a(3), Z => n1375);
   U1022 : EXOR2D1 port map( A1 => a(6), A2 => a(5), Z => n1376);
   U1023 : EXOR2D1 port map( A1 => a(8), A2 => a(7), Z => n1377);
   U1024 : NAN2D1 port map( A1 => a(0), A2 => n1398, Z => n1378);
   U1025 : OAI21D1 port map( A1 => a(2), A2 => a(1), B => n1401, Z => n1379);
   U1026 : OAI21D1 port map( A1 => a(4), A2 => a(3), B => n1403, Z => n1380);
   U1027 : OAI21D1 port map( A1 => a(6), A2 => a(5), B => n1405, Z => n1381);
   U1028 : OAI21D1 port map( A1 => a(8), A2 => a(7), B => n1407, Z => n1382);
   U1029 : INVD1 port map( A => n1383, Z => n1384);
   U1030 : INVD1 port map( A => n1393, Z => n1392);
   U1031 : INVD1 port map( A => n1395, Z => n1394);
   U1032 : INVD1 port map( A => n1397, Z => n1396);
   U1033 : INVD1 port map( A => n1391, Z => n1389);
   U1034 : INVD1 port map( A => n1391, Z => n1390);
   U1035 : INVD1 port map( A => n953, Z => n1399);
   U1036 : INVD1 port map( A => n1386, Z => n1385);
   U1037 : INVD1 port map( A => n1388, Z => n1387);
   U1038 : INVD1 port map( A => n952, Z => n1400);
   U1039 : INVD1 port map( A => n951, Z => n1402);
   U1040 : INVD1 port map( A => n950, Z => n1404);
   U1041 : INVD1 port map( A => n949, Z => n1406);
   U1042 : INVD1 port map( A => n948, Z => n1408);
   U1043 : INVD1 port map( A => n947, Z => n1410);
   U1044 : INVD1 port map( A => n946, Z => n1412);
   U1045 : INVD1 port map( A => n945, Z => n1414);
   U1046 : INVD1 port map( A => n944, Z => n1416);
   U1047 : INVD1 port map( A => n943, Z => n1418);
   U1048 : INVD1 port map( A => n942, Z => n1420);
   U1049 : INVD1 port map( A => n941, Z => n1422);
   U1050 : INVD1 port map( A => n940, Z => n1425);
   U1051 : INVD1 port map( A => n939, Z => n1426);
   U1052 : INVD1 port map( A => a(1), Z => n1398);
   U1053 : EXNOR2D1 port map( A1 => a(2), A2 => a(1), Z => n1383);
   U1054 : INVD1 port map( A => b(2), Z => n1393);
   U1055 : INVD1 port map( A => b(1), Z => n1395);
   U1056 : INVD1 port map( A => b(0), Z => n1397);
   U1057 : INVD1 port map( A => b(3), Z => n1391);
   U1058 : INVD1 port map( A => b(4), Z => n1388);
   U1059 : INVD1 port map( A => a(3), Z => n1401);
   U1060 : INVD1 port map( A => a(5), Z => n1403);
   U1061 : INVD1 port map( A => b(5), Z => n1386);
   U1062 : INVD1 port map( A => a(7), Z => n1405);
   U1063 : INVD1 port map( A => a(9), Z => n1407);
   U1064 : EXOR2D1 port map( A1 => a(10), A2 => a(9), Z => n1447);
   U1065 : INVD1 port map( A => a(11), Z => n1409);
   U1066 : OAI21D1 port map( A1 => a(9), A2 => a(10), B => n1409, Z => n42);
   U1067 : EXOR2D1 port map( A1 => a(12), A2 => a(11), Z => n1448);
   U1068 : INVD1 port map( A => a(13), Z => n1411);
   U1069 : OAI21D1 port map( A1 => a(12), A2 => a(11), B => n1411, Z => n50);
   U1070 : EXOR2D1 port map( A1 => a(14), A2 => a(13), Z => n1449);
   U1071 : INVD1 port map( A => a(15), Z => n1413);
   U1072 : OAI21D1 port map( A1 => a(14), A2 => a(13), B => n1413, Z => n58);
   U1073 : EXOR2D1 port map( A1 => a(16), A2 => a(15), Z => n1450);
   U1074 : INVD1 port map( A => a(17), Z => n1415);
   U1075 : OAI21D1 port map( A1 => a(16), A2 => a(15), B => n1415, Z => n66);
   U1076 : EXOR2D1 port map( A1 => a(18), A2 => a(17), Z => n1451);
   U1077 : INVD1 port map( A => a(19), Z => n1417);
   U1078 : OAI21D1 port map( A1 => a(18), A2 => a(17), B => n1417, Z => n73);
   U1079 : EXOR2D1 port map( A1 => a(20), A2 => a(19), Z => n1452);
   U1080 : INVD1 port map( A => a(21), Z => n1419);
   U1081 : OAI21D1 port map( A1 => a(20), A2 => a(19), B => n1419, Z => n80);
   U1082 : EXOR2D1 port map( A1 => a(22), A2 => a(21), Z => n1453);
   U1083 : INVD1 port map( A => a(23), Z => n1421);
   U1084 : OAI21D1 port map( A1 => a(22), A2 => a(21), B => n1421, Z => n84);
   U1085 : INVD1 port map( A => a(25), Z => n1423);
   U1086 : INVD1 port map( A => a(27), Z => n1424);
   U1087 : INVD1 port map( A => a(29), Z => n1427);
   U1088 : MUXB2DL port map( A0 => b(29), A1 => b(28), SL => n1383, Z => n862);
   U1089 : INVD1 port map( A => a(31), Z => n1428);
   U1090 : EXOR3D1 port map( A1 => n1429, A2 => n1430, A3 => n1431, Z => 
                           product(31));
   U1091 : EXOR3D1 port map( A1 => n208, A2 => n206, A3 => n1432, Z => n1431);
   U1092 : EXOR2D1 port map( A1 => n214, A2 => n212, Z => n1432);
   U1093 : EXOR2D1 port map( A1 => n202, A2 => n156, Z => n1430);
   U1094 : EXOR3D1 port map( A1 => n1433, A2 => n1434, A3 => n1435, Z => n1429)
                           ;
   U1095 : EXOR3D1 port map( A1 => n957, A2 => n955, A3 => n1436, Z => n1435);
   U1096 : EXNOR2D1 port map( A1 => n997, A2 => n975, Z => n1436);
   U1097 : EXOR3D1 port map( A1 => n1437, A2 => n204, A3 => n1438, Z => n1434);
   U1098 : EXOR3D1 port map( A1 => n1087, A2 => n1065, A3 => n1439, Z => n1438)
                           ;
   U1099 : EXNOR2D1 port map( A1 => n210, A2 => n1111, Z => n1439);
   U1100 : EXOR3D1 port map( A1 => n961, A2 => n218, A3 => n1440, Z => n1437);
   U1101 : EXOR2D1 port map( A1 => n985, A2 => n967, Z => n1440);
   U1102 : EXOR3D1 port map( A1 => n1441, A2 => n1442, A3 => n1443, Z => n1433)
                           ;
   U1103 : EXOR3D1 port map( A1 => n1027, A2 => n1011, A3 => n1444, Z => n1443)
                           ;
   U1104 : EXOR3D1 port map( A1 => n1165, A2 => n1137, A3 => n1045, Z => n1444)
                           ;
   U1105 : EXOR3D1 port map( A1 => n216, A2 => n1195, A3 => n1445, Z => n1442);
   U1106 : EXOR2D1 port map( A1 => n222, A2 => n220, Z => n1445);
   U1107 : EXOR3D1 port map( A1 => n226, A2 => n224, A3 => n1446, Z => n1441);
   U1108 : EXOR2D1 port map( A1 => n230, A2 => n228, Z => n1446);
   U1109 : OAI21D1 port map( A1 => a(28), A2 => a(27), B => n1427, Z => n99);
   U1110 : AOI21D1 port map( A1 => a(25), A2 => a(26), B => n1424, Z => n941);
   U1111 : OAI21D1 port map( A1 => a(26), A2 => a(25), B => n1424, Z => n94);
   U1112 : NAN2D1 port map( A1 => n1396, A2 => a(0), Z => n923);
   U1113 : MUXB2DL port map( A0 => n1396, A1 => b(1), SL => a(0), Z => n922);
   U1114 : MUXB2DL port map( A0 => n1394, A1 => n1392, SL => a(0), Z => n921);
   U1115 : MUXB2DL port map( A0 => n1392, A1 => n1390, SL => a(0), Z => n920);
   U1116 : MUXB2DL port map( A0 => n1389, A1 => b(4), SL => a(0), Z => n919);
   U1117 : MUXB2DL port map( A0 => n1387, A1 => n1385, SL => a(0), Z => n918);
   U1118 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => a(0), Z => n917);
   U1119 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => a(0), Z => n916);
   U1120 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => a(0), Z => n915);
   U1121 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => a(0), Z => n914);
   U1122 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => a(0), Z => n913);
   U1123 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => a(0), Z => n912);
   U1124 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => a(0), Z => n911);
   U1125 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => a(0), Z => n910);
   U1126 : AOI21D1 port map( A1 => a(23), A2 => a(24), B => n1423, Z => n942);
   U1127 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => a(0), Z => n909);
   U1128 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => a(0), Z => n908);
   U1129 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => a(0), Z => n907);
   U1130 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => a(0), Z => n906);
   U1131 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => a(0), Z => n905);
   U1132 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => a(0), Z => n904);
   U1133 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => a(0), Z => n903);
   U1134 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => a(0), Z => n902);
   U1135 : MUXB2DL port map( A0 => b(21), A1 => b(22), SL => a(0), Z => n901);
   U1136 : MUXB2DL port map( A0 => b(22), A1 => b(23), SL => a(0), Z => n900);
   U1137 : MUXB2DL port map( A0 => b(23), A1 => b(24), SL => a(0), Z => n899);
   U1138 : MUXB2DL port map( A0 => b(24), A1 => b(25), SL => a(0), Z => n898);
   U1139 : MUXB2DL port map( A0 => b(25), A1 => b(26), SL => a(0), Z => n897);
   U1140 : MUXB2DL port map( A0 => b(26), A1 => b(27), SL => a(0), Z => n896);
   U1141 : MUXB2DL port map( A0 => b(27), A1 => b(28), SL => a(0), Z => n895);
   U1142 : MUXB2DL port map( A0 => b(28), A1 => b(29), SL => a(0), Z => n894);
   U1143 : MUXB2DL port map( A0 => b(29), A1 => b(30), SL => a(0), Z => n893);
   U1144 : MUXB2DL port map( A0 => b(30), A1 => b(31), SL => a(0), Z => n892);
   U1145 : NAN2D1 port map( A1 => n1396, A2 => n1384, Z => n891);
   U1146 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1384, Z => n890);
   U1147 : OAI21D1 port map( A1 => a(24), A2 => a(23), B => n1423, Z => n89);
   U1148 : MUXB2DL port map( A0 => n1394, A1 => n1392, SL => n1384, Z => n889);
   U1149 : MUXB2DL port map( A0 => b(2), A1 => n1390, SL => n1384, Z => n888);
   U1150 : MUXB2DL port map( A0 => n1389, A1 => n1387, SL => n1384, Z => n887);
   U1151 : MUXB2DL port map( A0 => n1387, A1 => n1385, SL => n1384, Z => n886);
   U1152 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1384, Z => n885);
   U1153 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1384, Z => n884);
   U1154 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1384, Z => n883);
   U1155 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1384, Z => n882);
   U1156 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1384, Z => n881);
   U1157 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1384, Z => n880);
   U1158 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1384, Z => n879);
   U1159 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1384, Z => n878);
   U1160 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1384, Z => n877);
   U1161 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1384, Z => n876);
   U1162 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1384, Z => n875);
   U1163 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1384, Z => n874);
   U1164 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1384, Z => n873);
   U1165 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1384, Z => n872);
   U1166 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => n1384, Z => n871);
   U1167 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => n1384, Z => n870);
   U1168 : MUXB2DL port map( A0 => b(21), A1 => b(22), SL => n1384, Z => n869);
   U1169 : MUXB2DL port map( A0 => b(22), A1 => b(23), SL => n1384, Z => n868);
   U1170 : MUXB2DL port map( A0 => b(23), A1 => b(24), SL => n1384, Z => n867);
   U1171 : MUXB2DL port map( A0 => b(24), A1 => b(25), SL => n1384, Z => n866);
   U1172 : MUXB2DL port map( A0 => b(25), A1 => b(26), SL => n1384, Z => n865);
   U1173 : MUXB2DL port map( A0 => b(26), A1 => b(27), SL => n1384, Z => n864);
   U1174 : MUXB2DL port map( A0 => b(27), A1 => b(28), SL => n1384, Z => n863);
   U1175 : NAN2D1 port map( A1 => n1396, A2 => n1375, Z => n861);
   U1176 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1375, Z => n860);
   U1177 : AOI21D1 port map( A1 => a(21), A2 => a(22), B => n1421, Z => n943);
   U1178 : MUXB2DL port map( A0 => n1394, A1 => n1392, SL => n1375, Z => n859);
   U1179 : MUXB2DL port map( A0 => b(2), A1 => n1390, SL => n1375, Z => n858);
   U1180 : MUXB2DL port map( A0 => n1389, A1 => n1387, SL => n1375, Z => n857);
   U1181 : MUXB2DL port map( A0 => n1387, A1 => n1385, SL => n1375, Z => n856);
   U1182 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1375, Z => n855);
   U1183 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1375, Z => n854);
   U1184 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1375, Z => n853);
   U1185 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1375, Z => n852);
   U1186 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1375, Z => n851);
   U1187 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1375, Z => n850);
   U1188 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1375, Z => n849);
   U1189 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1375, Z => n848);
   U1190 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1375, Z => n847);
   U1191 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1375, Z => n846);
   U1192 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1375, Z => n845);
   U1193 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1375, Z => n844);
   U1194 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1375, Z => n843);
   U1195 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1375, Z => n842);
   U1196 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => n1375, Z => n841);
   U1197 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => n1375, Z => n840);
   U1198 : MUXB2DL port map( A0 => b(21), A1 => b(22), SL => n1375, Z => n839);
   U1199 : MUXB2DL port map( A0 => b(22), A1 => b(23), SL => n1375, Z => n838);
   U1200 : MUXB2DL port map( A0 => b(23), A1 => b(24), SL => n1375, Z => n837);
   U1201 : MUXB2DL port map( A0 => b(24), A1 => b(25), SL => n1375, Z => n836);
   U1202 : MUXB2DL port map( A0 => b(25), A1 => b(26), SL => n1375, Z => n835);
   U1203 : MUXB2DL port map( A0 => b(26), A1 => b(27), SL => n1375, Z => n834);
   U1204 : NAN2D1 port map( A1 => n1396, A2 => n1376, Z => n833);
   U1205 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1376, Z => n832);
   U1206 : MUXB2DL port map( A0 => n1394, A1 => n1392, SL => n1376, Z => n831);
   U1207 : MUXB2DL port map( A0 => n1392, A1 => n1390, SL => n1376, Z => n830);
   U1208 : MUXB2DL port map( A0 => n1389, A1 => n1387, SL => n1376, Z => n829);
   U1209 : MUXB2DL port map( A0 => n1387, A1 => n1385, SL => n1376, Z => n828);
   U1210 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1376, Z => n827);
   U1211 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1376, Z => n826);
   U1212 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1376, Z => n825);
   U1213 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1376, Z => n824);
   U1214 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1376, Z => n823);
   U1215 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1376, Z => n822);
   U1216 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1376, Z => n821);
   U1217 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1376, Z => n820);
   U1218 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1376, Z => n819);
   U1219 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1376, Z => n818);
   U1220 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1376, Z => n817);
   U1221 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1376, Z => n816);
   U1222 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1376, Z => n815);
   U1223 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1376, Z => n814);
   U1224 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => n1376, Z => n813);
   U1225 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => n1376, Z => n812);
   U1226 : MUXB2DL port map( A0 => b(21), A1 => b(22), SL => n1376, Z => n811);
   U1227 : MUXB2DL port map( A0 => b(22), A1 => b(23), SL => n1376, Z => n810);
   U1228 : AOI21D1 port map( A1 => a(19), A2 => a(20), B => n1419, Z => n944);
   U1229 : MUXB2DL port map( A0 => b(23), A1 => b(24), SL => n1376, Z => n809);
   U1230 : MUXB2DL port map( A0 => b(24), A1 => b(25), SL => n1376, Z => n808);
   U1231 : NAN2D1 port map( A1 => n1396, A2 => n1377, Z => n807);
   U1232 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1377, Z => n806);
   U1233 : MUXB2DL port map( A0 => b(1), A1 => n1392, SL => n1377, Z => n805);
   U1234 : MUXB2DL port map( A0 => b(2), A1 => n1390, SL => n1377, Z => n804);
   U1235 : MUXB2DL port map( A0 => n1389, A1 => n1387, SL => n1377, Z => n803);
   U1236 : MUXB2DL port map( A0 => n1387, A1 => n1385, SL => n1377, Z => n802);
   U1237 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1377, Z => n801);
   U1238 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1377, Z => n800);
   U1239 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1377, Z => n799);
   U1240 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1377, Z => n798);
   U1241 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1377, Z => n797);
   U1242 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1377, Z => n796);
   U1243 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1377, Z => n795);
   U1244 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1377, Z => n794);
   U1245 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1377, Z => n793);
   U1246 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1377, Z => n792);
   U1247 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1377, Z => n791);
   U1248 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1377, Z => n790);
   U1249 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1377, Z => n789);
   U1250 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1377, Z => n788);
   U1251 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => n1377, Z => n787);
   U1252 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => n1377, Z => n786);
   U1253 : MUXB2DL port map( A0 => b(21), A1 => b(22), SL => n1377, Z => n785);
   U1254 : MUXB2DL port map( A0 => b(22), A1 => b(23), SL => n1377, Z => n784);
   U1255 : NAN2D1 port map( A1 => n1396, A2 => n1447, Z => n783);
   U1256 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1447, Z => n782);
   U1257 : MUXB2DL port map( A0 => n1394, A1 => n1392, SL => n1447, Z => n781);
   U1258 : MUXB2DL port map( A0 => n1392, A1 => n1390, SL => n1447, Z => n780);
   U1259 : MUXB2DL port map( A0 => n1390, A1 => b(4), SL => n1447, Z => n779);
   U1260 : MUXB2DL port map( A0 => n1387, A1 => n1385, SL => n1447, Z => n778);
   U1261 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1447, Z => n777);
   U1262 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1447, Z => n776);
   U1263 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1447, Z => n775);
   U1264 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1447, Z => n774);
   U1265 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1447, Z => n773);
   U1266 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1447, Z => n772);
   U1267 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1447, Z => n771);
   U1268 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1447, Z => n770);
   U1269 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1447, Z => n769);
   U1270 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1447, Z => n768);
   U1271 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1447, Z => n767);
   U1272 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1447, Z => n766);
   U1273 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1447, Z => n765);
   U1274 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1447, Z => n764);
   U1275 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => n1447, Z => n763);
   U1276 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => n1447, Z => n762);
   U1277 : NAN2D1 port map( A1 => n1396, A2 => n1448, Z => n761);
   U1278 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1448, Z => n760);
   U1279 : MUXB2DL port map( A0 => b(1), A1 => n1392, SL => n1448, Z => n759);
   U1280 : MUXB2DL port map( A0 => b(2), A1 => n1390, SL => n1448, Z => n758);
   U1281 : MUXB2DL port map( A0 => n1389, A1 => b(4), SL => n1448, Z => n757);
   U1282 : MUXB2DL port map( A0 => n1387, A1 => n1385, SL => n1448, Z => n756);
   U1283 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1448, Z => n755);
   U1284 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1448, Z => n754);
   U1285 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1448, Z => n753);
   U1286 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1448, Z => n752);
   U1287 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1448, Z => n751);
   U1288 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1448, Z => n750);
   U1289 : AOI21D1 port map( A1 => a(17), A2 => a(18), B => n1417, Z => n945);
   U1290 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1448, Z => n749);
   U1291 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1448, Z => n748);
   U1292 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1448, Z => n747);
   U1293 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1448, Z => n746);
   U1294 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1448, Z => n745);
   U1295 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1448, Z => n744);
   U1296 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1448, Z => n743);
   U1297 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1448, Z => n742);
   U1298 : NAN2D1 port map( A1 => n1396, A2 => n1449, Z => n741);
   U1299 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1449, Z => n740);
   U1300 : MUXB2DL port map( A0 => n1394, A1 => n1392, SL => n1449, Z => n739);
   U1301 : MUXB2DL port map( A0 => b(2), A1 => n1390, SL => n1449, Z => n738);
   U1302 : MUXB2DL port map( A0 => n1389, A1 => b(4), SL => n1449, Z => n737);
   U1303 : MUXB2DL port map( A0 => n1387, A1 => n1385, SL => n1449, Z => n736);
   U1304 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1449, Z => n735);
   U1305 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1449, Z => n734);
   U1306 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1449, Z => n733);
   U1307 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1449, Z => n732);
   U1308 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1449, Z => n731);
   U1309 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1449, Z => n730);
   U1310 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1449, Z => n729);
   U1311 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1449, Z => n728);
   U1312 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1449, Z => n727);
   U1313 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1449, Z => n726);
   U1314 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1449, Z => n725);
   U1315 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1449, Z => n724);
   U1316 : NAN2D1 port map( A1 => n1396, A2 => n1450, Z => n723);
   U1317 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1450, Z => n722);
   U1318 : MUXB2DL port map( A0 => n1394, A1 => n1392, SL => n1450, Z => n721);
   U1319 : MUXB2DL port map( A0 => b(2), A1 => n1390, SL => n1450, Z => n720);
   U1320 : MUXB2DL port map( A0 => n1389, A1 => b(4), SL => n1450, Z => n719);
   U1321 : MUXB2DL port map( A0 => n1387, A1 => n1385, SL => n1450, Z => n718);
   U1322 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1450, Z => n717);
   U1323 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1450, Z => n716);
   U1324 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1450, Z => n715);
   U1325 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1450, Z => n714);
   U1326 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1450, Z => n713);
   U1327 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1450, Z => n712);
   U1328 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1450, Z => n711);
   U1329 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1450, Z => n710);
   U1330 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1450, Z => n709);
   U1331 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1450, Z => n708);
   U1332 : NAN2D1 port map( A1 => n1396, A2 => n1451, Z => n707);
   U1333 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1451, Z => n706);
   U1334 : MUXB2DL port map( A0 => n1394, A1 => n1392, SL => n1451, Z => n705);
   U1335 : MUXB2DL port map( A0 => b(2), A1 => n1390, SL => n1451, Z => n704);
   U1336 : MUXB2DL port map( A0 => n1389, A1 => b(4), SL => n1451, Z => n703);
   U1337 : MUXB2DL port map( A0 => n1387, A1 => n1385, SL => n1451, Z => n702);
   U1338 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1451, Z => n701);
   U1339 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1451, Z => n700);
   U1340 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1451, Z => n699);
   U1341 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1451, Z => n698);
   U1342 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1451, Z => n697);
   U1343 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1451, Z => n696);
   U1344 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1451, Z => n695);
   U1345 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1451, Z => n694);
   U1346 : NAN2D1 port map( A1 => n1396, A2 => n1452, Z => n693);
   U1347 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1452, Z => n692);
   U1348 : MUXB2DL port map( A0 => n1394, A1 => b(2), SL => n1452, Z => n691);
   U1349 : MUXB2DL port map( A0 => b(2), A1 => n1390, SL => n1452, Z => n690);
   U1350 : MUXB2DL port map( A0 => n1389, A1 => b(4), SL => n1452, Z => n689);
   U1351 : MUXB2DL port map( A0 => n1387, A1 => n1385, SL => n1452, Z => n688);
   U1352 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1452, Z => n687);
   U1353 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1452, Z => n686);
   U1354 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1452, Z => n685);
   U1355 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1452, Z => n684);
   U1356 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1452, Z => n683);
   U1357 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1452, Z => n682);
   U1358 : NAN2D1 port map( A1 => n1396, A2 => n1453, Z => n681);
   U1359 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1453, Z => n680);
   U1360 : AOI21D1 port map( A1 => a(15), A2 => a(16), B => n1415, Z => n946);
   U1361 : MUXB2DL port map( A0 => n1394, A1 => b(2), SL => n1453, Z => n679);
   U1362 : MUXB2DL port map( A0 => b(2), A1 => n1390, SL => n1453, Z => n678);
   U1363 : MUXB2DL port map( A0 => n1389, A1 => b(4), SL => n1453, Z => n677);
   U1364 : MUXB2DL port map( A0 => b(4), A1 => n1385, SL => n1453, Z => n676);
   U1365 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1453, Z => n675);
   U1366 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1453, Z => n674);
   U1367 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1453, Z => n673);
   U1368 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1453, Z => n672);
   U1369 : NAN2D1 port map( A1 => b(0), A2 => n1454, Z => n671);
   U1370 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1454, Z => n670);
   U1371 : MUXB2DL port map( A0 => n1394, A1 => b(2), SL => n1454, Z => n669);
   U1372 : MUXB2DL port map( A0 => b(2), A1 => n1390, SL => n1454, Z => n668);
   U1373 : MUXB2DL port map( A0 => n1389, A1 => b(4), SL => n1454, Z => n667);
   U1374 : MUXB2DL port map( A0 => n1387, A1 => b(5), SL => n1454, Z => n666);
   U1375 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1454, Z => n665);
   U1376 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1454, Z => n664);
   U1377 : EXOR2D1 port map( A1 => a(24), A2 => a(23), Z => n1454);
   U1378 : NAN2D1 port map( A1 => b(0), A2 => n1455, Z => n663);
   U1379 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1455, Z => n662);
   U1380 : MUXB2DL port map( A0 => n1394, A1 => b(2), SL => n1455, Z => n661);
   U1381 : MUXB2DL port map( A0 => b(2), A1 => n1390, SL => n1455, Z => n660);
   U1382 : MUXB2DL port map( A0 => n1389, A1 => b(4), SL => n1455, Z => n659);
   U1383 : MUXB2DL port map( A0 => n1387, A1 => n1385, SL => n1455, Z => n658);
   U1384 : EXOR2D1 port map( A1 => a(26), A2 => a(25), Z => n1455);
   U1385 : NAN2D1 port map( A1 => b(0), A2 => n1456, Z => n657);
   U1386 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1456, Z => n656);
   U1387 : MUXB2DL port map( A0 => n1394, A1 => n1392, SL => n1456, Z => n655);
   U1388 : MUXB2DL port map( A0 => b(2), A1 => n1390, SL => n1456, Z => n654);
   U1389 : EXOR2D1 port map( A1 => a(28), A2 => a(27), Z => n1456);
   U1390 : NAN2D1 port map( A1 => b(0), A2 => n1457, Z => n653);
   U1391 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1457, Z => n652);
   U1392 : EXOR2D1 port map( A1 => a(30), A2 => a(29), Z => n1457);
   U1393 : AOI21D1 port map( A1 => a(13), A2 => a(14), B => n1413, Z => n947);
   U1394 : AOI21D1 port map( A1 => a(11), A2 => a(12), B => n1411, Z => n948);
   U1395 : AOI21D1 port map( A1 => a(9), A2 => a(10), B => n1409, Z => n949);
   U1396 : AOI21D1 port map( A1 => a(7), A2 => a(8), B => n1407, Z => n950);
   U1397 : AOI21D1 port map( A1 => a(5), A2 => a(6), B => n1405, Z => n951);
   U1398 : AOI21D1 port map( A1 => a(3), A2 => a(4), B => n1403, Z => n952);
   U1399 : AOI21D1 port map( A1 => a(1), A2 => a(2), B => n1401, Z => n953);
   U1400 : AOI21D1 port map( A1 => a(29), A2 => a(30), B => n1428, Z => n939);
   U1401 : OAI21D1 port map( A1 => a(30), A2 => a(29), B => n1428, Z => n104);
   U1402 : AOI21D1 port map( A1 => a(27), A2 => a(28), B => n1427, Z => n940);

end hier_filter_none_20;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_gp_custom.all;

architecture hier_filter_none_20 of gp_custom_DW_mult_tc_0 is

   component AOI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component MUXB2DL
      port( A0, A1, SL : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal n42, n50, n58, n66, n73, n80, n84, n89, n94, n99, n104, n156, n157, 
      n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, 
      n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, 
      n182, n183, n184, n185, n186, n202, n203, n204, n205, n206, n207, n208, 
      n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, 
      n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, 
      n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, 
      n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, 
      n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, 
      n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, 
      n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
      n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, 
      n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, 
      n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, 
      n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, 
      n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, 
      n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, 
      n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, 
      n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, 
      n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, 
      n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, 
      n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, 
      n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, 
      n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, 
      n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, 
      n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, 
      n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, 
      n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, 
      n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, 
      n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, 
      n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
      n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, 
      n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, 
      n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, 
      n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
      n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, 
      n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, 
      n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, 
      n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, 
      n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, 
      n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, 
      n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, 
      n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, 
      n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, 
      n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, 
      n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, 
      n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, 
      n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, 
      n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, 
      n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, 
      n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, 
      n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, 
      n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, 
      n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, 
      n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, 
      n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, 
      n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, 
      n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, 
      n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, 
      n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, 
      n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, 
      n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, 
      n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, 
      n917, n918, n919, n920, n921, n922, n923, n939, n940, n941, n942, n943, 
      n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n955, n956, 
      n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, 
      n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, 
      n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, 
      n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, 
      n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, 
      n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, 
      n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, 
      n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, 
      n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, 
      n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, 
      n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, 
      n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, 
      n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, 
      n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, 
      n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, 
      n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, 
      n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, 
      n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, 
      n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, 
      n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, 
      n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, 
      n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, 
      n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, 
      n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, 
      n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, 
      n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, 
      n1224, n1225, n1226, n1375, n1376, n1377, n1378, n1379, n1380, n1381, 
      n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, 
      n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, 
      n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, 
      n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, 
      n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, 
      n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, 
      n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, 
      n1452, n1453, n1454 : std_logic;

begin
   
   U125 : ADFULD1 port map( A => n203, B => n232, CI => n157, CO => n156, S => 
                           product(30));
   U126 : ADFULD1 port map( A => n233, B => n260, CI => n158, CO => n157, S => 
                           product(29));
   U127 : ADFULD1 port map( A => n261, B => n288, CI => n159, CO => n158, S => 
                           product(28));
   U128 : ADFULD1 port map( A => n289, B => n314, CI => n160, CO => n159, S => 
                           product(27));
   U129 : ADFULD1 port map( A => n315, B => n340, CI => n161, CO => n160, S => 
                           product(26));
   U130 : ADFULD1 port map( A => n341, B => n364, CI => n162, CO => n161, S => 
                           product(25));
   U131 : ADFULD1 port map( A => n365, B => n388, CI => n163, CO => n162, S => 
                           product(24));
   U132 : ADFULD1 port map( A => n389, B => n410, CI => n164, CO => n163, S => 
                           product(23));
   U133 : ADFULD1 port map( A => n411, B => n432, CI => n165, CO => n164, S => 
                           product(22));
   U134 : ADFULD1 port map( A => n433, B => n452, CI => n166, CO => n165, S => 
                           product(21));
   U135 : ADFULD1 port map( A => n453, B => n472, CI => n167, CO => n166, S => 
                           product(20));
   U136 : ADFULD1 port map( A => n473, B => n490, CI => n168, CO => n167, S => 
                           product(19));
   U137 : ADFULD1 port map( A => n491, B => n508, CI => n169, CO => n168, S => 
                           product(18));
   U138 : ADFULD1 port map( A => n509, B => n524, CI => n170, CO => n169, S => 
                           product(17));
   U139 : ADFULD1 port map( A => n525, B => n540, CI => n171, CO => n170, S => 
                           product(16));
   U140 : ADFULD1 port map( A => n541, B => n554, CI => n172, CO => n171, S => 
                           product(15));
   U141 : ADFULD1 port map( A => n555, B => n568, CI => n173, CO => n172, S => 
                           product(14));
   U142 : ADFULD1 port map( A => n569, B => n580, CI => n174, CO => n173, S => 
                           product(13));
   U143 : ADFULD1 port map( A => n581, B => n592, CI => n175, CO => n174, S => 
                           product(12));
   U144 : ADFULD1 port map( A => n593, B => n602, CI => n176, CO => n175, S => 
                           product(11));
   U145 : ADFULD1 port map( A => n603, B => n612, CI => n177, CO => n176, S => 
                           product(10));
   U146 : ADFULD1 port map( A => n613, B => n620, CI => n178, CO => n177, S => 
                           product(9));
   U147 : ADFULD1 port map( A => n621, B => n628, CI => n179, CO => n178, S => 
                           product(8));
   U148 : ADFULD1 port map( A => n629, B => n634, CI => n180, CO => n179, S => 
                           product(7));
   U149 : ADFULD1 port map( A => n635, B => n640, CI => n181, CO => n180, S => 
                           product(6));
   U150 : ADFULD1 port map( A => n641, B => n644, CI => n182, CO => n181, S => 
                           product(5));
   U151 : ADFULD1 port map( A => n645, B => n648, CI => n183, CO => n182, S => 
                           product(4));
   U152 : ADFULD1 port map( A => n649, B => n1193, CI => n184, CO => n183, S =>
                           product(3));
   U153 : ADFULD1 port map( A => n651, B => n1194, CI => n185, CO => n184, S =>
                           product(2));
   U154 : ADHALFDL port map( A => n186, B => n1225, CO => n185, S => product(1)
                           );
   U155 : ADHALFDL port map( A => n1226, B => a(1), CO => n186, S => product(0)
                           );
   U171 : ADFULD1 port map( A => n234, B => n207, CI => n205, CO => n202, S => 
                           n203);
   U172 : ADFULD1 port map( A => n209, B => n211, CI => n236, CO => n204, S => 
                           n205);
   U173 : ADFULD1 port map( A => n240, B => n213, CI => n238, CO => n206, S => 
                           n207);
   U174 : ADFULD1 port map( A => n217, B => n242, CI => n215, CO => n208, S => 
                           n209);
   U175 : ADFULD1 port map( A => n244, B => n246, CI => n219, CO => n210, S => 
                           n211);
   U176 : ADFULD1 port map( A => n225, B => n223, CI => n248, CO => n212, S => 
                           n213);
   U177 : ADFULD1 port map( A => n221, B => n229, CI => n227, CO => n214, S => 
                           n215);
   U178 : ADFULD1 port map( A => n256, B => n252, CI => n254, CO => n216, S => 
                           n217);
   U179 : ADFULD1 port map( A => n258, B => n1088, CI => n250, CO => n218, S =>
                           n219);
   U180 : ADFULD1 port map( A => n1046, B => n1112, CI => n1066, CO => n220, S 
                           => n221);
   U181 : ADFULD1 port map( A => n986, B => n976, CI => n998, CO => n222, S => 
                           n223);
   U182 : ADFULD1 port map( A => n962, B => n1138, CI => n968, CO => n224, S =>
                           n225);
   U183 : ADFULD1 port map( A => n1166, B => n1012, CI => n231, CO => n226, S 
                           => n227);
   U184 : ADFULD1 port map( A => n1028, B => n956, CI => n958, CO => n228, S =>
                           n229);
   U185 : ADHALFDL port map( A => n1196, B => n939, CO => n230, S => n231);
   U186 : ADFULD1 port map( A => n262, B => n237, CI => n235, CO => n232, S => 
                           n233);
   U187 : ADFULD1 port map( A => n239, B => n266, CI => n264, CO => n234, S => 
                           n235);
   U188 : ADFULD1 port map( A => n268, B => n243, CI => n241, CO => n236, S => 
                           n237);
   U189 : ADFULD1 port map( A => n270, B => n247, CI => n245, CO => n238, S => 
                           n239);
   U190 : ADFULD1 port map( A => n274, B => n249, CI => n272, CO => n240, S => 
                           n241);
   U191 : ADFULD1 port map( A => n253, B => n255, CI => n257, CO => n242, S => 
                           n243);
   U192 : ADFULD1 port map( A => n280, B => n276, CI => n251, CO => n244, S => 
                           n245);
   U193 : ADFULD1 port map( A => n278, B => n284, CI => n282, CO => n246, S => 
                           n247);
   U194 : ADFULD1 port map( A => n1047, B => n1013, CI => n259, CO => n248, S 
                           => n249);
   U195 : ADFULD1 port map( A => n977, B => n1067, CI => n999, CO => n250, S =>
                           n251);
   U196 : ADFULD1 port map( A => n959, B => n969, CI => n963, CO => n252, S => 
                           n253);
   U197 : ADFULD1 port map( A => n1113, B => n987, CI => n1089, CO => n254, S 
                           => n255);
   U198 : ADFULD1 port map( A => n1167, B => n1029, CI => n1139, CO => n256, S 
                           => n257);
   U199 : ADHALFDL port map( A => n286, B => n1197, CO => n258, S => n259);
   U200 : ADFULD1 port map( A => n290, B => n265, CI => n263, CO => n260, S => 
                           n261);
   U201 : ADFULD1 port map( A => n267, B => n294, CI => n292, CO => n262, S => 
                           n263);
   U202 : ADFULD1 port map( A => n296, B => n271, CI => n269, CO => n264, S => 
                           n265);
   U203 : ADFULD1 port map( A => n275, B => n298, CI => n273, CO => n266, S => 
                           n267);
   U204 : ADFULD1 port map( A => n302, B => n281, CI => n300, CO => n268, S => 
                           n269);
   U205 : ADFULD1 port map( A => n283, B => n277, CI => n279, CO => n270, S => 
                           n271);
   U206 : ADFULD1 port map( A => n310, B => n308, CI => n285, CO => n272, S => 
                           n273);
   U207 : ADFULD1 port map( A => n304, B => n312, CI => n306, CO => n274, S => 
                           n275);
   U208 : ADFULD1 port map( A => n1014, B => n1068, CI => n1048, CO => n276, S 
                           => n277);
   U209 : ADFULD1 port map( A => n978, B => n1090, CI => n988, CO => n278, S =>
                           n279);
   U210 : ADFULD1 port map( A => n964, B => n1114, CI => n970, CO => n280, S =>
                           n281);
   U211 : ADFULD1 port map( A => n1140, B => n1000, CI => n287, CO => n282, S 
                           => n283);
   U212 : ADFULD1 port map( A => n1030, B => n960, CI => n1168, CO => n284, S 
                           => n285);
   U213 : ADHALFDL port map( A => n1198, B => n940, CO => n286, S => n287);
   U214 : ADFULD1 port map( A => n316, B => n293, CI => n291, CO => n288, S => 
                           n289);
   U215 : ADFULD1 port map( A => n318, B => n297, CI => n295, CO => n290, S => 
                           n291);
   U216 : ADFULD1 port map( A => n299, B => n322, CI => n320, CO => n292, S => 
                           n293);
   U217 : ADFULD1 port map( A => n324, B => n303, CI => n301, CO => n294, S => 
                           n295);
   U218 : ADFULD1 port map( A => n307, B => n309, CI => n326, CO => n296, S => 
                           n297);
   U219 : ADFULD1 port map( A => n305, B => n328, CI => n311, CO => n298, S => 
                           n299);
   U220 : ADFULD1 port map( A => n332, B => n330, CI => n334, CO => n300, S => 
                           n301);
   U221 : ADFULD1 port map( A => n313, B => n1091, CI => n336, CO => n302, S =>
                           n303);
   U222 : ADFULD1 port map( A => n1015, B => n1115, CI => n1069, CO => n304, S 
                           => n305);
   U223 : ADFULD1 port map( A => n1141, B => n1001, CI => n989, CO => n306, S 
                           => n307);
   U224 : ADFULD1 port map( A => n979, B => n1049, CI => n1169, CO => n308, S 
                           => n309);
   U225 : ADFULD1 port map( A => n965, B => n1031, CI => n971, CO => n310, S =>
                           n311);
   U226 : ADHALFDL port map( A => n338, B => n1199, CO => n312, S => n313);
   U227 : ADFULD1 port map( A => n342, B => n319, CI => n317, CO => n314, S => 
                           n315);
   U228 : ADFULD1 port map( A => n344, B => n346, CI => n321, CO => n316, S => 
                           n317);
   U229 : ADFULD1 port map( A => n325, B => n327, CI => n323, CO => n318, S => 
                           n319);
   U230 : ADFULD1 port map( A => n350, B => n352, CI => n348, CO => n320, S => 
                           n321);
   U231 : ADFULD1 port map( A => n333, B => n335, CI => n329, CO => n322, S => 
                           n323);
   U232 : ADFULD1 port map( A => n337, B => n358, CI => n331, CO => n324, S => 
                           n325);
   U233 : ADFULD1 port map( A => n354, B => n360, CI => n356, CO => n326, S => 
                           n327);
   U234 : ADFULD1 port map( A => n1092, B => n1116, CI => n362, CO => n328, S 
                           => n329);
   U235 : ADFULD1 port map( A => n1016, B => n1142, CI => n1070, CO => n330, S 
                           => n331);
   U236 : ADFULD1 port map( A => n990, B => n1170, CI => n1002, CO => n332, S 
                           => n333);
   U237 : ADFULD1 port map( A => n980, B => n1032, CI => n339, CO => n334, S =>
                           n335);
   U238 : ADFULD1 port map( A => n1050, B => n966, CI => n972, CO => n336, S =>
                           n337);
   U239 : ADHALFDL port map( A => n1200, B => n941, CO => n338, S => n339);
   U240 : ADFULD1 port map( A => n366, B => n345, CI => n343, CO => n340, S => 
                           n341);
   U241 : ADFULD1 port map( A => n347, B => n370, CI => n368, CO => n342, S => 
                           n343);
   U242 : ADFULD1 port map( A => n351, B => n372, CI => n349, CO => n344, S => 
                           n345);
   U243 : ADFULD1 port map( A => n374, B => n376, CI => n353, CO => n346, S => 
                           n347);
   U244 : ADFULD1 port map( A => n361, B => n357, CI => n359, CO => n348, S => 
                           n349);
   U245 : ADFULD1 port map( A => n378, B => n380, CI => n355, CO => n350, S => 
                           n351);
   U246 : ADFULD1 port map( A => n384, B => n363, CI => n382, CO => n352, S => 
                           n353);
   U247 : ADFULD1 port map( A => n1033, B => n1093, CI => n1071, CO => n354, S 
                           => n355);
   U248 : ADFULD1 port map( A => n991, B => n1117, CI => n1017, CO => n356, S 
                           => n357);
   U249 : ADFULD1 port map( A => n973, B => n1003, CI => n981, CO => n358, S =>
                           n359);
   U250 : ADFULD1 port map( A => n1171, B => n1051, CI => n1143, CO => n360, S 
                           => n361);
   U251 : ADHALFDL port map( A => n386, B => n1201, CO => n362, S => n363);
   U252 : ADFULD1 port map( A => n390, B => n369, CI => n367, CO => n364, S => 
                           n365);
   U253 : ADFULD1 port map( A => n371, B => n394, CI => n392, CO => n366, S => 
                           n367);
   U254 : ADFULD1 port map( A => n375, B => n396, CI => n373, CO => n368, S => 
                           n369);
   U255 : ADFULD1 port map( A => n398, B => n400, CI => n377, CO => n370, S => 
                           n371);
   U256 : ADFULD1 port map( A => n383, B => n379, CI => n381, CO => n372, S => 
                           n373);
   U257 : ADFULD1 port map( A => n402, B => n404, CI => n385, CO => n374, S => 
                           n375);
   U258 : ADFULD1 port map( A => n408, B => n1072, CI => n406, CO => n376, S =>
                           n377);
   U259 : ADFULD1 port map( A => n1004, B => n1094, CI => n1034, CO => n378, S 
                           => n379);
   U260 : ADFULD1 port map( A => n992, B => n1144, CI => n1118, CO => n380, S 
                           => n381);
   U261 : ADFULD1 port map( A => n982, B => n1018, CI => n387, CO => n382, S =>
                           n383);
   U262 : ADFULD1 port map( A => n1052, B => n974, CI => n1172, CO => n384, S 
                           => n385);
   U263 : ADHALFDL port map( A => n1202, B => n942, CO => n386, S => n387);
   U264 : ADFULD1 port map( A => n412, B => n393, CI => n391, CO => n388, S => 
                           n389);
   U265 : ADFULD1 port map( A => n395, B => n397, CI => n414, CO => n390, S => 
                           n391);
   U266 : ADFULD1 port map( A => n399, B => n418, CI => n416, CO => n392, S => 
                           n393);
   U267 : ADFULD1 port map( A => n401, B => n407, CI => n420, CO => n394, S => 
                           n395);
   U268 : ADFULD1 port map( A => n403, B => n424, CI => n405, CO => n396, S => 
                           n397);
   U269 : ADFULD1 port map( A => n426, B => n428, CI => n422, CO => n398, S => 
                           n399);
   U270 : ADFULD1 port map( A => n1073, B => n1095, CI => n409, CO => n400, S 
                           => n401);
   U271 : ADFULD1 port map( A => n1005, B => n1119, CI => n1019, CO => n402, S 
                           => n403);
   U272 : ADFULD1 port map( A => n1173, B => n1035, CI => n1145, CO => n404, S 
                           => n405);
   U273 : ADFULD1 port map( A => n983, B => n1053, CI => n993, CO => n406, S =>
                           n407);
   U274 : ADHALFDL port map( A => n430, B => n1203, CO => n408, S => n409);
   U275 : ADFULD1 port map( A => n434, B => n415, CI => n413, CO => n410, S => 
                           n411);
   U276 : ADFULD1 port map( A => n417, B => n419, CI => n436, CO => n412, S => 
                           n413);
   U277 : ADFULD1 port map( A => n421, B => n440, CI => n438, CO => n414, S => 
                           n415);
   U278 : ADFULD1 port map( A => n427, B => n425, CI => n442, CO => n416, S => 
                           n417);
   U279 : ADFULD1 port map( A => n429, B => n444, CI => n423, CO => n418, S => 
                           n419);
   U280 : ADFULD1 port map( A => n448, B => n450, CI => n446, CO => n420, S => 
                           n421);
   U281 : ADFULD1 port map( A => n1074, B => n1120, CI => n1096, CO => n422, S 
                           => n423);
   U282 : ADFULD1 port map( A => n1006, B => n1146, CI => n1020, CO => n424, S 
                           => n425);
   U283 : ADFULD1 port map( A => n1174, B => n1036, CI => n431, CO => n426, S 
                           => n427);
   U284 : ADFULD1 port map( A => n1054, B => n984, CI => n994, CO => n428, S =>
                           n429);
   U285 : ADHALFDL port map( A => n1204, B => n943, CO => n430, S => n431);
   U286 : ADFULD1 port map( A => n454, B => n437, CI => n435, CO => n432, S => 
                           n433);
   U287 : ADFULD1 port map( A => n439, B => n441, CI => n456, CO => n434, S => 
                           n435);
   U288 : ADFULD1 port map( A => n443, B => n460, CI => n458, CO => n436, S => 
                           n437);
   U289 : ADFULD1 port map( A => n449, B => n445, CI => n447, CO => n438, S => 
                           n439);
   U290 : ADFULD1 port map( A => n464, B => n466, CI => n462, CO => n440, S => 
                           n441);
   U291 : ADFULD1 port map( A => n451, B => n1037, CI => n468, CO => n442, S =>
                           n443);
   U292 : ADFULD1 port map( A => n995, B => n1075, CI => n1007, CO => n444, S 
                           => n445);
   U293 : ADFULD1 port map( A => n1121, B => n1021, CI => n1097, CO => n446, S 
                           => n447);
   U294 : ADFULD1 port map( A => n1175, B => n1055, CI => n1147, CO => n448, S 
                           => n449);
   U295 : ADHALFDL port map( A => n470, B => n1205, CO => n450, S => n451);
   U296 : ADFULD1 port map( A => n474, B => n457, CI => n455, CO => n452, S => 
                           n453);
   U297 : ADFULD1 port map( A => n459, B => n461, CI => n476, CO => n454, S => 
                           n455);
   U298 : ADFULD1 port map( A => n480, B => n463, CI => n478, CO => n456, S => 
                           n457);
   U299 : ADFULD1 port map( A => n465, B => n469, CI => n467, CO => n458, S => 
                           n459);
   U300 : ADFULD1 port map( A => n482, B => n486, CI => n484, CO => n460, S => 
                           n461);
   U301 : ADFULD1 port map( A => n1098, B => n1122, CI => n488, CO => n462, S 
                           => n463);
   U302 : ADFULD1 port map( A => n1022, B => n1148, CI => n1056, CO => n464, S 
                           => n465);
   U303 : ADFULD1 port map( A => n1008, B => n1038, CI => n471, CO => n466, S 
                           => n467);
   U304 : ADFULD1 port map( A => n1076, B => n996, CI => n1176, CO => n468, S 
                           => n469);
   U305 : ADHALFDL port map( A => n1206, B => n944, CO => n470, S => n471);
   U306 : ADFULD1 port map( A => n492, B => n477, CI => n475, CO => n472, S => 
                           n473);
   U307 : ADFULD1 port map( A => n479, B => n481, CI => n494, CO => n474, S => 
                           n475);
   U308 : ADFULD1 port map( A => n498, B => n487, CI => n496, CO => n476, S => 
                           n477);
   U309 : ADFULD1 port map( A => n483, B => n500, CI => n485, CO => n478, S => 
                           n479);
   U310 : ADFULD1 port map( A => n504, B => n489, CI => n502, CO => n480, S => 
                           n481);
   U311 : ADFULD1 port map( A => n1057, B => n1149, CI => n1123, CO => n482, S 
                           => n483);
   U312 : ADFULD1 port map( A => n1177, B => n1099, CI => n1039, CO => n484, S 
                           => n485);
   U313 : ADFULD1 port map( A => n1009, B => n1077, CI => n1023, CO => n486, S 
                           => n487);
   U314 : ADHALFDL port map( A => n506, B => n1207, CO => n488, S => n489);
   U315 : ADFULD1 port map( A => n510, B => n495, CI => n493, CO => n490, S => 
                           n491);
   U316 : ADFULD1 port map( A => n497, B => n499, CI => n512, CO => n492, S => 
                           n493);
   U317 : ADFULD1 port map( A => n516, B => n503, CI => n514, CO => n494, S => 
                           n495);
   U318 : ADFULD1 port map( A => n505, B => n518, CI => n501, CO => n496, S => 
                           n497);
   U319 : ADFULD1 port map( A => n522, B => n1124, CI => n520, CO => n498, S =>
                           n499);
   U320 : ADFULD1 port map( A => n1040, B => n1150, CI => n1058, CO => n500, S 
                           => n501);
   U321 : ADFULD1 port map( A => n1178, B => n1100, CI => n507, CO => n502, S 
                           => n503);
   U322 : ADFULD1 port map( A => n1078, B => n1010, CI => n1024, CO => n504, S 
                           => n505);
   U323 : ADHALFDL port map( A => n1208, B => n945, CO => n506, S => n507);
   U324 : ADFULD1 port map( A => n526, B => n513, CI => n511, CO => n508, S => 
                           n509);
   U325 : ADFULD1 port map( A => n528, B => n530, CI => n515, CO => n510, S => 
                           n511);
   U326 : ADFULD1 port map( A => n521, B => n519, CI => n517, CO => n512, S => 
                           n513);
   U327 : ADFULD1 port map( A => n534, B => n536, CI => n532, CO => n514, S => 
                           n515);
   U328 : ADFULD1 port map( A => n1101, B => n1125, CI => n523, CO => n516, S 
                           => n517);
   U329 : ADFULD1 port map( A => n1025, B => n1041, CI => n1059, CO => n518, S 
                           => n519);
   U330 : ADFULD1 port map( A => n1179, B => n1079, CI => n1151, CO => n520, S 
                           => n521);
   U331 : ADHALFDL port map( A => n538, B => n1209, CO => n522, S => n523);
   U332 : ADFULD1 port map( A => n542, B => n529, CI => n527, CO => n524, S => 
                           n525);
   U333 : ADFULD1 port map( A => n544, B => n546, CI => n531, CO => n526, S => 
                           n527);
   U334 : ADFULD1 port map( A => n533, B => n537, CI => n535, CO => n528, S => 
                           n529);
   U335 : ADFULD1 port map( A => n550, B => n552, CI => n548, CO => n530, S => 
                           n531);
   U336 : ADFULD1 port map( A => n1080, B => n1152, CI => n1126, CO => n532, S 
                           => n533);
   U337 : ADFULD1 port map( A => n1042, B => n1060, CI => n539, CO => n534, S 
                           => n535);
   U338 : ADFULD1 port map( A => n1102, B => n1026, CI => n1180, CO => n536, S 
                           => n537);
   U339 : ADHALFDL port map( A => n1210, B => n946, CO => n538, S => n539);
   U340 : ADFULD1 port map( A => n556, B => n545, CI => n543, CO => n540, S => 
                           n541);
   U341 : ADFULD1 port map( A => n547, B => n551, CI => n558, CO => n542, S => 
                           n543);
   U342 : ADFULD1 port map( A => n560, B => n562, CI => n549, CO => n544, S => 
                           n545);
   U343 : ADFULD1 port map( A => n553, B => n1153, CI => n564, CO => n546, S =>
                           n547);
   U344 : ADFULD1 port map( A => n1181, B => n1081, CI => n1127, CO => n548, S 
                           => n549);
   U345 : ADFULD1 port map( A => n1043, B => n1103, CI => n1061, CO => n550, S 
                           => n551);
   U346 : ADHALFDL port map( A => n566, B => n1211, CO => n552, S => n553);
   U347 : ADFULD1 port map( A => n570, B => n559, CI => n557, CO => n554, S => 
                           n555);
   U348 : ADFULD1 port map( A => n561, B => n563, CI => n572, CO => n556, S => 
                           n557);
   U349 : ADFULD1 port map( A => n574, B => n576, CI => n565, CO => n558, S => 
                           n559);
   U350 : ADFULD1 port map( A => n1062, B => n1128, CI => n578, CO => n560, S 
                           => n561);
   U351 : ADFULD1 port map( A => n1154, B => n1082, CI => n567, CO => n562, S 
                           => n563);
   U352 : ADFULD1 port map( A => n1104, B => n1044, CI => n1182, CO => n564, S 
                           => n565);
   U353 : ADHALFDL port map( A => n1212, B => n947, CO => n566, S => n567);
   U354 : ADFULD1 port map( A => n582, B => n573, CI => n571, CO => n568, S => 
                           n569);
   U355 : ADFULD1 port map( A => n577, B => n575, CI => n584, CO => n570, S => 
                           n571);
   U356 : ADFULD1 port map( A => n588, B => n579, CI => n586, CO => n572, S => 
                           n573);
   U357 : ADFULD1 port map( A => n1063, B => n1129, CI => n1083, CO => n574, S 
                           => n575);
   U358 : ADFULD1 port map( A => n1183, B => n1105, CI => n1155, CO => n576, S 
                           => n577);
   U359 : ADHALFDL port map( A => n590, B => n1213, CO => n578, S => n579);
   U360 : ADFULD1 port map( A => n585, B => n594, CI => n583, CO => n580, S => 
                           n581);
   U361 : ADFULD1 port map( A => n587, B => n589, CI => n596, CO => n582, S => 
                           n583);
   U362 : ADFULD1 port map( A => n600, B => n1106, CI => n598, CO => n584, S =>
                           n585);
   U363 : ADFULD1 port map( A => n1084, B => n1156, CI => n591, CO => n586, S 
                           => n587);
   U364 : ADFULD1 port map( A => n1130, B => n1064, CI => n1184, CO => n588, S 
                           => n589);
   U365 : ADHALFDL port map( A => n1214, B => n948, CO => n590, S => n591);
   U366 : ADFULD1 port map( A => n604, B => n597, CI => n595, CO => n592, S => 
                           n593);
   U367 : ADFULD1 port map( A => n606, B => n608, CI => n599, CO => n594, S => 
                           n595);
   U368 : ADFULD1 port map( A => n1107, B => n1157, CI => n601, CO => n596, S 
                           => n597);
   U369 : ADFULD1 port map( A => n1085, B => n1131, CI => n1185, CO => n598, S 
                           => n599);
   U370 : ADHALFDL port map( A => n610, B => n1215, CO => n600, S => n601);
   U371 : ADFULD1 port map( A => n614, B => n607, CI => n605, CO => n602, S => 
                           n603);
   U372 : ADFULD1 port map( A => n616, B => n618, CI => n609, CO => n604, S => 
                           n605);
   U373 : ADFULD1 port map( A => n1108, B => n1158, CI => n611, CO => n606, S 
                           => n607);
   U374 : ADFULD1 port map( A => n1132, B => n1086, CI => n1186, CO => n608, S 
                           => n609);
   U375 : ADHALFDL port map( A => n1216, B => n949, CO => n610, S => n611);
   U376 : ADFULD1 port map( A => n617, B => n622, CI => n615, CO => n612, S => 
                           n613);
   U377 : ADFULD1 port map( A => n619, B => n1187, CI => n624, CO => n614, S =>
                           n615);
   U378 : ADFULD1 port map( A => n1109, B => n1133, CI => n1159, CO => n616, S 
                           => n617);
   U379 : ADHALFDL port map( A => n626, B => n1217, CO => n618, S => n619);
   U380 : ADFULD1 port map( A => n625, B => n630, CI => n623, CO => n620, S => 
                           n621);
   U381 : ADFULD1 port map( A => n627, B => n1160, CI => n632, CO => n622, S =>
                           n623);
   U382 : ADFULD1 port map( A => n1188, B => n1110, CI => n1134, CO => n624, S 
                           => n625);
   U383 : ADHALFDL port map( A => n1218, B => n950, CO => n626, S => n627);
   U384 : ADFULD1 port map( A => n636, B => n633, CI => n631, CO => n628, S => 
                           n629);
   U385 : ADFULD1 port map( A => n1135, B => n1189, CI => n1161, CO => n630, S 
                           => n631);
   U386 : ADHALFDL port map( A => n638, B => n1219, CO => n632, S => n633);
   U387 : ADFULD1 port map( A => n642, B => n639, CI => n637, CO => n634, S => 
                           n635);
   U388 : ADFULD1 port map( A => n1190, B => n1136, CI => n1162, CO => n636, S 
                           => n637);
   U389 : ADHALFDL port map( A => n1220, B => n951, CO => n638, S => n639);
   U390 : ADFULD1 port map( A => n1163, B => n1191, CI => n643, CO => n640, S 
                           => n641);
   U391 : ADHALFDL port map( A => n646, B => n1221, CO => n642, S => n643);
   U392 : ADFULD1 port map( A => n1192, B => n1164, CI => n647, CO => n644, S 
                           => n645);
   U393 : ADHALFDL port map( A => n1222, B => n952, CO => n646, S => n647);
   U394 : ADHALFDL port map( A => n650, B => n1223, CO => n648, S => n649);
   U395 : ADHALFDL port map( A => n1224, B => n953, CO => n650, S => n651);
   U397 : MUXB2DL port map( A0 => n104, A1 => n1423, SL => n652, Z => n955);
   U399 : MUXB2DL port map( A0 => n104, A1 => n1423, SL => n653, Z => n956);
   U402 : MUXB2DL port map( A0 => n99, A1 => n1422, SL => n654, Z => n957);
   U404 : MUXB2DL port map( A0 => n99, A1 => n1422, SL => n655, Z => n958);
   U406 : MUXB2DL port map( A0 => n99, A1 => n1422, SL => n656, Z => n959);
   U408 : MUXB2DL port map( A0 => n99, A1 => n1422, SL => n657, Z => n960);
   U411 : MUXB2DL port map( A0 => n94, A1 => n1419, SL => n658, Z => n961);
   U413 : MUXB2DL port map( A0 => n94, A1 => n1419, SL => n659, Z => n962);
   U415 : MUXB2DL port map( A0 => n94, A1 => n1419, SL => n660, Z => n963);
   U417 : MUXB2DL port map( A0 => n94, A1 => n1419, SL => n661, Z => n964);
   U419 : MUXB2DL port map( A0 => n94, A1 => n1419, SL => n662, Z => n965);
   U421 : MUXB2DL port map( A0 => n94, A1 => n1419, SL => n663, Z => n966);
   U424 : MUXB2DL port map( A0 => n89, A1 => n1417, SL => n664, Z => n967);
   U426 : MUXB2DL port map( A0 => n89, A1 => n1417, SL => n665, Z => n968);
   U428 : MUXB2DL port map( A0 => n89, A1 => n1417, SL => n666, Z => n969);
   U430 : MUXB2DL port map( A0 => n89, A1 => n1417, SL => n667, Z => n970);
   U432 : MUXB2DL port map( A0 => n89, A1 => n1417, SL => n668, Z => n971);
   U434 : MUXB2DL port map( A0 => n89, A1 => n1417, SL => n669, Z => n972);
   U436 : MUXB2DL port map( A0 => n89, A1 => n1417, SL => n670, Z => n973);
   U438 : MUXB2DL port map( A0 => n89, A1 => n1417, SL => n671, Z => n974);
   U441 : MUXB2DL port map( A0 => n84, A1 => n1415, SL => n672, Z => n975);
   U443 : MUXB2DL port map( A0 => n84, A1 => n1415, SL => n673, Z => n976);
   U445 : MUXB2DL port map( A0 => n84, A1 => n1415, SL => n674, Z => n977);
   U447 : MUXB2DL port map( A0 => n84, A1 => n1415, SL => n675, Z => n978);
   U449 : MUXB2DL port map( A0 => n84, A1 => n1415, SL => n676, Z => n979);
   U451 : MUXB2DL port map( A0 => n84, A1 => n1415, SL => n677, Z => n980);
   U453 : MUXB2DL port map( A0 => n84, A1 => n1415, SL => n678, Z => n981);
   U455 : MUXB2DL port map( A0 => n84, A1 => n1415, SL => n679, Z => n982);
   U457 : MUXB2DL port map( A0 => n84, A1 => n1415, SL => n680, Z => n983);
   U459 : MUXB2DL port map( A0 => n84, A1 => n1415, SL => n681, Z => n984);
   U462 : MUXB2DL port map( A0 => n80, A1 => n1413, SL => n682, Z => n985);
   U464 : MUXB2DL port map( A0 => n80, A1 => n1413, SL => n683, Z => n986);
   U466 : MUXB2DL port map( A0 => n80, A1 => n1413, SL => n684, Z => n987);
   U468 : MUXB2DL port map( A0 => n80, A1 => n1413, SL => n685, Z => n988);
   U470 : MUXB2DL port map( A0 => n80, A1 => n1413, SL => n686, Z => n989);
   U472 : MUXB2DL port map( A0 => n80, A1 => n1413, SL => n687, Z => n990);
   U474 : MUXB2DL port map( A0 => n80, A1 => n1413, SL => n688, Z => n991);
   U476 : MUXB2DL port map( A0 => n80, A1 => n1413, SL => n689, Z => n992);
   U478 : MUXB2DL port map( A0 => n80, A1 => n1413, SL => n690, Z => n993);
   U480 : MUXB2DL port map( A0 => n80, A1 => n1413, SL => n691, Z => n994);
   U482 : MUXB2DL port map( A0 => n80, A1 => n1413, SL => n692, Z => n995);
   U484 : MUXB2DL port map( A0 => n80, A1 => n1413, SL => n693, Z => n996);
   U487 : MUXB2DL port map( A0 => n73, A1 => n1411, SL => n694, Z => n997);
   U489 : MUXB2DL port map( A0 => n73, A1 => n1411, SL => n695, Z => n998);
   U491 : MUXB2DL port map( A0 => n73, A1 => n1411, SL => n696, Z => n999);
   U493 : MUXB2DL port map( A0 => n73, A1 => n1411, SL => n697, Z => n1000);
   U495 : MUXB2DL port map( A0 => n73, A1 => n1411, SL => n698, Z => n1001);
   U497 : MUXB2DL port map( A0 => n73, A1 => n1411, SL => n699, Z => n1002);
   U499 : MUXB2DL port map( A0 => n73, A1 => n1411, SL => n700, Z => n1003);
   U501 : MUXB2DL port map( A0 => n73, A1 => n1411, SL => n701, Z => n1004);
   U503 : MUXB2DL port map( A0 => n73, A1 => n1411, SL => n702, Z => n1005);
   U505 : MUXB2DL port map( A0 => n73, A1 => n1411, SL => n703, Z => n1006);
   U507 : MUXB2DL port map( A0 => n73, A1 => n1411, SL => n704, Z => n1007);
   U509 : MUXB2DL port map( A0 => n73, A1 => n1411, SL => n705, Z => n1008);
   U511 : MUXB2DL port map( A0 => n73, A1 => n1411, SL => n706, Z => n1009);
   U513 : MUXB2DL port map( A0 => n73, A1 => n1411, SL => n707, Z => n1010);
   U516 : MUXB2DL port map( A0 => n66, A1 => n1409, SL => n708, Z => n1011);
   U518 : MUXB2DL port map( A0 => n66, A1 => n1409, SL => n709, Z => n1012);
   U520 : MUXB2DL port map( A0 => n66, A1 => n1409, SL => n710, Z => n1013);
   U522 : MUXB2DL port map( A0 => n66, A1 => n1409, SL => n711, Z => n1014);
   U524 : MUXB2DL port map( A0 => n66, A1 => n1409, SL => n712, Z => n1015);
   U526 : MUXB2DL port map( A0 => n66, A1 => n1409, SL => n713, Z => n1016);
   U528 : MUXB2DL port map( A0 => n66, A1 => n1409, SL => n714, Z => n1017);
   U530 : MUXB2DL port map( A0 => n66, A1 => n1409, SL => n715, Z => n1018);
   U532 : MUXB2DL port map( A0 => n66, A1 => n1409, SL => n716, Z => n1019);
   U534 : MUXB2DL port map( A0 => n66, A1 => n1409, SL => n717, Z => n1020);
   U536 : MUXB2DL port map( A0 => n66, A1 => n1409, SL => n718, Z => n1021);
   U538 : MUXB2DL port map( A0 => n66, A1 => n1409, SL => n719, Z => n1022);
   U540 : MUXB2DL port map( A0 => n66, A1 => n1409, SL => n720, Z => n1023);
   U542 : MUXB2DL port map( A0 => n66, A1 => n1409, SL => n721, Z => n1024);
   U544 : MUXB2DL port map( A0 => n66, A1 => n1409, SL => n722, Z => n1025);
   U546 : MUXB2DL port map( A0 => n66, A1 => n1409, SL => n723, Z => n1026);
   U549 : MUXB2DL port map( A0 => n58, A1 => n1407, SL => n724, Z => n1027);
   U551 : MUXB2DL port map( A0 => n58, A1 => n1407, SL => n725, Z => n1028);
   U553 : MUXB2DL port map( A0 => n58, A1 => n1407, SL => n726, Z => n1029);
   U555 : MUXB2DL port map( A0 => n58, A1 => n1407, SL => n727, Z => n1030);
   U557 : MUXB2DL port map( A0 => n58, A1 => n1407, SL => n728, Z => n1031);
   U559 : MUXB2DL port map( A0 => n58, A1 => n1407, SL => n729, Z => n1032);
   U561 : MUXB2DL port map( A0 => n58, A1 => n1407, SL => n730, Z => n1033);
   U563 : MUXB2DL port map( A0 => n58, A1 => n1407, SL => n731, Z => n1034);
   U565 : MUXB2DL port map( A0 => n58, A1 => n1407, SL => n732, Z => n1035);
   U567 : MUXB2DL port map( A0 => n58, A1 => n1407, SL => n733, Z => n1036);
   U569 : MUXB2DL port map( A0 => n58, A1 => n1407, SL => n734, Z => n1037);
   U571 : MUXB2DL port map( A0 => n58, A1 => n1407, SL => n735, Z => n1038);
   U573 : MUXB2DL port map( A0 => n58, A1 => n1407, SL => n736, Z => n1039);
   U575 : MUXB2DL port map( A0 => n58, A1 => n1407, SL => n737, Z => n1040);
   U577 : MUXB2DL port map( A0 => n58, A1 => n1407, SL => n738, Z => n1041);
   U579 : MUXB2DL port map( A0 => n58, A1 => n1407, SL => n739, Z => n1042);
   U581 : MUXB2DL port map( A0 => n58, A1 => n1407, SL => n740, Z => n1043);
   U583 : MUXB2DL port map( A0 => n58, A1 => n1407, SL => n741, Z => n1044);
   U586 : MUXB2DL port map( A0 => n50, A1 => n1405, SL => n742, Z => n1045);
   U588 : MUXB2DL port map( A0 => n50, A1 => n1405, SL => n743, Z => n1046);
   U590 : MUXB2DL port map( A0 => n50, A1 => n1405, SL => n744, Z => n1047);
   U592 : MUXB2DL port map( A0 => n50, A1 => n1405, SL => n745, Z => n1048);
   U594 : MUXB2DL port map( A0 => n50, A1 => n1405, SL => n746, Z => n1049);
   U596 : MUXB2DL port map( A0 => n50, A1 => n1405, SL => n747, Z => n1050);
   U598 : MUXB2DL port map( A0 => n50, A1 => n1405, SL => n748, Z => n1051);
   U600 : MUXB2DL port map( A0 => n50, A1 => n1405, SL => n749, Z => n1052);
   U602 : MUXB2DL port map( A0 => n50, A1 => n1405, SL => n750, Z => n1053);
   U604 : MUXB2DL port map( A0 => n50, A1 => n1405, SL => n751, Z => n1054);
   U606 : MUXB2DL port map( A0 => n50, A1 => n1405, SL => n752, Z => n1055);
   U608 : MUXB2DL port map( A0 => n50, A1 => n1405, SL => n753, Z => n1056);
   U610 : MUXB2DL port map( A0 => n50, A1 => n1405, SL => n754, Z => n1057);
   U612 : MUXB2DL port map( A0 => n50, A1 => n1405, SL => n755, Z => n1058);
   U614 : MUXB2DL port map( A0 => n50, A1 => n1405, SL => n756, Z => n1059);
   U616 : MUXB2DL port map( A0 => n50, A1 => n1405, SL => n757, Z => n1060);
   U618 : MUXB2DL port map( A0 => n50, A1 => n1405, SL => n758, Z => n1061);
   U620 : MUXB2DL port map( A0 => n50, A1 => n1405, SL => n759, Z => n1062);
   U622 : MUXB2DL port map( A0 => n50, A1 => n1405, SL => n760, Z => n1063);
   U624 : MUXB2DL port map( A0 => n50, A1 => n1405, SL => n761, Z => n1064);
   U627 : MUXB2DL port map( A0 => n42, A1 => n1403, SL => n762, Z => n1065);
   U629 : MUXB2DL port map( A0 => n42, A1 => n1403, SL => n763, Z => n1066);
   U631 : MUXB2DL port map( A0 => n42, A1 => n1403, SL => n764, Z => n1067);
   U633 : MUXB2DL port map( A0 => n42, A1 => n1403, SL => n765, Z => n1068);
   U635 : MUXB2DL port map( A0 => n42, A1 => n1403, SL => n766, Z => n1069);
   U637 : MUXB2DL port map( A0 => n42, A1 => n1403, SL => n767, Z => n1070);
   U639 : MUXB2DL port map( A0 => n42, A1 => n1403, SL => n768, Z => n1071);
   U641 : MUXB2DL port map( A0 => n42, A1 => n1403, SL => n769, Z => n1072);
   U643 : MUXB2DL port map( A0 => n42, A1 => n1403, SL => n770, Z => n1073);
   U645 : MUXB2DL port map( A0 => n42, A1 => n1403, SL => n771, Z => n1074);
   U647 : MUXB2DL port map( A0 => n42, A1 => n1403, SL => n772, Z => n1075);
   U649 : MUXB2DL port map( A0 => n42, A1 => n1403, SL => n773, Z => n1076);
   U651 : MUXB2DL port map( A0 => n42, A1 => n1403, SL => n774, Z => n1077);
   U653 : MUXB2DL port map( A0 => n42, A1 => n1403, SL => n775, Z => n1078);
   U655 : MUXB2DL port map( A0 => n42, A1 => n1403, SL => n776, Z => n1079);
   U657 : MUXB2DL port map( A0 => n42, A1 => n1403, SL => n777, Z => n1080);
   U659 : MUXB2DL port map( A0 => n42, A1 => n1403, SL => n778, Z => n1081);
   U661 : MUXB2DL port map( A0 => n42, A1 => n1403, SL => n779, Z => n1082);
   U663 : MUXB2DL port map( A0 => n42, A1 => n1403, SL => n780, Z => n1083);
   U665 : MUXB2DL port map( A0 => n42, A1 => n1403, SL => n781, Z => n1084);
   U667 : MUXB2DL port map( A0 => n42, A1 => n1403, SL => n782, Z => n1085);
   U669 : MUXB2DL port map( A0 => n42, A1 => n1403, SL => n783, Z => n1086);
   U672 : MUXB2DL port map( A0 => n1382, A1 => n1401, SL => n784, Z => n1087);
   U674 : MUXB2DL port map( A0 => n1382, A1 => n1401, SL => n785, Z => n1088);
   U676 : MUXB2DL port map( A0 => n1382, A1 => n1401, SL => n786, Z => n1089);
   U678 : MUXB2DL port map( A0 => n1382, A1 => n1401, SL => n787, Z => n1090);
   U680 : MUXB2DL port map( A0 => n1382, A1 => n1401, SL => n788, Z => n1091);
   U682 : MUXB2DL port map( A0 => n1382, A1 => n1401, SL => n789, Z => n1092);
   U684 : MUXB2DL port map( A0 => n1382, A1 => n1401, SL => n790, Z => n1093);
   U686 : MUXB2DL port map( A0 => n1382, A1 => n1401, SL => n791, Z => n1094);
   U688 : MUXB2DL port map( A0 => n1382, A1 => n1401, SL => n792, Z => n1095);
   U690 : MUXB2DL port map( A0 => n1382, A1 => n1401, SL => n793, Z => n1096);
   U692 : MUXB2DL port map( A0 => n1382, A1 => n1401, SL => n794, Z => n1097);
   U694 : MUXB2DL port map( A0 => n1382, A1 => n1401, SL => n795, Z => n1098);
   U696 : MUXB2DL port map( A0 => n1382, A1 => n1401, SL => n796, Z => n1099);
   U698 : MUXB2DL port map( A0 => n1382, A1 => n1401, SL => n797, Z => n1100);
   U700 : MUXB2DL port map( A0 => n1382, A1 => n1401, SL => n798, Z => n1101);
   U702 : MUXB2DL port map( A0 => n1382, A1 => n1401, SL => n799, Z => n1102);
   U704 : MUXB2DL port map( A0 => n1382, A1 => n1401, SL => n800, Z => n1103);
   U706 : MUXB2DL port map( A0 => n1382, A1 => n1401, SL => n801, Z => n1104);
   U708 : MUXB2DL port map( A0 => n1382, A1 => n1401, SL => n802, Z => n1105);
   U710 : MUXB2DL port map( A0 => n1382, A1 => n1401, SL => n803, Z => n1106);
   U712 : MUXB2DL port map( A0 => n1382, A1 => n1401, SL => n804, Z => n1107);
   U714 : MUXB2DL port map( A0 => n1382, A1 => n1401, SL => n805, Z => n1108);
   U716 : MUXB2DL port map( A0 => n1382, A1 => n1401, SL => n806, Z => n1109);
   U718 : MUXB2DL port map( A0 => n1382, A1 => n1401, SL => n807, Z => n1110);
   U721 : MUXB2DL port map( A0 => n1381, A1 => n1399, SL => n808, Z => n1111);
   U723 : MUXB2DL port map( A0 => n1381, A1 => n1399, SL => n809, Z => n1112);
   U725 : MUXB2DL port map( A0 => n1381, A1 => n1399, SL => n810, Z => n1113);
   U727 : MUXB2DL port map( A0 => n1381, A1 => n1399, SL => n811, Z => n1114);
   U729 : MUXB2DL port map( A0 => n1381, A1 => n1399, SL => n812, Z => n1115);
   U731 : MUXB2DL port map( A0 => n1381, A1 => n1399, SL => n813, Z => n1116);
   U733 : MUXB2DL port map( A0 => n1381, A1 => n1399, SL => n814, Z => n1117);
   U735 : MUXB2DL port map( A0 => n1381, A1 => n1399, SL => n815, Z => n1118);
   U737 : MUXB2DL port map( A0 => n1381, A1 => n1399, SL => n816, Z => n1119);
   U739 : MUXB2DL port map( A0 => n1381, A1 => n1399, SL => n817, Z => n1120);
   U741 : MUXB2DL port map( A0 => n1381, A1 => n1399, SL => n818, Z => n1121);
   U743 : MUXB2DL port map( A0 => n1381, A1 => n1399, SL => n819, Z => n1122);
   U745 : MUXB2DL port map( A0 => n1381, A1 => n1399, SL => n820, Z => n1123);
   U747 : MUXB2DL port map( A0 => n1381, A1 => n1399, SL => n821, Z => n1124);
   U749 : MUXB2DL port map( A0 => n1381, A1 => n1399, SL => n822, Z => n1125);
   U751 : MUXB2DL port map( A0 => n1381, A1 => n1399, SL => n823, Z => n1126);
   U753 : MUXB2DL port map( A0 => n1381, A1 => n1399, SL => n824, Z => n1127);
   U755 : MUXB2DL port map( A0 => n1381, A1 => n1399, SL => n825, Z => n1128);
   U757 : MUXB2DL port map( A0 => n1381, A1 => n1399, SL => n826, Z => n1129);
   U759 : MUXB2DL port map( A0 => n1381, A1 => n1399, SL => n827, Z => n1130);
   U761 : MUXB2DL port map( A0 => n1381, A1 => n1399, SL => n828, Z => n1131);
   U763 : MUXB2DL port map( A0 => n1381, A1 => n1399, SL => n829, Z => n1132);
   U765 : MUXB2DL port map( A0 => n1381, A1 => n1399, SL => n830, Z => n1133);
   U767 : MUXB2DL port map( A0 => n1381, A1 => n1399, SL => n831, Z => n1134);
   U769 : MUXB2DL port map( A0 => n1381, A1 => n1399, SL => n832, Z => n1135);
   U771 : MUXB2DL port map( A0 => n1381, A1 => n1399, SL => n833, Z => n1136);
   U774 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n834, Z => n1137);
   U776 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n835, Z => n1138);
   U778 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n836, Z => n1139);
   U780 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n837, Z => n1140);
   U782 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n838, Z => n1141);
   U784 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n839, Z => n1142);
   U786 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n840, Z => n1143);
   U788 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n841, Z => n1144);
   U790 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n842, Z => n1145);
   U792 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n843, Z => n1146);
   U794 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n844, Z => n1147);
   U796 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n845, Z => n1148);
   U798 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n846, Z => n1149);
   U800 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n847, Z => n1150);
   U802 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n848, Z => n1151);
   U804 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n849, Z => n1152);
   U806 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n850, Z => n1153);
   U808 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n851, Z => n1154);
   U810 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n852, Z => n1155);
   U812 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n853, Z => n1156);
   U814 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n854, Z => n1157);
   U816 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n855, Z => n1158);
   U818 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n856, Z => n1159);
   U820 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n857, Z => n1160);
   U822 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n858, Z => n1161);
   U824 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n859, Z => n1162);
   U826 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n860, Z => n1163);
   U828 : MUXB2DL port map( A0 => n1380, A1 => n1397, SL => n861, Z => n1164);
   U831 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n862, Z => n1165);
   U833 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n863, Z => n1166);
   U835 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n864, Z => n1167);
   U837 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n865, Z => n1168);
   U839 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n866, Z => n1169);
   U841 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n867, Z => n1170);
   U843 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n868, Z => n1171);
   U845 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n869, Z => n1172);
   U847 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n870, Z => n1173);
   U849 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n871, Z => n1174);
   U851 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n872, Z => n1175);
   U853 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n873, Z => n1176);
   U855 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n874, Z => n1177);
   U857 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n875, Z => n1178);
   U859 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n876, Z => n1179);
   U861 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n877, Z => n1180);
   U863 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n878, Z => n1181);
   U865 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n879, Z => n1182);
   U867 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n880, Z => n1183);
   U869 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n881, Z => n1184);
   U871 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n882, Z => n1185);
   U873 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n883, Z => n1186);
   U875 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n884, Z => n1187);
   U877 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n885, Z => n1188);
   U879 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n886, Z => n1189);
   U881 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n887, Z => n1190);
   U883 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n888, Z => n1191);
   U885 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n889, Z => n1192);
   U887 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n890, Z => n1193);
   U889 : MUXB2DL port map( A0 => n1379, A1 => n1396, SL => n891, Z => n1194);
   U892 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n892, Z => n1195);
   U894 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n893, Z => n1196);
   U896 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n894, Z => n1197);
   U898 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n895, Z => n1198);
   U900 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n896, Z => n1199);
   U902 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n897, Z => n1200);
   U904 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n898, Z => n1201);
   U906 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n899, Z => n1202);
   U908 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n900, Z => n1203);
   U910 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n901, Z => n1204);
   U912 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n902, Z => n1205);
   U914 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n903, Z => n1206);
   U916 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n904, Z => n1207);
   U918 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n905, Z => n1208);
   U920 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n906, Z => n1209);
   U922 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n907, Z => n1210);
   U924 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n908, Z => n1211);
   U926 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n909, Z => n1212);
   U928 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n910, Z => n1213);
   U930 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n911, Z => n1214);
   U932 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n912, Z => n1215);
   U934 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n913, Z => n1216);
   U936 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n914, Z => n1217);
   U938 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n915, Z => n1218);
   U940 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n916, Z => n1219);
   U942 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n917, Z => n1220);
   U944 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n918, Z => n1221);
   U946 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n919, Z => n1222);
   U948 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n920, Z => n1223);
   U950 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n921, Z => n1224);
   U952 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n922, Z => n1225);
   U954 : MUXB2DL port map( A0 => n1378, A1 => n1395, SL => n923, Z => n1226);
   U1021 : EXOR2D1 port map( A1 => a(4), A2 => a(3), Z => n1375);
   U1022 : EXOR2D1 port map( A1 => a(6), A2 => a(5), Z => n1376);
   U1023 : EXOR2D1 port map( A1 => a(8), A2 => a(7), Z => n1377);
   U1024 : NAN2D1 port map( A1 => a(0), A2 => n1395, Z => n1378);
   U1025 : OAI21D1 port map( A1 => a(2), A2 => a(1), B => n1398, Z => n1379);
   U1026 : OAI21D1 port map( A1 => a(4), A2 => a(3), B => n1400, Z => n1380);
   U1027 : OAI21D1 port map( A1 => a(6), A2 => a(5), B => n1402, Z => n1381);
   U1028 : OAI21D1 port map( A1 => a(8), A2 => a(7), B => n1404, Z => n1382);
   U1029 : INVD1 port map( A => n1383, Z => n1384);
   U1030 : INVD1 port map( A => n1390, Z => n1389);
   U1031 : INVD1 port map( A => n1392, Z => n1391);
   U1032 : INVD1 port map( A => n1394, Z => n1393);
   U1033 : INVD1 port map( A => n1388, Z => n1387);
   U1034 : INVD1 port map( A => n953, Z => n1396);
   U1035 : INVD1 port map( A => n1386, Z => n1385);
   U1036 : INVD1 port map( A => n952, Z => n1397);
   U1037 : INVD1 port map( A => n951, Z => n1399);
   U1038 : INVD1 port map( A => n950, Z => n1401);
   U1039 : INVD1 port map( A => n949, Z => n1403);
   U1040 : INVD1 port map( A => n948, Z => n1405);
   U1041 : INVD1 port map( A => n947, Z => n1407);
   U1042 : INVD1 port map( A => n946, Z => n1409);
   U1043 : INVD1 port map( A => n945, Z => n1411);
   U1044 : INVD1 port map( A => n944, Z => n1413);
   U1045 : INVD1 port map( A => n943, Z => n1415);
   U1046 : INVD1 port map( A => n942, Z => n1417);
   U1047 : INVD1 port map( A => n941, Z => n1419);
   U1048 : INVD1 port map( A => n940, Z => n1422);
   U1049 : INVD1 port map( A => n939, Z => n1423);
   U1050 : INVD1 port map( A => a(1), Z => n1395);
   U1051 : EXNOR2D1 port map( A1 => a(2), A2 => a(1), Z => n1383);
   U1052 : INVD1 port map( A => b(2), Z => n1390);
   U1053 : INVD1 port map( A => b(1), Z => n1392);
   U1054 : INVD1 port map( A => b(0), Z => n1394);
   U1055 : INVD1 port map( A => b(3), Z => n1388);
   U1056 : INVD1 port map( A => a(3), Z => n1398);
   U1057 : INVD1 port map( A => a(5), Z => n1400);
   U1058 : INVD1 port map( A => b(5), Z => n1386);
   U1059 : INVD1 port map( A => a(7), Z => n1402);
   U1060 : INVD1 port map( A => a(9), Z => n1404);
   U1061 : EXOR2D1 port map( A1 => a(10), A2 => a(9), Z => n1444);
   U1062 : INVD1 port map( A => a(11), Z => n1406);
   U1063 : OAI21D1 port map( A1 => a(9), A2 => a(10), B => n1406, Z => n42);
   U1064 : EXOR2D1 port map( A1 => a(12), A2 => a(11), Z => n1445);
   U1065 : INVD1 port map( A => a(13), Z => n1408);
   U1066 : OAI21D1 port map( A1 => a(12), A2 => a(11), B => n1408, Z => n50);
   U1067 : EXOR2D1 port map( A1 => a(14), A2 => a(13), Z => n1446);
   U1068 : INVD1 port map( A => a(15), Z => n1410);
   U1069 : OAI21D1 port map( A1 => a(14), A2 => a(13), B => n1410, Z => n58);
   U1070 : EXOR2D1 port map( A1 => a(16), A2 => a(15), Z => n1447);
   U1071 : INVD1 port map( A => a(17), Z => n1412);
   U1072 : OAI21D1 port map( A1 => a(16), A2 => a(15), B => n1412, Z => n66);
   U1073 : EXOR2D1 port map( A1 => a(18), A2 => a(17), Z => n1448);
   U1074 : INVD1 port map( A => a(19), Z => n1414);
   U1075 : OAI21D1 port map( A1 => a(18), A2 => a(17), B => n1414, Z => n73);
   U1076 : EXOR2D1 port map( A1 => a(20), A2 => a(19), Z => n1449);
   U1077 : INVD1 port map( A => a(21), Z => n1416);
   U1078 : OAI21D1 port map( A1 => a(20), A2 => a(19), B => n1416, Z => n80);
   U1079 : EXOR2D1 port map( A1 => a(22), A2 => a(21), Z => n1450);
   U1080 : INVD1 port map( A => a(23), Z => n1418);
   U1081 : OAI21D1 port map( A1 => a(22), A2 => a(21), B => n1418, Z => n84);
   U1082 : INVD1 port map( A => a(25), Z => n1420);
   U1083 : INVD1 port map( A => a(27), Z => n1421);
   U1084 : INVD1 port map( A => a(29), Z => n1424);
   U1085 : MUXB2DL port map( A0 => b(29), A1 => b(28), SL => n1383, Z => n862);
   U1086 : INVD1 port map( A => a(31), Z => n1425);
   U1087 : EXOR3D1 port map( A1 => n1426, A2 => n1427, A3 => n1428, Z => 
                           product(31));
   U1088 : EXOR3D1 port map( A1 => n208, A2 => n206, A3 => n1429, Z => n1428);
   U1089 : EXOR2D1 port map( A1 => n214, A2 => n212, Z => n1429);
   U1090 : EXOR2D1 port map( A1 => n202, A2 => n156, Z => n1427);
   U1091 : EXOR3D1 port map( A1 => n1430, A2 => n1431, A3 => n1432, Z => n1426)
                           ;
   U1092 : EXOR3D1 port map( A1 => n957, A2 => n955, A3 => n1433, Z => n1432);
   U1093 : EXNOR2D1 port map( A1 => n997, A2 => n975, Z => n1433);
   U1094 : EXOR3D1 port map( A1 => n1434, A2 => n204, A3 => n1435, Z => n1431);
   U1095 : EXOR3D1 port map( A1 => n1087, A2 => n1065, A3 => n1436, Z => n1435)
                           ;
   U1096 : EXNOR2D1 port map( A1 => n210, A2 => n1111, Z => n1436);
   U1097 : EXOR3D1 port map( A1 => n961, A2 => n218, A3 => n1437, Z => n1434);
   U1098 : EXOR2D1 port map( A1 => n985, A2 => n967, Z => n1437);
   U1099 : EXOR3D1 port map( A1 => n1438, A2 => n1439, A3 => n1440, Z => n1430)
                           ;
   U1100 : EXOR3D1 port map( A1 => n1027, A2 => n1011, A3 => n1441, Z => n1440)
                           ;
   U1101 : EXOR3D1 port map( A1 => n1165, A2 => n1137, A3 => n1045, Z => n1441)
                           ;
   U1102 : EXOR3D1 port map( A1 => n216, A2 => n1195, A3 => n1442, Z => n1439);
   U1103 : EXOR2D1 port map( A1 => n222, A2 => n220, Z => n1442);
   U1104 : EXOR3D1 port map( A1 => n226, A2 => n224, A3 => n1443, Z => n1438);
   U1105 : EXOR2D1 port map( A1 => n230, A2 => n228, Z => n1443);
   U1106 : OAI21D1 port map( A1 => a(28), A2 => a(27), B => n1424, Z => n99);
   U1107 : AOI21D1 port map( A1 => a(25), A2 => a(26), B => n1421, Z => n941);
   U1108 : OAI21D1 port map( A1 => a(26), A2 => a(25), B => n1421, Z => n94);
   U1109 : NAN2D1 port map( A1 => n1393, A2 => a(0), Z => n923);
   U1110 : MUXB2DL port map( A0 => b(0), A1 => n1391, SL => a(0), Z => n922);
   U1111 : MUXB2DL port map( A0 => n1391, A1 => n1389, SL => a(0), Z => n921);
   U1112 : MUXB2DL port map( A0 => b(2), A1 => n1387, SL => a(0), Z => n920);
   U1113 : MUXB2DL port map( A0 => n1387, A1 => b(4), SL => a(0), Z => n919);
   U1114 : MUXB2DL port map( A0 => b(4), A1 => n1385, SL => a(0), Z => n918);
   U1115 : MUXB2DL port map( A0 => n1385, A1 => b(6), SL => a(0), Z => n917);
   U1116 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => a(0), Z => n916);
   U1117 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => a(0), Z => n915);
   U1118 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => a(0), Z => n914);
   U1119 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => a(0), Z => n913);
   U1120 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => a(0), Z => n912);
   U1121 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => a(0), Z => n911);
   U1122 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => a(0), Z => n910);
   U1123 : AOI21D1 port map( A1 => a(23), A2 => a(24), B => n1420, Z => n942);
   U1124 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => a(0), Z => n909);
   U1125 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => a(0), Z => n908);
   U1126 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => a(0), Z => n907);
   U1127 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => a(0), Z => n906);
   U1128 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => a(0), Z => n905);
   U1129 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => a(0), Z => n904);
   U1130 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => a(0), Z => n903);
   U1131 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => a(0), Z => n902);
   U1132 : MUXB2DL port map( A0 => b(21), A1 => b(22), SL => a(0), Z => n901);
   U1133 : MUXB2DL port map( A0 => b(22), A1 => b(23), SL => a(0), Z => n900);
   U1134 : MUXB2DL port map( A0 => b(23), A1 => b(24), SL => a(0), Z => n899);
   U1135 : MUXB2DL port map( A0 => b(24), A1 => b(25), SL => a(0), Z => n898);
   U1136 : MUXB2DL port map( A0 => b(25), A1 => b(26), SL => a(0), Z => n897);
   U1137 : MUXB2DL port map( A0 => b(26), A1 => b(27), SL => a(0), Z => n896);
   U1138 : MUXB2DL port map( A0 => b(27), A1 => b(28), SL => a(0), Z => n895);
   U1139 : MUXB2DL port map( A0 => b(28), A1 => b(29), SL => a(0), Z => n894);
   U1140 : MUXB2DL port map( A0 => b(29), A1 => b(30), SL => a(0), Z => n893);
   U1141 : MUXB2DL port map( A0 => b(30), A1 => b(31), SL => a(0), Z => n892);
   U1142 : NAN2D1 port map( A1 => n1393, A2 => n1384, Z => n891);
   U1143 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1384, Z => n890);
   U1144 : OAI21D1 port map( A1 => a(24), A2 => a(23), B => n1420, Z => n89);
   U1145 : MUXB2DL port map( A0 => n1391, A1 => n1389, SL => n1384, Z => n889);
   U1146 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1384, Z => n888);
   U1147 : MUXB2DL port map( A0 => n1387, A1 => b(4), SL => n1384, Z => n887);
   U1148 : MUXB2DL port map( A0 => b(4), A1 => n1385, SL => n1384, Z => n886);
   U1149 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1384, Z => n885);
   U1150 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1384, Z => n884);
   U1151 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1384, Z => n883);
   U1152 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1384, Z => n882);
   U1153 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1384, Z => n881);
   U1154 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1384, Z => n880);
   U1155 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1384, Z => n879);
   U1156 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1384, Z => n878);
   U1157 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1384, Z => n877);
   U1158 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1384, Z => n876);
   U1159 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1384, Z => n875);
   U1160 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1384, Z => n874);
   U1161 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1384, Z => n873);
   U1162 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1384, Z => n872);
   U1163 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => n1384, Z => n871);
   U1164 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => n1384, Z => n870);
   U1165 : MUXB2DL port map( A0 => b(21), A1 => b(22), SL => n1384, Z => n869);
   U1166 : MUXB2DL port map( A0 => b(22), A1 => b(23), SL => n1384, Z => n868);
   U1167 : MUXB2DL port map( A0 => b(23), A1 => b(24), SL => n1384, Z => n867);
   U1168 : MUXB2DL port map( A0 => b(24), A1 => b(25), SL => n1384, Z => n866);
   U1169 : MUXB2DL port map( A0 => b(25), A1 => b(26), SL => n1384, Z => n865);
   U1170 : MUXB2DL port map( A0 => b(26), A1 => b(27), SL => n1384, Z => n864);
   U1171 : MUXB2DL port map( A0 => b(27), A1 => b(28), SL => n1384, Z => n863);
   U1172 : NAN2D1 port map( A1 => n1393, A2 => n1375, Z => n861);
   U1173 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1375, Z => n860);
   U1174 : AOI21D1 port map( A1 => a(21), A2 => a(22), B => n1418, Z => n943);
   U1175 : MUXB2DL port map( A0 => n1391, A1 => n1389, SL => n1375, Z => n859);
   U1176 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1375, Z => n858);
   U1177 : MUXB2DL port map( A0 => n1387, A1 => b(4), SL => n1375, Z => n857);
   U1178 : MUXB2DL port map( A0 => b(4), A1 => n1385, SL => n1375, Z => n856);
   U1179 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1375, Z => n855);
   U1180 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1375, Z => n854);
   U1181 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1375, Z => n853);
   U1182 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1375, Z => n852);
   U1183 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1375, Z => n851);
   U1184 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1375, Z => n850);
   U1185 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1375, Z => n849);
   U1186 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1375, Z => n848);
   U1187 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1375, Z => n847);
   U1188 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1375, Z => n846);
   U1189 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1375, Z => n845);
   U1190 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1375, Z => n844);
   U1191 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1375, Z => n843);
   U1192 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1375, Z => n842);
   U1193 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => n1375, Z => n841);
   U1194 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => n1375, Z => n840);
   U1195 : MUXB2DL port map( A0 => b(21), A1 => b(22), SL => n1375, Z => n839);
   U1196 : MUXB2DL port map( A0 => b(22), A1 => b(23), SL => n1375, Z => n838);
   U1197 : MUXB2DL port map( A0 => b(23), A1 => b(24), SL => n1375, Z => n837);
   U1198 : MUXB2DL port map( A0 => b(24), A1 => b(25), SL => n1375, Z => n836);
   U1199 : MUXB2DL port map( A0 => b(25), A1 => b(26), SL => n1375, Z => n835);
   U1200 : MUXB2DL port map( A0 => b(26), A1 => b(27), SL => n1375, Z => n834);
   U1201 : NAN2D1 port map( A1 => n1393, A2 => n1376, Z => n833);
   U1202 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1376, Z => n832);
   U1203 : MUXB2DL port map( A0 => n1391, A1 => n1389, SL => n1376, Z => n831);
   U1204 : MUXB2DL port map( A0 => n1389, A1 => b(3), SL => n1376, Z => n830);
   U1205 : MUXB2DL port map( A0 => n1387, A1 => b(4), SL => n1376, Z => n829);
   U1206 : MUXB2DL port map( A0 => b(4), A1 => n1385, SL => n1376, Z => n828);
   U1207 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1376, Z => n827);
   U1208 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1376, Z => n826);
   U1209 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1376, Z => n825);
   U1210 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1376, Z => n824);
   U1211 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1376, Z => n823);
   U1212 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1376, Z => n822);
   U1213 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1376, Z => n821);
   U1214 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1376, Z => n820);
   U1215 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1376, Z => n819);
   U1216 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1376, Z => n818);
   U1217 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1376, Z => n817);
   U1218 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1376, Z => n816);
   U1219 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1376, Z => n815);
   U1220 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1376, Z => n814);
   U1221 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => n1376, Z => n813);
   U1222 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => n1376, Z => n812);
   U1223 : MUXB2DL port map( A0 => b(21), A1 => b(22), SL => n1376, Z => n811);
   U1224 : MUXB2DL port map( A0 => b(22), A1 => b(23), SL => n1376, Z => n810);
   U1225 : AOI21D1 port map( A1 => a(19), A2 => a(20), B => n1416, Z => n944);
   U1226 : MUXB2DL port map( A0 => b(23), A1 => b(24), SL => n1376, Z => n809);
   U1227 : MUXB2DL port map( A0 => b(24), A1 => b(25), SL => n1376, Z => n808);
   U1228 : NAN2D1 port map( A1 => n1393, A2 => n1377, Z => n807);
   U1229 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1377, Z => n806);
   U1230 : MUXB2DL port map( A0 => b(1), A1 => n1389, SL => n1377, Z => n805);
   U1231 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1377, Z => n804);
   U1232 : MUXB2DL port map( A0 => n1387, A1 => b(4), SL => n1377, Z => n803);
   U1233 : MUXB2DL port map( A0 => b(4), A1 => n1385, SL => n1377, Z => n802);
   U1234 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1377, Z => n801);
   U1235 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1377, Z => n800);
   U1236 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1377, Z => n799);
   U1237 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1377, Z => n798);
   U1238 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1377, Z => n797);
   U1239 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1377, Z => n796);
   U1240 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1377, Z => n795);
   U1241 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1377, Z => n794);
   U1242 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1377, Z => n793);
   U1243 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1377, Z => n792);
   U1244 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1377, Z => n791);
   U1245 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1377, Z => n790);
   U1246 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1377, Z => n789);
   U1247 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1377, Z => n788);
   U1248 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => n1377, Z => n787);
   U1249 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => n1377, Z => n786);
   U1250 : MUXB2DL port map( A0 => b(21), A1 => b(22), SL => n1377, Z => n785);
   U1251 : MUXB2DL port map( A0 => b(22), A1 => b(23), SL => n1377, Z => n784);
   U1252 : NAN2D1 port map( A1 => n1393, A2 => n1444, Z => n783);
   U1253 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1444, Z => n782);
   U1254 : MUXB2DL port map( A0 => n1391, A1 => n1389, SL => n1444, Z => n781);
   U1255 : MUXB2DL port map( A0 => n1389, A1 => b(3), SL => n1444, Z => n780);
   U1256 : MUXB2DL port map( A0 => b(3), A1 => b(4), SL => n1444, Z => n779);
   U1257 : MUXB2DL port map( A0 => b(4), A1 => n1385, SL => n1444, Z => n778);
   U1258 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1444, Z => n777);
   U1259 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1444, Z => n776);
   U1260 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1444, Z => n775);
   U1261 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1444, Z => n774);
   U1262 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1444, Z => n773);
   U1263 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1444, Z => n772);
   U1264 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1444, Z => n771);
   U1265 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1444, Z => n770);
   U1266 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1444, Z => n769);
   U1267 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1444, Z => n768);
   U1268 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1444, Z => n767);
   U1269 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1444, Z => n766);
   U1270 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1444, Z => n765);
   U1271 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1444, Z => n764);
   U1272 : MUXB2DL port map( A0 => b(19), A1 => b(20), SL => n1444, Z => n763);
   U1273 : MUXB2DL port map( A0 => b(20), A1 => b(21), SL => n1444, Z => n762);
   U1274 : NAN2D1 port map( A1 => n1393, A2 => n1445, Z => n761);
   U1275 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1445, Z => n760);
   U1276 : MUXB2DL port map( A0 => b(1), A1 => n1389, SL => n1445, Z => n759);
   U1277 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1445, Z => n758);
   U1278 : MUXB2DL port map( A0 => n1387, A1 => b(4), SL => n1445, Z => n757);
   U1279 : MUXB2DL port map( A0 => b(4), A1 => n1385, SL => n1445, Z => n756);
   U1280 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1445, Z => n755);
   U1281 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1445, Z => n754);
   U1282 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1445, Z => n753);
   U1283 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1445, Z => n752);
   U1284 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1445, Z => n751);
   U1285 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1445, Z => n750);
   U1286 : AOI21D1 port map( A1 => a(17), A2 => a(18), B => n1414, Z => n945);
   U1287 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1445, Z => n749);
   U1288 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1445, Z => n748);
   U1289 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1445, Z => n747);
   U1290 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1445, Z => n746);
   U1291 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1445, Z => n745);
   U1292 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1445, Z => n744);
   U1293 : MUXB2DL port map( A0 => b(17), A1 => b(18), SL => n1445, Z => n743);
   U1294 : MUXB2DL port map( A0 => b(18), A1 => b(19), SL => n1445, Z => n742);
   U1295 : NAN2D1 port map( A1 => n1393, A2 => n1446, Z => n741);
   U1296 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1446, Z => n740);
   U1297 : MUXB2DL port map( A0 => n1391, A1 => n1389, SL => n1446, Z => n739);
   U1298 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1446, Z => n738);
   U1299 : MUXB2DL port map( A0 => n1387, A1 => b(4), SL => n1446, Z => n737);
   U1300 : MUXB2DL port map( A0 => b(4), A1 => n1385, SL => n1446, Z => n736);
   U1301 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1446, Z => n735);
   U1302 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1446, Z => n734);
   U1303 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1446, Z => n733);
   U1304 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1446, Z => n732);
   U1305 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1446, Z => n731);
   U1306 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1446, Z => n730);
   U1307 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1446, Z => n729);
   U1308 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1446, Z => n728);
   U1309 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1446, Z => n727);
   U1310 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1446, Z => n726);
   U1311 : MUXB2DL port map( A0 => b(15), A1 => b(16), SL => n1446, Z => n725);
   U1312 : MUXB2DL port map( A0 => b(16), A1 => b(17), SL => n1446, Z => n724);
   U1313 : NAN2D1 port map( A1 => n1393, A2 => n1447, Z => n723);
   U1314 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1447, Z => n722);
   U1315 : MUXB2DL port map( A0 => n1391, A1 => n1389, SL => n1447, Z => n721);
   U1316 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1447, Z => n720);
   U1317 : MUXB2DL port map( A0 => n1387, A1 => b(4), SL => n1447, Z => n719);
   U1318 : MUXB2DL port map( A0 => b(4), A1 => n1385, SL => n1447, Z => n718);
   U1319 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1447, Z => n717);
   U1320 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1447, Z => n716);
   U1321 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1447, Z => n715);
   U1322 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1447, Z => n714);
   U1323 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1447, Z => n713);
   U1324 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1447, Z => n712);
   U1325 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1447, Z => n711);
   U1326 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1447, Z => n710);
   U1327 : MUXB2DL port map( A0 => b(13), A1 => b(14), SL => n1447, Z => n709);
   U1328 : MUXB2DL port map( A0 => b(14), A1 => b(15), SL => n1447, Z => n708);
   U1329 : NAN2D1 port map( A1 => n1393, A2 => n1448, Z => n707);
   U1330 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1448, Z => n706);
   U1331 : MUXB2DL port map( A0 => n1391, A1 => n1389, SL => n1448, Z => n705);
   U1332 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1448, Z => n704);
   U1333 : MUXB2DL port map( A0 => n1387, A1 => b(4), SL => n1448, Z => n703);
   U1334 : MUXB2DL port map( A0 => b(4), A1 => n1385, SL => n1448, Z => n702);
   U1335 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1448, Z => n701);
   U1336 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1448, Z => n700);
   U1337 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1448, Z => n699);
   U1338 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1448, Z => n698);
   U1339 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1448, Z => n697);
   U1340 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1448, Z => n696);
   U1341 : MUXB2DL port map( A0 => b(11), A1 => b(12), SL => n1448, Z => n695);
   U1342 : MUXB2DL port map( A0 => b(12), A1 => b(13), SL => n1448, Z => n694);
   U1343 : NAN2D1 port map( A1 => n1393, A2 => n1449, Z => n693);
   U1344 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1449, Z => n692);
   U1345 : MUXB2DL port map( A0 => n1391, A1 => b(2), SL => n1449, Z => n691);
   U1346 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1449, Z => n690);
   U1347 : MUXB2DL port map( A0 => n1387, A1 => b(4), SL => n1449, Z => n689);
   U1348 : MUXB2DL port map( A0 => b(4), A1 => n1385, SL => n1449, Z => n688);
   U1349 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1449, Z => n687);
   U1350 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1449, Z => n686);
   U1351 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1449, Z => n685);
   U1352 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1449, Z => n684);
   U1353 : MUXB2DL port map( A0 => b(9), A1 => b(10), SL => n1449, Z => n683);
   U1354 : MUXB2DL port map( A0 => b(10), A1 => b(11), SL => n1449, Z => n682);
   U1355 : NAN2D1 port map( A1 => n1393, A2 => n1450, Z => n681);
   U1356 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1450, Z => n680);
   U1357 : AOI21D1 port map( A1 => a(15), A2 => a(16), B => n1412, Z => n946);
   U1358 : MUXB2DL port map( A0 => n1391, A1 => b(2), SL => n1450, Z => n679);
   U1359 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1450, Z => n678);
   U1360 : MUXB2DL port map( A0 => n1387, A1 => b(4), SL => n1450, Z => n677);
   U1361 : MUXB2DL port map( A0 => b(4), A1 => n1385, SL => n1450, Z => n676);
   U1362 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1450, Z => n675);
   U1363 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1450, Z => n674);
   U1364 : MUXB2DL port map( A0 => b(7), A1 => b(8), SL => n1450, Z => n673);
   U1365 : MUXB2DL port map( A0 => b(8), A1 => b(9), SL => n1450, Z => n672);
   U1366 : NAN2D1 port map( A1 => b(0), A2 => n1451, Z => n671);
   U1367 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1451, Z => n670);
   U1368 : MUXB2DL port map( A0 => n1391, A1 => b(2), SL => n1451, Z => n669);
   U1369 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1451, Z => n668);
   U1370 : MUXB2DL port map( A0 => n1387, A1 => b(4), SL => n1451, Z => n667);
   U1371 : MUXB2DL port map( A0 => b(4), A1 => b(5), SL => n1451, Z => n666);
   U1372 : MUXB2DL port map( A0 => b(5), A1 => b(6), SL => n1451, Z => n665);
   U1373 : MUXB2DL port map( A0 => b(6), A1 => b(7), SL => n1451, Z => n664);
   U1374 : EXOR2D1 port map( A1 => a(24), A2 => a(23), Z => n1451);
   U1375 : NAN2D1 port map( A1 => b(0), A2 => n1452, Z => n663);
   U1376 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1452, Z => n662);
   U1377 : MUXB2DL port map( A0 => n1391, A1 => b(2), SL => n1452, Z => n661);
   U1378 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1452, Z => n660);
   U1379 : MUXB2DL port map( A0 => n1387, A1 => b(4), SL => n1452, Z => n659);
   U1380 : MUXB2DL port map( A0 => b(4), A1 => n1385, SL => n1452, Z => n658);
   U1381 : EXOR2D1 port map( A1 => a(26), A2 => a(25), Z => n1452);
   U1382 : NAN2D1 port map( A1 => b(0), A2 => n1453, Z => n657);
   U1383 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1453, Z => n656);
   U1384 : MUXB2DL port map( A0 => n1391, A1 => n1389, SL => n1453, Z => n655);
   U1385 : MUXB2DL port map( A0 => b(2), A1 => b(3), SL => n1453, Z => n654);
   U1386 : EXOR2D1 port map( A1 => a(28), A2 => a(27), Z => n1453);
   U1387 : NAN2D1 port map( A1 => b(0), A2 => n1454, Z => n653);
   U1388 : MUXB2DL port map( A0 => b(0), A1 => b(1), SL => n1454, Z => n652);
   U1389 : EXOR2D1 port map( A1 => a(30), A2 => a(29), Z => n1454);
   U1390 : AOI21D1 port map( A1 => a(13), A2 => a(14), B => n1410, Z => n947);
   U1391 : AOI21D1 port map( A1 => a(11), A2 => a(12), B => n1408, Z => n948);
   U1392 : AOI21D1 port map( A1 => a(9), A2 => a(10), B => n1406, Z => n949);
   U1393 : AOI21D1 port map( A1 => a(7), A2 => a(8), B => n1404, Z => n950);
   U1394 : AOI21D1 port map( A1 => a(5), A2 => a(6), B => n1402, Z => n951);
   U1395 : AOI21D1 port map( A1 => a(3), A2 => a(4), B => n1400, Z => n952);
   U1396 : AOI21D1 port map( A1 => a(1), A2 => a(2), B => n1398, Z => n953);
   U1397 : AOI21D1 port map( A1 => a(29), A2 => a(30), B => n1425, Z => n939);
   U1398 : OAI21D1 port map( A1 => a(30), A2 => a(29), B => n1425, Z => n104);
   U1399 : AOI21D1 port map( A1 => a(27), A2 => a(28), B => n1424, Z => n940);

end hier_filter_none_20;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_gp_custom.all;

architecture hier_filter_none_20 of gp_custom is

   component NOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN4D1
      port( A1, A2, A3, A4 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AO22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AO31D1
      port( A1, A2, A3, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22M10D1
      port( B1, B2, A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3M1D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211D1
      port( A1, A2, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFBD2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFRPQ1
      port( D, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component DFERPQ1
      port( D, CEB, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFSPQ1
      port( D, CK, SB : in std_logic;  Q : out std_logic);
   end component;
   
   component gp_custom_DW_mult_tc_0
      port( a, b : in std_logic_vector (31 downto 0);  product : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component gp_custom_DW_mult_tc_1
      port( a, b : in std_logic_vector (31 downto 0);  product : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component gp_custom_DW_mult_tc_4
      port( a, b : in std_logic_vector (31 downto 0);  product : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component gp_custom_DW_mult_tc_3
      port( a, b : in std_logic_vector (31 downto 0);  product : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component gp_custom_DW_mult_tc_2
      port( a, b : in std_logic_vector (31 downto 0);  product : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component OA21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI32D1
      port( A1, A2, A3, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal N62, N63, N64, avs_readdata_31_port, avs_readdata_30_port, 
      avs_readdata_29_port, avs_readdata_28_port, avs_readdata_27_port, 
      avs_readdata_26_port, avs_readdata_25_port, avs_readdata_24_port, 
      avs_readdata_23_port, avs_readdata_22_port, avs_readdata_21_port, 
      avs_readdata_20_port, avs_readdata_19_port, avs_readdata_18_port, 
      avs_readdata_17_port, avs_readdata_16_port, avs_readdata_15_port, 
      avs_readdata_14_port, avs_readdata_13_port, avs_readdata_12_port, 
      avs_readdata_11_port, avs_readdata_10_port, avs_readdata_9_port, 
      avs_readdata_8_port, avs_readdata_7_port, avs_readdata_6_port, 
      avs_readdata_5_port, avs_readdata_4_port, avs_readdata_3_port, 
      avs_readdata_2_port, avs_readdata_1_port, avs_readdata_0_port, 
      stop_sim_port, out_buf_255_port, out_buf_254_port, out_buf_253_port, 
      out_buf_252_port, out_buf_251_port, out_buf_250_port, out_buf_249_port, 
      out_buf_248_port, out_buf_247_port, out_buf_246_port, out_buf_245_port, 
      out_buf_244_port, out_buf_243_port, out_buf_242_port, out_buf_241_port, 
      out_buf_240_port, out_buf_239_port, out_buf_238_port, out_buf_237_port, 
      out_buf_236_port, out_buf_235_port, out_buf_234_port, out_buf_233_port, 
      out_buf_232_port, out_buf_231_port, out_buf_230_port, out_buf_229_port, 
      out_buf_228_port, out_buf_227_port, out_buf_226_port, out_buf_225_port, 
      out_buf_224_port, out_buf_223_port, out_buf_222_port, out_buf_221_port, 
      out_buf_220_port, out_buf_219_port, out_buf_218_port, out_buf_217_port, 
      out_buf_216_port, out_buf_215_port, out_buf_214_port, out_buf_213_port, 
      out_buf_212_port, out_buf_211_port, out_buf_210_port, out_buf_209_port, 
      out_buf_208_port, out_buf_207_port, out_buf_206_port, out_buf_205_port, 
      out_buf_204_port, out_buf_203_port, out_buf_202_port, out_buf_201_port, 
      out_buf_200_port, out_buf_199_port, out_buf_198_port, out_buf_197_port, 
      out_buf_196_port, out_buf_195_port, out_buf_194_port, out_buf_193_port, 
      out_buf_192_port, out_buf_191_port, out_buf_190_port, out_buf_189_port, 
      out_buf_188_port, out_buf_187_port, out_buf_186_port, out_buf_185_port, 
      out_buf_184_port, out_buf_183_port, out_buf_182_port, out_buf_181_port, 
      out_buf_180_port, out_buf_179_port, out_buf_178_port, out_buf_177_port, 
      out_buf_176_port, out_buf_175_port, out_buf_174_port, out_buf_173_port, 
      out_buf_172_port, out_buf_171_port, out_buf_170_port, out_buf_169_port, 
      out_buf_168_port, out_buf_167_port, out_buf_166_port, out_buf_165_port, 
      out_buf_164_port, out_buf_163_port, out_buf_162_port, out_buf_161_port, 
      out_buf_160_port, out_buf_159_port, out_buf_158_port, out_buf_157_port, 
      out_buf_156_port, out_buf_155_port, out_buf_154_port, out_buf_153_port, 
      out_buf_152_port, out_buf_151_port, out_buf_150_port, out_buf_149_port, 
      out_buf_148_port, out_buf_147_port, out_buf_146_port, out_buf_145_port, 
      out_buf_144_port, out_buf_143_port, out_buf_142_port, out_buf_141_port, 
      out_buf_140_port, out_buf_139_port, out_buf_138_port, out_buf_137_port, 
      out_buf_136_port, out_buf_135_port, out_buf_134_port, out_buf_133_port, 
      out_buf_132_port, out_buf_131_port, out_buf_130_port, out_buf_129_port, 
      out_buf_128_port, out_buf_127_port, out_buf_126_port, out_buf_125_port, 
      out_buf_124_port, out_buf_123_port, out_buf_122_port, out_buf_121_port, 
      out_buf_120_port, out_buf_119_port, out_buf_118_port, out_buf_117_port, 
      out_buf_116_port, out_buf_115_port, out_buf_114_port, out_buf_113_port, 
      out_buf_112_port, out_buf_111_port, out_buf_110_port, out_buf_109_port, 
      out_buf_108_port, out_buf_107_port, out_buf_106_port, out_buf_105_port, 
      out_buf_104_port, out_buf_103_port, out_buf_102_port, out_buf_101_port, 
      out_buf_100_port, out_buf_99_port, out_buf_98_port, out_buf_97_port, 
      out_buf_96_port, out_buf_95_port, out_buf_94_port, out_buf_93_port, 
      out_buf_92_port, out_buf_91_port, out_buf_90_port, out_buf_89_port, 
      out_buf_88_port, out_buf_87_port, out_buf_86_port, out_buf_85_port, 
      out_buf_84_port, out_buf_83_port, out_buf_82_port, out_buf_81_port, 
      out_buf_80_port, out_buf_79_port, out_buf_78_port, out_buf_77_port, 
      out_buf_76_port, out_buf_75_port, out_buf_74_port, out_buf_73_port, 
      out_buf_72_port, out_buf_71_port, out_buf_70_port, out_buf_69_port, 
      out_buf_68_port, out_buf_67_port, out_buf_66_port, out_buf_65_port, 
      out_buf_64_port, out_buf_63_port, out_buf_62_port, out_buf_61_port, 
      out_buf_60_port, out_buf_59_port, out_buf_58_port, out_buf_57_port, 
      out_buf_56_port, out_buf_55_port, out_buf_54_port, out_buf_53_port, 
      out_buf_52_port, out_buf_51_port, out_buf_50_port, out_buf_49_port, 
      out_buf_48_port, out_buf_47_port, out_buf_46_port, out_buf_45_port, 
      out_buf_44_port, out_buf_43_port, out_buf_42_port, out_buf_41_port, 
      out_buf_40_port, out_buf_39_port, out_buf_38_port, out_buf_37_port, 
      out_buf_36_port, out_buf_35_port, out_buf_34_port, out_buf_33_port, 
      out_buf_32_port, out_buf_31_port, out_buf_30_port, out_buf_29_port, 
      out_buf_28_port, out_buf_27_port, out_buf_26_port, out_buf_25_port, 
      out_buf_24_port, out_buf_23_port, out_buf_22_port, out_buf_21_port, 
      out_buf_20_port, out_buf_19_port, out_buf_18_port, out_buf_17_port, 
      out_buf_16_port, out_buf_15_port, out_buf_14_port, out_buf_13_port, 
      out_buf_12_port, out_buf_11_port, out_buf_10_port, out_buf_9_port, 
      out_buf_8_port, out_buf_7_port, out_buf_6_port, out_buf_5_port, 
      out_buf_4_port, out_buf_3_port, out_buf_2_port, out_buf_1_port, 
      out_buf_0_port, coeff_memory_0_31_port, coeff_memory_0_30_port, 
      coeff_memory_0_29_port, coeff_memory_0_28_port, coeff_memory_0_27_port, 
      coeff_memory_0_26_port, coeff_memory_0_25_port, coeff_memory_0_24_port, 
      coeff_memory_0_23_port, coeff_memory_0_22_port, coeff_memory_0_21_port, 
      coeff_memory_0_20_port, coeff_memory_0_19_port, coeff_memory_0_18_port, 
      coeff_memory_0_17_port, coeff_memory_0_16_port, coeff_memory_0_15_port, 
      coeff_memory_0_14_port, coeff_memory_0_13_port, coeff_memory_0_12_port, 
      coeff_memory_0_11_port, coeff_memory_0_10_port, coeff_memory_0_9_port, 
      coeff_memory_0_8_port, coeff_memory_0_7_port, coeff_memory_0_6_port, 
      coeff_memory_0_5_port, coeff_memory_0_4_port, coeff_memory_0_3_port, 
      coeff_memory_0_2_port, coeff_memory_0_1_port, coeff_memory_0_0_port, 
      coeff_memory_1_31_port, coeff_memory_1_30_port, coeff_memory_1_29_port, 
      coeff_memory_1_28_port, coeff_memory_1_27_port, coeff_memory_1_26_port, 
      coeff_memory_1_25_port, coeff_memory_1_24_port, coeff_memory_1_23_port, 
      coeff_memory_1_22_port, coeff_memory_1_21_port, coeff_memory_1_20_port, 
      coeff_memory_1_19_port, coeff_memory_1_18_port, coeff_memory_1_17_port, 
      coeff_memory_1_16_port, coeff_memory_1_15_port, coeff_memory_1_14_port, 
      coeff_memory_1_13_port, coeff_memory_1_12_port, coeff_memory_1_11_port, 
      coeff_memory_1_10_port, coeff_memory_1_9_port, coeff_memory_1_8_port, 
      coeff_memory_1_7_port, coeff_memory_1_6_port, coeff_memory_1_5_port, 
      coeff_memory_1_4_port, coeff_memory_1_3_port, coeff_memory_1_2_port, 
      coeff_memory_1_1_port, coeff_memory_1_0_port, coeff_memory_2_31_port, 
      coeff_memory_2_30_port, coeff_memory_2_29_port, coeff_memory_2_28_port, 
      coeff_memory_2_27_port, coeff_memory_2_26_port, coeff_memory_2_25_port, 
      coeff_memory_2_24_port, coeff_memory_2_23_port, coeff_memory_2_22_port, 
      coeff_memory_2_21_port, coeff_memory_2_20_port, coeff_memory_2_19_port, 
      coeff_memory_2_18_port, coeff_memory_2_17_port, coeff_memory_2_16_port, 
      coeff_memory_2_15_port, coeff_memory_2_14_port, coeff_memory_2_13_port, 
      coeff_memory_2_12_port, coeff_memory_2_11_port, coeff_memory_2_10_port, 
      coeff_memory_2_9_port, coeff_memory_2_8_port, coeff_memory_2_7_port, 
      coeff_memory_2_6_port, coeff_memory_2_5_port, coeff_memory_2_4_port, 
      coeff_memory_2_3_port, coeff_memory_2_2_port, coeff_memory_2_1_port, 
      coeff_memory_2_0_port, coeff_memory_3_31_port, coeff_memory_3_30_port, 
      coeff_memory_3_29_port, coeff_memory_3_28_port, coeff_memory_3_27_port, 
      coeff_memory_3_26_port, coeff_memory_3_25_port, coeff_memory_3_24_port, 
      coeff_memory_3_23_port, coeff_memory_3_22_port, coeff_memory_3_21_port, 
      coeff_memory_3_20_port, coeff_memory_3_19_port, coeff_memory_3_18_port, 
      coeff_memory_3_17_port, coeff_memory_3_16_port, coeff_memory_3_15_port, 
      coeff_memory_3_14_port, coeff_memory_3_13_port, coeff_memory_3_12_port, 
      coeff_memory_3_11_port, coeff_memory_3_10_port, coeff_memory_3_9_port, 
      coeff_memory_3_8_port, coeff_memory_3_7_port, coeff_memory_3_6_port, 
      coeff_memory_3_5_port, coeff_memory_3_4_port, coeff_memory_3_3_port, 
      coeff_memory_3_2_port, coeff_memory_3_1_port, coeff_memory_3_0_port, 
      coeff_memory_4_31_port, coeff_memory_4_30_port, coeff_memory_4_29_port, 
      coeff_memory_4_28_port, coeff_memory_4_27_port, coeff_memory_4_26_port, 
      coeff_memory_4_25_port, coeff_memory_4_24_port, coeff_memory_4_23_port, 
      coeff_memory_4_22_port, coeff_memory_4_21_port, coeff_memory_4_20_port, 
      coeff_memory_4_19_port, coeff_memory_4_18_port, coeff_memory_4_17_port, 
      coeff_memory_4_16_port, coeff_memory_4_15_port, coeff_memory_4_14_port, 
      coeff_memory_4_13_port, coeff_memory_4_12_port, coeff_memory_4_11_port, 
      coeff_memory_4_10_port, coeff_memory_4_9_port, coeff_memory_4_8_port, 
      coeff_memory_4_7_port, coeff_memory_4_6_port, coeff_memory_4_5_port, 
      coeff_memory_4_4_port, coeff_memory_4_3_port, coeff_memory_4_2_port, 
      coeff_memory_4_1_port, coeff_memory_4_0_port, operand_regs_255_port, 
      operand_regs_254_port, operand_regs_253_port, operand_regs_252_port, 
      operand_regs_251_port, operand_regs_250_port, operand_regs_249_port, 
      operand_regs_248_port, operand_regs_247_port, operand_regs_246_port, 
      operand_regs_245_port, operand_regs_244_port, operand_regs_243_port, 
      operand_regs_242_port, operand_regs_241_port, operand_regs_240_port, 
      operand_regs_239_port, operand_regs_238_port, operand_regs_237_port, 
      operand_regs_236_port, operand_regs_235_port, operand_regs_234_port, 
      operand_regs_233_port, operand_regs_232_port, operand_regs_231_port, 
      operand_regs_230_port, operand_regs_229_port, operand_regs_228_port, 
      operand_regs_227_port, operand_regs_226_port, operand_regs_225_port, 
      operand_regs_224_port, operand_regs_223_port, operand_regs_222_port, 
      operand_regs_221_port, operand_regs_220_port, operand_regs_219_port, 
      operand_regs_218_port, operand_regs_217_port, operand_regs_216_port, 
      operand_regs_215_port, operand_regs_214_port, operand_regs_213_port, 
      operand_regs_212_port, operand_regs_211_port, operand_regs_210_port, 
      operand_regs_209_port, operand_regs_208_port, operand_regs_207_port, 
      operand_regs_206_port, operand_regs_205_port, operand_regs_204_port, 
      operand_regs_203_port, operand_regs_202_port, operand_regs_201_port, 
      operand_regs_200_port, operand_regs_199_port, operand_regs_198_port, 
      operand_regs_197_port, operand_regs_196_port, operand_regs_195_port, 
      operand_regs_194_port, operand_regs_193_port, operand_regs_192_port, 
      operand_regs_191_port, operand_regs_190_port, operand_regs_189_port, 
      operand_regs_188_port, operand_regs_187_port, operand_regs_186_port, 
      operand_regs_185_port, operand_regs_184_port, operand_regs_183_port, 
      operand_regs_182_port, operand_regs_181_port, operand_regs_180_port, 
      operand_regs_179_port, operand_regs_178_port, operand_regs_177_port, 
      operand_regs_176_port, operand_regs_175_port, operand_regs_174_port, 
      operand_regs_173_port, operand_regs_172_port, operand_regs_171_port, 
      operand_regs_170_port, operand_regs_169_port, operand_regs_168_port, 
      operand_regs_167_port, operand_regs_166_port, operand_regs_165_port, 
      operand_regs_164_port, operand_regs_163_port, operand_regs_162_port, 
      operand_regs_161_port, operand_regs_160_port, operand_regs_159_port, 
      operand_regs_158_port, operand_regs_157_port, operand_regs_156_port, 
      operand_regs_155_port, operand_regs_154_port, operand_regs_153_port, 
      operand_regs_152_port, operand_regs_151_port, operand_regs_150_port, 
      operand_regs_149_port, operand_regs_148_port, operand_regs_147_port, 
      operand_regs_146_port, operand_regs_145_port, operand_regs_144_port, 
      operand_regs_143_port, operand_regs_142_port, operand_regs_141_port, 
      operand_regs_140_port, operand_regs_139_port, operand_regs_138_port, 
      operand_regs_137_port, operand_regs_136_port, operand_regs_135_port, 
      operand_regs_134_port, operand_regs_133_port, operand_regs_132_port, 
      operand_regs_131_port, operand_regs_130_port, operand_regs_129_port, 
      operand_regs_128_port, operand_regs_127_port, operand_regs_126_port, 
      operand_regs_125_port, operand_regs_124_port, operand_regs_123_port, 
      operand_regs_122_port, operand_regs_121_port, operand_regs_120_port, 
      operand_regs_119_port, operand_regs_118_port, operand_regs_117_port, 
      operand_regs_116_port, operand_regs_115_port, operand_regs_114_port, 
      operand_regs_113_port, operand_regs_112_port, operand_regs_111_port, 
      operand_regs_110_port, operand_regs_109_port, operand_regs_108_port, 
      operand_regs_107_port, operand_regs_106_port, operand_regs_105_port, 
      operand_regs_104_port, operand_regs_103_port, operand_regs_102_port, 
      operand_regs_101_port, operand_regs_100_port, operand_regs_99_port, 
      operand_regs_98_port, operand_regs_97_port, operand_regs_96_port, 
      operand_regs_95_port, operand_regs_94_port, operand_regs_93_port, 
      operand_regs_92_port, operand_regs_91_port, operand_regs_90_port, 
      operand_regs_89_port, operand_regs_88_port, operand_regs_87_port, 
      operand_regs_86_port, operand_regs_85_port, operand_regs_84_port, 
      operand_regs_83_port, operand_regs_82_port, operand_regs_81_port, 
      operand_regs_80_port, operand_regs_79_port, operand_regs_78_port, 
      operand_regs_77_port, operand_regs_76_port, operand_regs_75_port, 
      operand_regs_74_port, operand_regs_73_port, operand_regs_72_port, 
      operand_regs_71_port, operand_regs_70_port, operand_regs_69_port, 
      operand_regs_68_port, operand_regs_67_port, operand_regs_66_port, 
      operand_regs_65_port, operand_regs_64_port, operand_regs_63_port, 
      operand_regs_62_port, operand_regs_61_port, operand_regs_60_port, 
      operand_regs_59_port, operand_regs_58_port, operand_regs_57_port, 
      operand_regs_56_port, operand_regs_55_port, operand_regs_54_port, 
      operand_regs_53_port, operand_regs_52_port, operand_regs_51_port, 
      operand_regs_50_port, operand_regs_49_port, operand_regs_48_port, 
      operand_regs_47_port, operand_regs_46_port, operand_regs_45_port, 
      operand_regs_44_port, operand_regs_43_port, operand_regs_42_port, 
      operand_regs_41_port, operand_regs_40_port, operand_regs_39_port, 
      operand_regs_38_port, operand_regs_37_port, operand_regs_36_port, 
      operand_regs_35_port, operand_regs_34_port, operand_regs_33_port, 
      operand_regs_32_port, operand_regs_31_port, operand_regs_30_port, 
      operand_regs_29_port, operand_regs_28_port, operand_regs_27_port, 
      operand_regs_26_port, operand_regs_25_port, operand_regs_24_port, 
      operand_regs_23_port, operand_regs_22_port, operand_regs_21_port, 
      operand_regs_20_port, operand_regs_19_port, operand_regs_18_port, 
      operand_regs_17_port, operand_regs_16_port, operand_regs_15_port, 
      operand_regs_14_port, operand_regs_13_port, operand_regs_12_port, 
      operand_regs_11_port, operand_regs_10_port, operand_regs_9_port, 
      operand_regs_8_port, operand_regs_7_port, operand_regs_6_port, 
      operand_regs_5_port, operand_regs_4_port, operand_regs_3_port, 
      operand_regs_2_port, operand_regs_1_port, operand_regs_0_port, in_trigger
      , out_trigger, coeff_load, operand_load, read_comp_res, filt_mult_inputs,
      N66, comp_res_159_port, comp_res_158_port, comp_res_157_port, 
      comp_res_156_port, comp_res_155_port, comp_res_154_port, 
      comp_res_153_port, comp_res_152_port, comp_res_151_port, 
      comp_res_150_port, comp_res_149_port, comp_res_148_port, 
      comp_res_147_port, comp_res_146_port, comp_res_145_port, 
      comp_res_144_port, comp_res_143_port, comp_res_142_port, 
      comp_res_141_port, comp_res_140_port, comp_res_139_port, 
      comp_res_138_port, comp_res_137_port, comp_res_136_port, 
      comp_res_135_port, comp_res_134_port, comp_res_133_port, 
      comp_res_132_port, comp_res_131_port, comp_res_130_port, 
      comp_res_129_port, comp_res_128_port, comp_res_127_port, 
      comp_res_126_port, comp_res_125_port, comp_res_124_port, 
      comp_res_123_port, comp_res_122_port, comp_res_121_port, 
      comp_res_120_port, comp_res_119_port, comp_res_118_port, 
      comp_res_117_port, comp_res_116_port, comp_res_115_port, 
      comp_res_114_port, comp_res_113_port, comp_res_112_port, 
      comp_res_111_port, comp_res_110_port, comp_res_109_port, 
      comp_res_108_port, comp_res_107_port, comp_res_106_port, 
      comp_res_105_port, comp_res_104_port, comp_res_103_port, 
      comp_res_102_port, comp_res_101_port, comp_res_100_port, comp_res_99_port
      , comp_res_98_port, comp_res_97_port, comp_res_96_port, comp_res_95_port,
      comp_res_94_port, comp_res_93_port, comp_res_92_port, comp_res_91_port, 
      comp_res_90_port, comp_res_89_port, comp_res_88_port, comp_res_87_port, 
      comp_res_86_port, comp_res_85_port, comp_res_84_port, comp_res_83_port, 
      comp_res_82_port, comp_res_81_port, comp_res_80_port, comp_res_79_port, 
      comp_res_78_port, comp_res_77_port, comp_res_76_port, comp_res_75_port, 
      comp_res_74_port, comp_res_73_port, comp_res_72_port, comp_res_71_port, 
      comp_res_70_port, comp_res_69_port, comp_res_68_port, comp_res_67_port, 
      comp_res_66_port, comp_res_65_port, comp_res_64_port, comp_res_63_port, 
      comp_res_62_port, comp_res_61_port, comp_res_60_port, comp_res_59_port, 
      comp_res_58_port, comp_res_57_port, comp_res_56_port, comp_res_55_port, 
      comp_res_54_port, comp_res_53_port, comp_res_52_port, comp_res_51_port, 
      comp_res_50_port, comp_res_49_port, comp_res_48_port, comp_res_47_port, 
      comp_res_46_port, comp_res_45_port, comp_res_44_port, comp_res_43_port, 
      comp_res_42_port, comp_res_41_port, comp_res_40_port, comp_res_39_port, 
      comp_res_38_port, comp_res_37_port, comp_res_36_port, comp_res_35_port, 
      comp_res_34_port, comp_res_33_port, comp_res_32_port, comp_res_31_port, 
      comp_res_30_port, comp_res_29_port, comp_res_28_port, comp_res_27_port, 
      comp_res_26_port, comp_res_25_port, comp_res_24_port, comp_res_23_port, 
      comp_res_22_port, comp_res_21_port, comp_res_20_port, comp_res_19_port, 
      comp_res_18_port, comp_res_17_port, comp_res_16_port, comp_res_15_port, 
      comp_res_14_port, comp_res_13_port, comp_res_12_port, comp_res_11_port, 
      comp_res_10_port, comp_res_9_port, comp_res_8_port, comp_res_7_port, 
      comp_res_6_port, comp_res_5_port, comp_res_4_port, comp_res_3_port, 
      comp_res_2_port, comp_res_1_port, comp_res_0_port, N1978, N1979, N1980, 
      N1981, N1982, N1983, N1984, N1985, N1986, N1987, N1988, N1989, N1990, 
      N1991, N1992, N1993, N1994, N1995, N1996, N1997, N1998, N1999, N2000, 
      N2001, N2002, N2003, N2004, N2005, N2006, N2007, N2008, N2009, 
      in_buf_255_port, in_buf_254_port, in_buf_253_port, in_buf_252_port, 
      in_buf_251_port, in_buf_250_port, in_buf_249_port, in_buf_248_port, 
      in_buf_247_port, in_buf_246_port, in_buf_245_port, in_buf_244_port, 
      in_buf_243_port, in_buf_242_port, in_buf_241_port, in_buf_240_port, 
      in_buf_239_port, in_buf_238_port, in_buf_237_port, in_buf_236_port, 
      in_buf_235_port, in_buf_234_port, in_buf_233_port, in_buf_232_port, 
      in_buf_231_port, in_buf_230_port, in_buf_229_port, in_buf_228_port, 
      in_buf_227_port, in_buf_226_port, in_buf_225_port, in_buf_224_port, 
      in_buf_223_port, in_buf_222_port, in_buf_221_port, in_buf_220_port, 
      in_buf_219_port, in_buf_218_port, in_buf_217_port, in_buf_216_port, 
      in_buf_215_port, in_buf_214_port, in_buf_213_port, in_buf_212_port, 
      in_buf_211_port, in_buf_210_port, in_buf_209_port, in_buf_208_port, 
      in_buf_207_port, in_buf_206_port, in_buf_205_port, in_buf_204_port, 
      in_buf_203_port, in_buf_202_port, in_buf_201_port, in_buf_200_port, 
      in_buf_199_port, in_buf_198_port, in_buf_197_port, in_buf_196_port, 
      in_buf_195_port, in_buf_194_port, in_buf_193_port, in_buf_192_port, 
      in_buf_191_port, in_buf_190_port, in_buf_189_port, in_buf_188_port, 
      in_buf_187_port, in_buf_186_port, in_buf_185_port, in_buf_184_port, 
      in_buf_183_port, in_buf_182_port, in_buf_181_port, in_buf_180_port, 
      in_buf_179_port, in_buf_178_port, in_buf_177_port, in_buf_176_port, 
      in_buf_175_port, in_buf_174_port, in_buf_173_port, in_buf_172_port, 
      in_buf_171_port, in_buf_170_port, in_buf_169_port, in_buf_168_port, 
      in_buf_167_port, in_buf_166_port, in_buf_165_port, in_buf_164_port, 
      in_buf_163_port, in_buf_162_port, in_buf_161_port, in_buf_160_port, 
      in_buf_159_port, in_buf_158_port, in_buf_157_port, in_buf_156_port, 
      in_buf_155_port, in_buf_154_port, in_buf_153_port, in_buf_152_port, 
      in_buf_151_port, in_buf_150_port, in_buf_149_port, in_buf_148_port, 
      in_buf_147_port, in_buf_146_port, in_buf_145_port, in_buf_144_port, 
      in_buf_143_port, in_buf_142_port, in_buf_141_port, in_buf_140_port, 
      in_buf_139_port, in_buf_138_port, in_buf_137_port, in_buf_136_port, 
      in_buf_135_port, in_buf_134_port, in_buf_133_port, in_buf_132_port, 
      in_buf_131_port, in_buf_130_port, in_buf_129_port, in_buf_128_port, 
      in_buf_127_port, in_buf_126_port, in_buf_125_port, in_buf_124_port, 
      in_buf_123_port, in_buf_122_port, in_buf_121_port, in_buf_120_port, 
      in_buf_119_port, in_buf_118_port, in_buf_117_port, in_buf_116_port, 
      in_buf_115_port, in_buf_114_port, in_buf_113_port, in_buf_112_port, 
      in_buf_111_port, in_buf_110_port, in_buf_109_port, in_buf_108_port, 
      in_buf_107_port, in_buf_106_port, in_buf_105_port, in_buf_104_port, 
      in_buf_103_port, in_buf_102_port, in_buf_101_port, in_buf_100_port, 
      in_buf_99_port, in_buf_98_port, in_buf_97_port, in_buf_96_port, 
      in_buf_95_port, in_buf_94_port, in_buf_93_port, in_buf_92_port, 
      in_buf_91_port, in_buf_90_port, in_buf_89_port, in_buf_88_port, 
      in_buf_87_port, in_buf_86_port, in_buf_85_port, in_buf_84_port, 
      in_buf_83_port, in_buf_82_port, in_buf_81_port, in_buf_80_port, 
      in_buf_79_port, in_buf_78_port, in_buf_77_port, in_buf_76_port, 
      in_buf_75_port, in_buf_74_port, in_buf_73_port, in_buf_72_port, 
      in_buf_71_port, in_buf_70_port, in_buf_69_port, in_buf_68_port, 
      in_buf_67_port, in_buf_66_port, in_buf_65_port, in_buf_64_port, 
      in_buf_63_port, in_buf_62_port, in_buf_61_port, in_buf_60_port, 
      in_buf_59_port, in_buf_58_port, in_buf_57_port, in_buf_56_port, 
      in_buf_55_port, in_buf_54_port, in_buf_53_port, in_buf_52_port, 
      in_buf_51_port, in_buf_50_port, in_buf_49_port, in_buf_48_port, 
      in_buf_47_port, in_buf_46_port, in_buf_45_port, in_buf_44_port, 
      in_buf_43_port, in_buf_42_port, in_buf_41_port, in_buf_40_port, 
      in_buf_39_port, in_buf_38_port, in_buf_37_port, in_buf_36_port, 
      in_buf_35_port, in_buf_34_port, in_buf_33_port, in_buf_32_port, 
      in_buf_31_port, in_buf_30_port, in_buf_29_port, in_buf_28_port, 
      in_buf_27_port, in_buf_26_port, in_buf_25_port, in_buf_24_port, 
      in_buf_23_port, in_buf_22_port, in_buf_21_port, in_buf_20_port, 
      in_buf_19_port, in_buf_18_port, in_buf_17_port, in_buf_16_port, 
      in_buf_15_port, in_buf_14_port, in_buf_13_port, in_buf_12_port, 
      in_buf_11_port, in_buf_10_port, in_buf_9_port, in_buf_8_port, 
      in_buf_7_port, in_buf_6_port, in_buf_5_port, in_buf_4_port, in_buf_3_port
      , in_buf_2_port, in_buf_1_port, in_buf_0_port, N2010, N2011, N2012, N2013
      , N2014, N2015, N2016, N2017, N2018, N2019, N2020, N2021, N2022, N2023, 
      N2024, N2025, N2026, N2027, N2028, N2029, N2030, N2031, N2032, N2033, 
      N2034, N2035, N2036, N2037, N2038, N2039, N2040, N2041, in_busy, out_busy
      , in_counter_2_port, in_counter_1_port, in_counter_0_port, odd, odd1, 
      N2850, N2851, N2852, N2853, N2854, N2855, N2856, N2857, N2858, N2859, 
      N2860, N2861, N2862, N2863, N2864, N2865, N2867, N2868, N2869, N2870, 
      N2871, N2872, N2873, N2874, N2875, N2876, N2877, N2878, N2879, N2880, 
      N2881, N2882, N2888, N2889, N2890, N2891, N2892, N2893, N2894, N2895, 
      N2896, N2897, N2898, N2899, N2900, N2901, N2902, N2903, N2913, N2914, 
      N2915, N2916, N2917, N2918, N2919, N2920, N2921, N2922, N2923, N2924, 
      N2925, N2926, N2927, N2928, N2929, N2930, N2931, N2932, N2933, N2934, 
      N2935, N2936, N2937, N2938, N2939, N2940, N2941, N2942, N2943, N2944, 
      N2945, N2946, N2947, N2948, N2949, N2950, N2951, N2952, N2953, N2954, 
      N2955, N2956, N2957, N2958, N2959, N2960, N2961, N2962, N2963, N2964, 
      N2965, N2966, N2967, N2968, N2969, N2970, N2971, N2972, N2973, N2974, 
      N2975, N2976, N2977, N2978, N2979, N2980, N2981, N2982, N2983, N2984, 
      N2985, N2986, N2987, N2988, N2989, N2990, N2991, N2992, N2993, N2994, 
      N2995, N2996, N2997, N2998, N2999, N3000, N3001, N3002, N3003, N3004, 
      N3005, N3006, N3007, N3008, N3009, N3010, N3011, N3012, N3013, N3014, 
      N3015, N3016, N3017, N3018, N3019, N3020, N3021, N3022, N3023, N3024, 
      N3025, N3026, N3027, N3028, N3029, N3030, N3031, N3032, N3033, N3034, 
      N3035, N3036, N3037, N3038, N3039, N3040, N3041, N3042, N3043, N3044, 
      N3045, N3046, N3047, N3048, N3049, N3050, N3051, N3052, N3053, N3054, 
      N3055, N3056, N3057, N3058, N3059, N3060, N3061, N3062, N3063, N3064, 
      N3065, N3066, N3067, N3068, N3069, N3070, N3071, N3072, N3073, N3074, 
      N3075, N3076, N3077, N3078, N3079, N3080, N3081, N3082, N3083, N3084, 
      N3085, N3086, N3087, N3088, N3089, N3090, N3091, N3092, N3093, N3094, 
      N3095, N3096, N3097, N3098, N3099, N3100, N3101, N3102, N3103, N3104, 
      N3105, N3106, N3107, N3108, N3109, N3110, N3111, N3112, N3113, N3114, 
      N3115, N3116, N3117, N3118, N3119, N3120, N3121, N3122, N3123, N3124, 
      N3125, N3126, N3127, N3128, N3129, N3130, N3131, N3132, N3133, N3134, 
      N3135, N3136, N3137, N3138, N3139, N3140, N3141, N3142, N3143, N3144, 
      N3145, N3146, N3147, N3148, N3149, N3150, N3151, N3152, N3153, N3154, 
      N3155, N3156, N3157, N3158, N3159, N3160, N3161, N3162, N3163, N3164, 
      N3165, N3166, N3167, N3168, N3201, N3202, N3203, N3204, N3205, N3206, 
      N3207, N3208, N3209, N3210, N3211, N3212, N3213, N3214, N3215, N3216, 
      N3217, N3218, N3219, N3220, N3221, N3222, N3223, N3224, N3225, N3226, 
      N3227, N3228, N3229, N3230, N3231, N3232, N3233, N3234, N3235, N3236, 
      N3237, N3238, N3239, N3240, N3241, N3242, N3243, N3244, N3245, N3246, 
      N3247, N3248, N3249, N3250, N3251, N3252, N3253, N3254, N3255, N3256, 
      N3257, N3258, N3259, N3260, N3261, N3262, N3263, N3264, N3265, N3266, 
      N3267, N3268, N3269, N3270, N3271, N3272, N3273, N3274, N3275, N3276, 
      N3277, N3278, N3279, N3280, N3281, N3282, N3283, N3284, N3285, N3286, 
      N3287, N3288, N3289, N3290, N3291, N3292, N3293, N3294, N3295, N3296, 
      N3297, N3298, N3299, N3300, N3301, N3302, N3303, N3304, N3305, N3306, 
      N3307, N3308, N3309, N3310, N3311, N3312, N3313, N3314, N3315, N3316, 
      N3317, N3318, N3319, N3320, N3321, N3322, N3323, N3324, N3325, N3326, 
      N3327, N3328, N3329, N3330, N3331, N3332, N3333, N3334, N3335, N3336, 
      N3337, N3338, N3339, N3340, N3341, N3342, N3343, N3344, N3345, N3346, 
      N3347, N3348, N3349, N3350, N3351, N3352, N3353, N3354, N3355, N3356, 
      N3357, N3358, N3359, N3360, N3361, N3362, N3363, N3364, N3365, N3366, 
      N3367, N3368, N3369, N3370, N3371, N3372, N3373, N3374, N3375, N3376, 
      N3377, N3378, N3379, N3380, N3381, N3382, N3383, N3384, N3385, N3386, 
      N3387, N3388, N3389, N3390, N3391, N3392, n4, n5, n10, n12, n13, n14, n15
      , n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44
      , n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, 
      n5900, n6000, n6100, n6300, n6400, n65, n68, n69, n70, n72, n73, n74, n76
      , n77, n78, n79, n81, n84, n85, n86, n87, n88, n89, n91, n92, n93, n95, 
      n96, n97, n99, n100, n101, n103, n104, n106, n107, n108, n109, n110, n111
      , n114, n115, n118, n119, n120, n122, n123, n124, n125, n126, n127, n128,
      n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, 
      n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, 
      n153, n154, n155, n156, n157, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, 
      n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, 
      n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, 
      n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, 
      n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, 
      n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, 
      n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, 
      n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, 
      n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, 
      n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, 
      n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, 
      n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, 
      n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, 
      n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, 
      n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, 
      n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, 
      n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, 
      n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, 
      n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, 
      n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, 
      n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, 
      n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, 
      n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, 
      n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, 
      n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, 
      n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, 
      n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, 
      n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, 
      n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, 
      n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, 
      n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, 
      n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, 
      n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, 
      n585, n586, n587, n588, n589, n5901, n591, n592, n593, n594, n595, n596, 
      n597, n598, n599, n6001, n601, n602, n603, n604, n605, n606, n607, n608, 
      n609, n6101, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, 
      n621, n622, n623, n624, n625, n626, n627, n628, n629, n6301, n631, n632, 
      n633, n634, n635, n636, n637, n638, n639, n6401, n641, n642, n643, n644, 
      n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, 
      n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, 
      n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, 
      n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, 
      n693, n694, n695, n696, n697, n_1160, n_1161, n_1162, n_1163, n_1164, 
      n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, 
      n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, 
      n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, 
      n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, 
      n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, 
      n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, 
      n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, 
      n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, 
      n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, 
      n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, 
      n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, 
      n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, 
      n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, 
      n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, 
      n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, 
      n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, 
      n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, 
      n_1318, n_1319 : std_logic;

begin
   avs_readdata <= ( avs_readdata_31_port, avs_readdata_30_port, 
      avs_readdata_29_port, avs_readdata_28_port, avs_readdata_27_port, 
      avs_readdata_26_port, avs_readdata_25_port, avs_readdata_24_port, 
      avs_readdata_23_port, avs_readdata_22_port, avs_readdata_21_port, 
      avs_readdata_20_port, avs_readdata_19_port, avs_readdata_18_port, 
      avs_readdata_17_port, avs_readdata_16_port, avs_readdata_15_port, 
      avs_readdata_14_port, avs_readdata_13_port, avs_readdata_12_port, 
      avs_readdata_11_port, avs_readdata_10_port, avs_readdata_9_port, 
      avs_readdata_8_port, avs_readdata_7_port, avs_readdata_6_port, 
      avs_readdata_5_port, avs_readdata_4_port, avs_readdata_3_port, 
      avs_readdata_2_port, avs_readdata_1_port, avs_readdata_0_port );
   clk_out <= clk;
   stop_sim <= stop_sim_port;
   
   U3 : OAI22D1 port map( A1 => N63, A2 => n4, B1 => n5, B2 => n697, Z => n201)
                           ;
   U4 : AOI21D1 port map( A1 => out_busy, A2 => n694, B => n684, Z => n5);
   U7 : AOI22D1 port map( A1 => N1978, A2 => n267, B1 => N2010, B2 => n674, Z 
                           => n10);
   U9 : AOI22D1 port map( A1 => N2011, A2 => n12, B1 => avs_readdata_30_port, 
                           B2 => n676, Z => n15);
   U12 : AOI22D1 port map( A1 => N1980, A2 => n267, B1 => N2012, B2 => n674, Z 
                           => n16);
   U14 : AOI22D1 port map( A1 => N2013, A2 => n674, B1 => avs_readdata_28_port,
                           B2 => n676, Z => n18);
   U17 : AOI22D1 port map( A1 => N1982, A2 => n267, B1 => N2014, B2 => n674, Z 
                           => n19);
   U19 : AOI22D1 port map( A1 => N2015, A2 => n674, B1 => avs_readdata_26_port,
                           B2 => n676, Z => n21);
   U22 : AOI22D1 port map( A1 => N1984, A2 => n267, B1 => N2016, B2 => n674, Z 
                           => n22);
   U24 : AOI22D1 port map( A1 => N2017, A2 => n674, B1 => avs_readdata_24_port,
                           B2 => n676, Z => n24);
   U27 : AOI22D1 port map( A1 => N1986, A2 => n267, B1 => N2018, B2 => n674, Z 
                           => n25);
   U29 : AOI22D1 port map( A1 => N2019, A2 => n12, B1 => avs_readdata_22_port, 
                           B2 => n676, Z => n27);
   U32 : AOI22D1 port map( A1 => N1988, A2 => n267, B1 => N2020, B2 => n674, Z 
                           => n28);
   U34 : AOI22D1 port map( A1 => N2021, A2 => n12, B1 => avs_readdata_20_port, 
                           B2 => n676, Z => n30);
   U37 : AOI22D1 port map( A1 => N1990, A2 => n267, B1 => N2022, B2 => n674, Z 
                           => n31);
   U39 : AOI22D1 port map( A1 => N2023, A2 => n12, B1 => avs_readdata_18_port, 
                           B2 => n676, Z => n33);
   U42 : AOI22D1 port map( A1 => N1992, A2 => n267, B1 => N2024, B2 => n674, Z 
                           => n34);
   U44 : AOI22D1 port map( A1 => N2025, A2 => n12, B1 => avs_readdata_16_port, 
                           B2 => n676, Z => n36);
   U47 : AOI22D1 port map( A1 => N1994, A2 => n267, B1 => N2026, B2 => n674, Z 
                           => n37);
   U49 : AOI22D1 port map( A1 => N2027, A2 => n12, B1 => avs_readdata_14_port, 
                           B2 => n676, Z => n39);
   U52 : AOI22D1 port map( A1 => N1996, A2 => n267, B1 => N2028, B2 => n12, Z 
                           => n40);
   U54 : AOI22D1 port map( A1 => N2029, A2 => n12, B1 => avs_readdata_12_port, 
                           B2 => n676, Z => n42);
   U57 : AOI22D1 port map( A1 => N1998, A2 => n267, B1 => N2030, B2 => n12, Z 
                           => n43);
   U59 : AOI22D1 port map( A1 => N2031, A2 => n12, B1 => avs_readdata_10_port, 
                           B2 => n676, Z => n45);
   U62 : AOI22D1 port map( A1 => N2000, A2 => n267, B1 => N2032, B2 => n12, Z 
                           => n46);
   U64 : AOI22D1 port map( A1 => N2033, A2 => n12, B1 => avs_readdata_8_port, 
                           B2 => n676, Z => n48);
   U67 : AOI22D1 port map( A1 => N2002, A2 => n267, B1 => N2034, B2 => n674, Z 
                           => n49);
   U69 : AOI22D1 port map( A1 => N2035, A2 => n12, B1 => avs_readdata_6_port, 
                           B2 => n676, Z => n51);
   U72 : AOI22D1 port map( A1 => N2004, A2 => n267, B1 => N2036, B2 => n674, Z 
                           => n52);
   U74 : AOI22D1 port map( A1 => N2037, A2 => n12, B1 => avs_readdata_4_port, 
                           B2 => n676, Z => n54);
   U77 : AOI22D1 port map( A1 => N2006, A2 => n267, B1 => N2038, B2 => n674, Z 
                           => n55);
   U79 : AOI22D1 port map( A1 => N2039, A2 => n12, B1 => avs_readdata_2_port, 
                           B2 => n676, Z => n57);
   U82 : AOI22D1 port map( A1 => N2008, A2 => n267, B1 => N2040, B2 => n674, Z 
                           => n58);
   U84 : AOI22D1 port map( A1 => N2041, A2 => n674, B1 => avs_readdata_0_port, 
                           B2 => n676, Z => n6100);
   U94 : AOI21D1 port map( A1 => n678, A2 => in_trigger, B => n72, Z => n70);
   U95 : OAI22D1 port map( A1 => n6400, A2 => n73, B1 => n74, B2 => n685, Z => 
                           n72);
   U96 : AOI22D1 port map( A1 => in_busy, A2 => n69, B1 => out_busy, B2 => n68,
                           Z => n73);
   U97 : EXNOR2D1 port map( A1 => n695, A2 => n76, Z => n234);
   U98 : AOI22D1 port map( A1 => n77, A2 => out_busy, B1 => n695, B2 => n685, Z
                           => n76);
   U100 : OAI22D1 port map( A1 => n697, A2 => n4, B1 => n79, B2 => n671, Z => 
                           n235);
   U103 : OAI32D1 port map( A1 => n684, A2 => N62, A3 => n695, B1 => n694, B2 
                           => n81, Z => n236);
   U105 : OAI32D1 port map( A1 => n696, A2 => n695, A3 => n78, B1 => out_busy, 
                           B2 => n685, Z => n81);
   U111 : OAI211D1 port map( A1 => n692, A2 => n84, B => n85, C => n86, Z => 
                           n237);
   U113 : OAI22D1 port map( A1 => n683, A2 => n88, B1 => n89, B2 => n693, Z => 
                           n238);
   U115 : EXNOR2D1 port map( A1 => in_busy, A2 => n161, Z => n239);
   U117 : AOI22D1 port map( A1 => avs_writedata(0), A2 => n677, B1 => 
                           out_trigger, B2 => n74, Z => n92);
   U122 : AOI22D1 port map( A1 => avs_writedata(0), A2 => n678, B1 => 
                           in_trigger, B2 => n96, Z => n95);
   U125 : EXNOR2D1 port map( A1 => n695, A2 => n672, Z => n154);
   U126 : EXNOR2D1 port map( A1 => n687, A2 => in_busy, Z => n156);
   U130 : AOI22D1 port map( A1 => odd, A2 => n91, B1 => n101, B2 => in_busy, Z 
                           => n100);
   U131 : OAI21D1 port map( A1 => in_counter_1_port, A2 => n690, B => n688, Z 
                           => n91);
   U200 : OA21M20D1 port map( A1 => n690, A2 => in_trigger, B => n176, Z => 
                           n161);
   mult_21_C241 : gp_custom_DW_mult_tc_2 port map( a(31) => N2944, a(30) => 
                           N2943, a(29) => N2942, a(28) => N2941, a(27) => 
                           N2940, a(26) => N2939, a(25) => N2938, a(24) => 
                           N2937, a(23) => N2936, a(22) => N2935, a(21) => 
                           N2934, a(20) => N2933, a(19) => N2932, a(18) => 
                           N2931, a(17) => N2930, a(16) => N2929, a(15) => 
                           N2928, a(14) => N2927, a(13) => N2926, a(12) => 
                           N2925, a(11) => N2924, a(10) => N2923, a(9) => N2922
                           , a(8) => N2921, a(7) => N2920, a(6) => N2919, a(5) 
                           => N2918, a(4) => N2917, a(3) => N2916, a(2) => 
                           N2915, a(1) => N2914, a(0) => N2913, b(31) => N3104,
                           b(30) => N3103, b(29) => N3102, b(28) => N3101, 
                           b(27) => N3100, b(26) => N3099, b(25) => N3098, 
                           b(24) => N3097, b(23) => N3096, b(22) => N3095, 
                           b(21) => N3094, b(20) => N3093, b(19) => N3092, 
                           b(18) => N3091, b(17) => N3090, b(16) => N3089, 
                           b(15) => N3088, b(14) => N3087, b(13) => N3086, 
                           b(12) => N3085, b(11) => N3084, b(10) => N3083, b(9)
                           => N3082, b(8) => N3081, b(7) => N3080, b(6) => 
                           N3079, b(5) => N3078, b(4) => N3077, b(3) => N3076, 
                           b(2) => N3075, b(1) => N3074, b(0) => N3073, 
                           product(63) => n_1160, product(62) => n_1161, 
                           product(61) => n_1162, product(60) => n_1163, 
                           product(59) => n_1164, product(58) => n_1165, 
                           product(57) => n_1166, product(56) => n_1167, 
                           product(55) => n_1168, product(54) => n_1169, 
                           product(53) => n_1170, product(52) => n_1171, 
                           product(51) => n_1172, product(50) => n_1173, 
                           product(49) => n_1174, product(48) => n_1175, 
                           product(47) => n_1176, product(46) => n_1177, 
                           product(45) => n_1178, product(44) => n_1179, 
                           product(43) => n_1180, product(42) => n_1181, 
                           product(41) => n_1182, product(40) => n_1183, 
                           product(39) => n_1184, product(38) => n_1185, 
                           product(37) => n_1186, product(36) => n_1187, 
                           product(35) => n_1188, product(34) => n_1189, 
                           product(33) => n_1190, product(32) => n_1191, 
                           product(31) => N3264, product(30) => N3263, 
                           product(29) => N3262, product(28) => N3261, 
                           product(27) => N3260, product(26) => N3259, 
                           product(25) => N3258, product(24) => N3257, 
                           product(23) => N3256, product(22) => N3255, 
                           product(21) => N3254, product(20) => N3253, 
                           product(19) => N3252, product(18) => N3251, 
                           product(17) => N3250, product(16) => N3249, 
                           product(15) => N3248, product(14) => N3247, 
                           product(13) => N3246, product(12) => N3245, 
                           product(11) => N3244, product(10) => N3243, 
                           product(9) => N3242, product(8) => N3241, product(7)
                           => N3240, product(6) => N3239, product(5) => N3238, 
                           product(4) => N3237, product(3) => N3236, product(2)
                           => N3235, product(1) => N3234, product(0) => N3233);
   mult_21_C243 : gp_custom_DW_mult_tc_3 port map( a(31) => N2976, a(30) => 
                           N2975, a(29) => N2974, a(28) => N2973, a(27) => 
                           N2972, a(26) => N2971, a(25) => N2970, a(24) => 
                           N2969, a(23) => N2968, a(22) => N2967, a(21) => 
                           N2966, a(20) => N2965, a(19) => N2964, a(18) => 
                           N2963, a(17) => N2962, a(16) => N2961, a(15) => 
                           N2960, a(14) => N2959, a(13) => N2958, a(12) => 
                           N2957, a(11) => N2956, a(10) => N2955, a(9) => N2954
                           , a(8) => N2953, a(7) => N2952, a(6) => N2951, a(5) 
                           => N2950, a(4) => N2949, a(3) => N2948, a(2) => 
                           N2947, a(1) => N2946, a(0) => N2945, b(31) => N3136,
                           b(30) => N3135, b(29) => N3134, b(28) => N3133, 
                           b(27) => N3132, b(26) => N3131, b(25) => N3130, 
                           b(24) => N3129, b(23) => N3128, b(22) => N3127, 
                           b(21) => N3126, b(20) => N3125, b(19) => N3124, 
                           b(18) => N3123, b(17) => N3122, b(16) => N3121, 
                           b(15) => N3120, b(14) => N3119, b(13) => N3118, 
                           b(12) => N3117, b(11) => N3116, b(10) => N3115, b(9)
                           => N3114, b(8) => N3113, b(7) => N3112, b(6) => 
                           N3111, b(5) => N3110, b(4) => N3109, b(3) => N3108, 
                           b(2) => N3107, b(1) => N3106, b(0) => N3105, 
                           product(63) => n_1192, product(62) => n_1193, 
                           product(61) => n_1194, product(60) => n_1195, 
                           product(59) => n_1196, product(58) => n_1197, 
                           product(57) => n_1198, product(56) => n_1199, 
                           product(55) => n_1200, product(54) => n_1201, 
                           product(53) => n_1202, product(52) => n_1203, 
                           product(51) => n_1204, product(50) => n_1205, 
                           product(49) => n_1206, product(48) => n_1207, 
                           product(47) => n_1208, product(46) => n_1209, 
                           product(45) => n_1210, product(44) => n_1211, 
                           product(43) => n_1212, product(42) => n_1213, 
                           product(41) => n_1214, product(40) => n_1215, 
                           product(39) => n_1216, product(38) => n_1217, 
                           product(37) => n_1218, product(36) => n_1219, 
                           product(35) => n_1220, product(34) => n_1221, 
                           product(33) => n_1222, product(32) => n_1223, 
                           product(31) => N3296, product(30) => N3295, 
                           product(29) => N3294, product(28) => N3293, 
                           product(27) => N3292, product(26) => N3291, 
                           product(25) => N3290, product(24) => N3289, 
                           product(23) => N3288, product(22) => N3287, 
                           product(21) => N3286, product(20) => N3285, 
                           product(19) => N3284, product(18) => N3283, 
                           product(17) => N3282, product(16) => N3281, 
                           product(15) => N3280, product(14) => N3279, 
                           product(13) => N3278, product(12) => N3277, 
                           product(11) => N3276, product(10) => N3275, 
                           product(9) => N3274, product(8) => N3273, product(7)
                           => N3272, product(6) => N3271, product(5) => N3270, 
                           product(4) => N3269, product(3) => N3268, product(2)
                           => N3267, product(1) => N3266, product(0) => N3265);
   mult_21_C245 : gp_custom_DW_mult_tc_4 port map( a(31) => N3008, a(30) => 
                           N3007, a(29) => N3006, a(28) => N3005, a(27) => 
                           N3004, a(26) => N3003, a(25) => N3002, a(24) => 
                           N3001, a(23) => N3000, a(22) => N2999, a(21) => 
                           N2998, a(20) => N2997, a(19) => N2996, a(18) => 
                           N2995, a(17) => N2994, a(16) => N2993, a(15) => 
                           N2992, a(14) => N2991, a(13) => N2990, a(12) => 
                           N2989, a(11) => N2988, a(10) => N2987, a(9) => N2986
                           , a(8) => N2985, a(7) => N2984, a(6) => N2983, a(5) 
                           => N2982, a(4) => N2981, a(3) => N2980, a(2) => 
                           N2979, a(1) => N2978, a(0) => N2977, b(31) => N3168,
                           b(30) => N3167, b(29) => N3166, b(28) => N3165, 
                           b(27) => N3164, b(26) => N3163, b(25) => N3162, 
                           b(24) => N3161, b(23) => N3160, b(22) => N3159, 
                           b(21) => N3158, b(20) => N3157, b(19) => N3156, 
                           b(18) => N3155, b(17) => N3154, b(16) => N3153, 
                           b(15) => N3152, b(14) => N3151, b(13) => N3150, 
                           b(12) => N3149, b(11) => N3148, b(10) => N3147, b(9)
                           => N3146, b(8) => N3145, b(7) => N3144, b(6) => 
                           N3143, b(5) => N3142, b(4) => N3141, b(3) => N3140, 
                           b(2) => N3139, b(1) => N3138, b(0) => N3137, 
                           product(63) => n_1224, product(62) => n_1225, 
                           product(61) => n_1226, product(60) => n_1227, 
                           product(59) => n_1228, product(58) => n_1229, 
                           product(57) => n_1230, product(56) => n_1231, 
                           product(55) => n_1232, product(54) => n_1233, 
                           product(53) => n_1234, product(52) => n_1235, 
                           product(51) => n_1236, product(50) => n_1237, 
                           product(49) => n_1238, product(48) => n_1239, 
                           product(47) => n_1240, product(46) => n_1241, 
                           product(45) => n_1242, product(44) => n_1243, 
                           product(43) => n_1244, product(42) => n_1245, 
                           product(41) => n_1246, product(40) => n_1247, 
                           product(39) => n_1248, product(38) => n_1249, 
                           product(37) => n_1250, product(36) => n_1251, 
                           product(35) => n_1252, product(34) => n_1253, 
                           product(33) => n_1254, product(32) => n_1255, 
                           product(31) => N3328, product(30) => N3327, 
                           product(29) => N3326, product(28) => N3325, 
                           product(27) => N3324, product(26) => N3323, 
                           product(25) => N3322, product(24) => N3321, 
                           product(23) => N3320, product(22) => N3319, 
                           product(21) => N3318, product(20) => N3317, 
                           product(19) => N3316, product(18) => N3315, 
                           product(17) => N3314, product(16) => N3313, 
                           product(15) => N3312, product(14) => N3311, 
                           product(13) => N3310, product(12) => N3309, 
                           product(11) => N3308, product(10) => N3307, 
                           product(9) => N3306, product(8) => N3305, product(7)
                           => N3304, product(6) => N3303, product(5) => N3302, 
                           product(4) => N3301, product(3) => N3300, product(2)
                           => N3299, product(1) => N3298, product(0) => N3297);
   mult_21_C247 : gp_custom_DW_mult_tc_1 port map( a(31) => N3040, a(30) => 
                           N3039, a(29) => N3038, a(28) => N3037, a(27) => 
                           N3036, a(26) => N3035, a(25) => N3034, a(24) => 
                           N3033, a(23) => N3032, a(22) => N3031, a(21) => 
                           N3030, a(20) => N3029, a(19) => N3028, a(18) => 
                           N3027, a(17) => N3026, a(16) => N3025, a(15) => 
                           N3024, a(14) => N3023, a(13) => N3022, a(12) => 
                           N3021, a(11) => N3020, a(10) => N3019, a(9) => N3018
                           , a(8) => N3017, a(7) => N3016, a(6) => N3015, a(5) 
                           => N3014, a(4) => N3013, a(3) => N3012, a(2) => 
                           N3011, a(1) => N3010, a(0) => N3009, b(31) => N3232,
                           b(30) => N3231, b(29) => N3230, b(28) => N3229, 
                           b(27) => N3228, b(26) => N3227, b(25) => N3226, 
                           b(24) => N3225, b(23) => N3224, b(22) => N3223, 
                           b(21) => N3222, b(20) => N3221, b(19) => N3220, 
                           b(18) => N3219, b(17) => N3218, b(16) => N3217, 
                           b(15) => N3216, b(14) => N3215, b(13) => N3214, 
                           b(12) => N3213, b(11) => N3212, b(10) => N3211, b(9)
                           => N3210, b(8) => N3209, b(7) => N3208, b(6) => 
                           N3207, b(5) => N3206, b(4) => N3205, b(3) => N3204, 
                           b(2) => N3203, b(1) => N3202, b(0) => N3201, 
                           product(63) => n_1256, product(62) => n_1257, 
                           product(61) => n_1258, product(60) => n_1259, 
                           product(59) => n_1260, product(58) => n_1261, 
                           product(57) => n_1262, product(56) => n_1263, 
                           product(55) => n_1264, product(54) => n_1265, 
                           product(53) => n_1266, product(52) => n_1267, 
                           product(51) => n_1268, product(50) => n_1269, 
                           product(49) => n_1270, product(48) => n_1271, 
                           product(47) => n_1272, product(46) => n_1273, 
                           product(45) => n_1274, product(44) => n_1275, 
                           product(43) => n_1276, product(42) => n_1277, 
                           product(41) => n_1278, product(40) => n_1279, 
                           product(39) => n_1280, product(38) => n_1281, 
                           product(37) => n_1282, product(36) => n_1283, 
                           product(35) => n_1284, product(34) => n_1285, 
                           product(33) => n_1286, product(32) => n_1287, 
                           product(31) => N3360, product(30) => N3359, 
                           product(29) => N3358, product(28) => N3357, 
                           product(27) => N3356, product(26) => N3355, 
                           product(25) => N3354, product(24) => N3353, 
                           product(23) => N3352, product(22) => N3351, 
                           product(21) => N3350, product(20) => N3349, 
                           product(19) => N3348, product(18) => N3347, 
                           product(17) => N3346, product(16) => N3345, 
                           product(15) => N3344, product(14) => N3343, 
                           product(13) => N3342, product(12) => N3341, 
                           product(11) => N3340, product(10) => N3339, 
                           product(9) => N3338, product(8) => N3337, product(7)
                           => N3336, product(6) => N3335, product(5) => N3334, 
                           product(4) => N3333, product(3) => N3332, product(2)
                           => N3331, product(1) => N3330, product(0) => N3329);
   mult_21_C249 : gp_custom_DW_mult_tc_0 port map( a(31) => N3072, a(30) => 
                           N3071, a(29) => N3070, a(28) => N3069, a(27) => 
                           N3068, a(26) => N3067, a(25) => N3066, a(24) => 
                           N3065, a(23) => N3064, a(22) => N3063, a(21) => 
                           N3062, a(20) => N3061, a(19) => N3060, a(18) => 
                           N3059, a(17) => N3058, a(16) => N3057, a(15) => 
                           N3056, a(14) => N3055, a(13) => N3054, a(12) => 
                           N3053, a(11) => N3052, a(10) => N3051, a(9) => N3050
                           , a(8) => N3049, a(7) => N3048, a(6) => N3047, a(5) 
                           => N3046, a(4) => N3045, a(3) => N3044, a(2) => 
                           N3043, a(1) => N3042, a(0) => N3041, b(31) => N3232,
                           b(30) => N3231, b(29) => N3230, b(28) => N3229, 
                           b(27) => N3228, b(26) => N3227, b(25) => N3226, 
                           b(24) => N3225, b(23) => N3224, b(22) => N3223, 
                           b(21) => N3222, b(20) => N3221, b(19) => N3220, 
                           b(18) => N3219, b(17) => N3218, b(16) => N3217, 
                           b(15) => N3216, b(14) => N3215, b(13) => N3214, 
                           b(12) => N3213, b(11) => N3212, b(10) => N3211, b(9)
                           => N3210, b(8) => N3209, b(7) => N3208, b(6) => 
                           N3207, b(5) => N3206, b(4) => N3205, b(3) => N3204, 
                           b(2) => N3203, b(1) => N3202, b(0) => N3201, 
                           product(63) => n_1288, product(62) => n_1289, 
                           product(61) => n_1290, product(60) => n_1291, 
                           product(59) => n_1292, product(58) => n_1293, 
                           product(57) => n_1294, product(56) => n_1295, 
                           product(55) => n_1296, product(54) => n_1297, 
                           product(53) => n_1298, product(52) => n_1299, 
                           product(51) => n_1300, product(50) => n_1301, 
                           product(49) => n_1302, product(48) => n_1303, 
                           product(47) => n_1304, product(46) => n_1305, 
                           product(45) => n_1306, product(44) => n_1307, 
                           product(43) => n_1308, product(42) => n_1309, 
                           product(41) => n_1310, product(40) => n_1311, 
                           product(39) => n_1312, product(38) => n_1313, 
                           product(37) => n_1314, product(36) => n_1315, 
                           product(35) => n_1316, product(34) => n_1317, 
                           product(33) => n_1318, product(32) => n_1319, 
                           product(31) => N3392, product(30) => N3391, 
                           product(29) => N3390, product(28) => N3389, 
                           product(27) => N3388, product(26) => N3387, 
                           product(25) => N3386, product(24) => N3385, 
                           product(23) => N3384, product(22) => N3383, 
                           product(21) => N3382, product(20) => N3381, 
                           product(19) => N3380, product(18) => N3379, 
                           product(17) => N3378, product(16) => N3377, 
                           product(15) => N3376, product(14) => N3375, 
                           product(13) => N3374, product(12) => N3373, 
                           product(11) => N3372, product(10) => N3371, 
                           product(9) => N3370, product(8) => N3369, product(7)
                           => N3368, product(6) => N3367, product(5) => N3366, 
                           product(4) => N3365, product(3) => N3364, product(2)
                           => N3363, product(1) => N3362, product(0) => N3361);
   comp_res_reg_4_30_inst : DFFRPQ1 port map( D => N3391, CK => clk, RB => 
                           resetn, Q => comp_res_30_port);
   comp_res_reg_4_28_inst : DFFRPQ1 port map( D => N3389, CK => clk, RB => 
                           resetn, Q => comp_res_28_port);
   comp_res_reg_4_26_inst : DFFRPQ1 port map( D => N3387, CK => clk, RB => 
                           resetn, Q => comp_res_26_port);
   comp_res_reg_4_24_inst : DFFRPQ1 port map( D => N3385, CK => clk, RB => 
                           resetn, Q => comp_res_24_port);
   comp_res_reg_4_22_inst : DFFRPQ1 port map( D => N3383, CK => clk, RB => 
                           resetn, Q => comp_res_22_port);
   comp_res_reg_4_20_inst : DFFRPQ1 port map( D => N3381, CK => clk, RB => 
                           resetn, Q => comp_res_20_port);
   comp_res_reg_4_18_inst : DFFRPQ1 port map( D => N3379, CK => clk, RB => 
                           resetn, Q => comp_res_18_port);
   comp_res_reg_4_16_inst : DFFRPQ1 port map( D => N3377, CK => clk, RB => 
                           resetn, Q => comp_res_16_port);
   comp_res_reg_4_14_inst : DFFRPQ1 port map( D => N3375, CK => clk, RB => 
                           resetn, Q => comp_res_14_port);
   comp_res_reg_4_12_inst : DFFRPQ1 port map( D => N3373, CK => clk, RB => 
                           resetn, Q => comp_res_12_port);
   comp_res_reg_4_10_inst : DFFRPQ1 port map( D => N3371, CK => clk, RB => 
                           resetn, Q => comp_res_10_port);
   comp_res_reg_4_8_inst : DFFRPQ1 port map( D => N3369, CK => clk, RB => 
                           resetn, Q => comp_res_8_port);
   comp_res_reg_4_6_inst : DFFRPQ1 port map( D => N3367, CK => clk, RB => 
                           resetn, Q => comp_res_6_port);
   comp_res_reg_4_4_inst : DFFRPQ1 port map( D => N3365, CK => clk, RB => 
                           resetn, Q => comp_res_4_port);
   comp_res_reg_4_2_inst : DFFRPQ1 port map( D => N3363, CK => clk, RB => 
                           resetn, Q => comp_res_2_port);
   comp_res_reg_4_0_inst : DFFRPQ1 port map( D => N3361, CK => clk, RB => 
                           resetn, Q => comp_res_0_port);
   comp_res_reg_4_31_inst : DFFRPQ1 port map( D => N3392, CK => clk, RB => 
                           resetn, Q => comp_res_31_port);
   comp_res_reg_4_29_inst : DFFRPQ1 port map( D => N3390, CK => clk, RB => 
                           resetn, Q => comp_res_29_port);
   comp_res_reg_4_27_inst : DFFRPQ1 port map( D => N3388, CK => clk, RB => 
                           resetn, Q => comp_res_27_port);
   comp_res_reg_4_25_inst : DFFRPQ1 port map( D => N3386, CK => clk, RB => 
                           resetn, Q => comp_res_25_port);
   comp_res_reg_4_23_inst : DFFRPQ1 port map( D => N3384, CK => clk, RB => 
                           resetn, Q => comp_res_23_port);
   comp_res_reg_4_21_inst : DFFRPQ1 port map( D => N3382, CK => clk, RB => 
                           resetn, Q => comp_res_21_port);
   comp_res_reg_4_19_inst : DFFRPQ1 port map( D => N3380, CK => clk, RB => 
                           resetn, Q => comp_res_19_port);
   comp_res_reg_4_17_inst : DFFRPQ1 port map( D => N3378, CK => clk, RB => 
                           resetn, Q => comp_res_17_port);
   comp_res_reg_4_15_inst : DFFRPQ1 port map( D => N3376, CK => clk, RB => 
                           resetn, Q => comp_res_15_port);
   comp_res_reg_4_13_inst : DFFRPQ1 port map( D => N3374, CK => clk, RB => 
                           resetn, Q => comp_res_13_port);
   comp_res_reg_4_11_inst : DFFRPQ1 port map( D => N3372, CK => clk, RB => 
                           resetn, Q => comp_res_11_port);
   comp_res_reg_4_9_inst : DFFRPQ1 port map( D => N3370, CK => clk, RB => 
                           resetn, Q => comp_res_9_port);
   comp_res_reg_4_7_inst : DFFRPQ1 port map( D => N3368, CK => clk, RB => 
                           resetn, Q => comp_res_7_port);
   comp_res_reg_4_5_inst : DFFRPQ1 port map( D => N3366, CK => clk, RB => 
                           resetn, Q => comp_res_5_port);
   comp_res_reg_4_3_inst : DFFRPQ1 port map( D => N3364, CK => clk, RB => 
                           resetn, Q => comp_res_3_port);
   comp_res_reg_4_1_inst : DFFRPQ1 port map( D => N3362, CK => clk, RB => 
                           resetn, Q => comp_res_1_port);
   comp_res_reg_3_30_inst : DFFRPQ1 port map( D => N3359, CK => clk, RB => 
                           resetn, Q => comp_res_62_port);
   comp_res_reg_3_28_inst : DFFRPQ1 port map( D => N3357, CK => clk, RB => 
                           resetn, Q => comp_res_60_port);
   comp_res_reg_3_26_inst : DFFRPQ1 port map( D => N3355, CK => clk, RB => 
                           resetn, Q => comp_res_58_port);
   comp_res_reg_3_24_inst : DFFRPQ1 port map( D => N3353, CK => clk, RB => 
                           resetn, Q => comp_res_56_port);
   comp_res_reg_3_22_inst : DFFRPQ1 port map( D => N3351, CK => clk, RB => 
                           resetn, Q => comp_res_54_port);
   comp_res_reg_3_20_inst : DFFRPQ1 port map( D => N3349, CK => clk, RB => 
                           resetn, Q => comp_res_52_port);
   comp_res_reg_3_18_inst : DFFRPQ1 port map( D => N3347, CK => clk, RB => 
                           resetn, Q => comp_res_50_port);
   comp_res_reg_3_16_inst : DFFRPQ1 port map( D => N3345, CK => clk, RB => 
                           resetn, Q => comp_res_48_port);
   comp_res_reg_3_14_inst : DFFRPQ1 port map( D => N3343, CK => clk, RB => 
                           resetn, Q => comp_res_46_port);
   comp_res_reg_3_12_inst : DFFRPQ1 port map( D => N3341, CK => clk, RB => 
                           resetn, Q => comp_res_44_port);
   comp_res_reg_3_10_inst : DFFRPQ1 port map( D => N3339, CK => clk, RB => 
                           resetn, Q => comp_res_42_port);
   comp_res_reg_3_8_inst : DFFRPQ1 port map( D => N3337, CK => clk, RB => 
                           resetn, Q => comp_res_40_port);
   comp_res_reg_3_6_inst : DFFRPQ1 port map( D => N3335, CK => clk, RB => 
                           resetn, Q => comp_res_38_port);
   comp_res_reg_3_4_inst : DFFRPQ1 port map( D => N3333, CK => clk, RB => 
                           resetn, Q => comp_res_36_port);
   comp_res_reg_3_2_inst : DFFRPQ1 port map( D => N3331, CK => clk, RB => 
                           resetn, Q => comp_res_34_port);
   comp_res_reg_2_30_inst : DFFRPQ1 port map( D => N3327, CK => clk, RB => 
                           resetn, Q => comp_res_94_port);
   comp_res_reg_2_28_inst : DFFRPQ1 port map( D => N3325, CK => clk, RB => 
                           resetn, Q => comp_res_92_port);
   comp_res_reg_2_26_inst : DFFRPQ1 port map( D => N3323, CK => clk, RB => 
                           resetn, Q => comp_res_90_port);
   comp_res_reg_2_24_inst : DFFRPQ1 port map( D => N3321, CK => clk, RB => 
                           resetn, Q => comp_res_88_port);
   comp_res_reg_2_22_inst : DFFRPQ1 port map( D => N3319, CK => clk, RB => 
                           resetn, Q => comp_res_86_port);
   comp_res_reg_2_20_inst : DFFRPQ1 port map( D => N3317, CK => clk, RB => 
                           resetn, Q => comp_res_84_port);
   comp_res_reg_2_18_inst : DFFRPQ1 port map( D => N3315, CK => clk, RB => 
                           resetn, Q => comp_res_82_port);
   comp_res_reg_2_16_inst : DFFRPQ1 port map( D => N3313, CK => clk, RB => 
                           resetn, Q => comp_res_80_port);
   comp_res_reg_2_14_inst : DFFRPQ1 port map( D => N3311, CK => clk, RB => 
                           resetn, Q => comp_res_78_port);
   comp_res_reg_2_12_inst : DFFRPQ1 port map( D => N3309, CK => clk, RB => 
                           resetn, Q => comp_res_76_port);
   comp_res_reg_2_10_inst : DFFRPQ1 port map( D => N3307, CK => clk, RB => 
                           resetn, Q => comp_res_74_port);
   comp_res_reg_2_8_inst : DFFRPQ1 port map( D => N3305, CK => clk, RB => 
                           resetn, Q => comp_res_72_port);
   comp_res_reg_2_6_inst : DFFRPQ1 port map( D => N3303, CK => clk, RB => 
                           resetn, Q => comp_res_70_port);
   comp_res_reg_2_4_inst : DFFRPQ1 port map( D => N3301, CK => clk, RB => 
                           resetn, Q => comp_res_68_port);
   comp_res_reg_2_2_inst : DFFRPQ1 port map( D => N3299, CK => clk, RB => 
                           resetn, Q => comp_res_66_port);
   comp_res_reg_1_30_inst : DFFRPQ1 port map( D => N3295, CK => clk, RB => 
                           resetn, Q => comp_res_126_port);
   comp_res_reg_1_28_inst : DFFRPQ1 port map( D => N3293, CK => clk, RB => 
                           resetn, Q => comp_res_124_port);
   comp_res_reg_1_26_inst : DFFRPQ1 port map( D => N3291, CK => clk, RB => 
                           resetn, Q => comp_res_122_port);
   comp_res_reg_1_24_inst : DFFRPQ1 port map( D => N3289, CK => clk, RB => 
                           resetn, Q => comp_res_120_port);
   comp_res_reg_1_22_inst : DFFRPQ1 port map( D => N3287, CK => clk, RB => 
                           resetn, Q => comp_res_118_port);
   comp_res_reg_1_20_inst : DFFRPQ1 port map( D => N3285, CK => clk, RB => 
                           resetn, Q => comp_res_116_port);
   comp_res_reg_1_18_inst : DFFRPQ1 port map( D => N3283, CK => clk, RB => 
                           resetn, Q => comp_res_114_port);
   comp_res_reg_1_16_inst : DFFRPQ1 port map( D => N3281, CK => clk, RB => 
                           resetn, Q => comp_res_112_port);
   comp_res_reg_1_14_inst : DFFRPQ1 port map( D => N3279, CK => clk, RB => 
                           resetn, Q => comp_res_110_port);
   comp_res_reg_1_12_inst : DFFRPQ1 port map( D => N3277, CK => clk, RB => 
                           resetn, Q => comp_res_108_port);
   comp_res_reg_1_10_inst : DFFRPQ1 port map( D => N3275, CK => clk, RB => 
                           resetn, Q => comp_res_106_port);
   comp_res_reg_1_8_inst : DFFRPQ1 port map( D => N3273, CK => clk, RB => 
                           resetn, Q => comp_res_104_port);
   comp_res_reg_1_6_inst : DFFRPQ1 port map( D => N3271, CK => clk, RB => 
                           resetn, Q => comp_res_102_port);
   comp_res_reg_1_4_inst : DFFRPQ1 port map( D => N3269, CK => clk, RB => 
                           resetn, Q => comp_res_100_port);
   comp_res_reg_1_2_inst : DFFRPQ1 port map( D => N3267, CK => clk, RB => 
                           resetn, Q => comp_res_98_port);
   comp_res_reg_0_30_inst : DFFRPQ1 port map( D => N3263, CK => clk, RB => 
                           resetn, Q => comp_res_158_port);
   comp_res_reg_0_28_inst : DFFRPQ1 port map( D => N3261, CK => clk, RB => 
                           resetn, Q => comp_res_156_port);
   comp_res_reg_0_26_inst : DFFRPQ1 port map( D => N3259, CK => clk, RB => 
                           resetn, Q => comp_res_154_port);
   comp_res_reg_0_24_inst : DFFRPQ1 port map( D => N3257, CK => clk, RB => 
                           resetn, Q => comp_res_152_port);
   comp_res_reg_0_22_inst : DFFRPQ1 port map( D => N3255, CK => clk, RB => 
                           resetn, Q => comp_res_150_port);
   comp_res_reg_0_20_inst : DFFRPQ1 port map( D => N3253, CK => clk, RB => 
                           resetn, Q => comp_res_148_port);
   comp_res_reg_0_18_inst : DFFRPQ1 port map( D => N3251, CK => clk, RB => 
                           resetn, Q => comp_res_146_port);
   comp_res_reg_0_16_inst : DFFRPQ1 port map( D => N3249, CK => clk, RB => 
                           resetn, Q => comp_res_144_port);
   comp_res_reg_0_14_inst : DFFRPQ1 port map( D => N3247, CK => clk, RB => 
                           resetn, Q => comp_res_142_port);
   comp_res_reg_0_12_inst : DFFRPQ1 port map( D => N3245, CK => clk, RB => 
                           resetn, Q => comp_res_140_port);
   comp_res_reg_0_10_inst : DFFRPQ1 port map( D => N3243, CK => clk, RB => 
                           resetn, Q => comp_res_138_port);
   comp_res_reg_0_8_inst : DFFRPQ1 port map( D => N3241, CK => clk, RB => 
                           resetn, Q => comp_res_136_port);
   comp_res_reg_0_6_inst : DFFRPQ1 port map( D => N3239, CK => clk, RB => 
                           resetn, Q => comp_res_134_port);
   comp_res_reg_0_4_inst : DFFRPQ1 port map( D => N3237, CK => clk, RB => 
                           resetn, Q => comp_res_132_port);
   comp_res_reg_0_2_inst : DFFRPQ1 port map( D => N3235, CK => clk, RB => 
                           resetn, Q => comp_res_130_port);
   comp_res_reg_3_0_inst : DFFRPQ1 port map( D => N3329, CK => clk, RB => 
                           resetn, Q => comp_res_32_port);
   comp_res_reg_2_0_inst : DFFRPQ1 port map( D => N3297, CK => clk, RB => 
                           resetn, Q => comp_res_64_port);
   comp_res_reg_1_0_inst : DFFRPQ1 port map( D => N3265, CK => clk, RB => 
                           resetn, Q => comp_res_96_port);
   comp_res_reg_0_0_inst : DFFRPQ1 port map( D => N3233, CK => clk, RB => 
                           resetn, Q => comp_res_128_port);
   in_buf_reg_7_31_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n176,
                           CK => clk, RB => resetn, Q => in_buf_31_port);
   in_buf_reg_7_29_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n176,
                           CK => clk, RB => resetn, Q => in_buf_29_port);
   in_buf_reg_7_27_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n176,
                           CK => clk, RB => resetn, Q => in_buf_27_port);
   in_buf_reg_7_25_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n176, 
                           CK => clk, RB => resetn, Q => in_buf_25_port);
   in_buf_reg_7_23_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n176, 
                           CK => clk, RB => resetn, Q => in_buf_23_port);
   in_buf_reg_7_21_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n176, 
                           CK => clk, RB => resetn, Q => in_buf_21_port);
   in_buf_reg_7_19_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n176, 
                           CK => clk, RB => resetn, Q => in_buf_19_port);
   in_buf_reg_7_17_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n176, 
                           CK => clk, RB => resetn, Q => in_buf_17_port);
   in_buf_reg_7_15_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n177,
                           CK => clk, RB => resetn, Q => in_buf_15_port);
   in_buf_reg_7_13_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n177,
                           CK => clk, RB => resetn, Q => in_buf_13_port);
   in_buf_reg_7_11_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n177,
                           CK => clk, RB => resetn, Q => in_buf_11_port);
   in_buf_reg_7_9_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n177, 
                           CK => clk, RB => resetn, Q => in_buf_9_port);
   in_buf_reg_7_7_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n177, 
                           CK => clk, RB => resetn, Q => in_buf_7_port);
   in_buf_reg_7_5_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n177, 
                           CK => clk, RB => resetn, Q => in_buf_5_port);
   in_buf_reg_7_3_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n177, 
                           CK => clk, RB => resetn, Q => in_buf_3_port);
   in_buf_reg_7_1_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n177, 
                           CK => clk, RB => resetn, Q => in_buf_1_port);
   comp_res_reg_3_31_inst : DFFRPQ1 port map( D => N3360, CK => clk, RB => 
                           resetn, Q => comp_res_63_port);
   comp_res_reg_3_29_inst : DFFRPQ1 port map( D => N3358, CK => clk, RB => 
                           resetn, Q => comp_res_61_port);
   comp_res_reg_3_27_inst : DFFRPQ1 port map( D => N3356, CK => clk, RB => 
                           resetn, Q => comp_res_59_port);
   comp_res_reg_3_25_inst : DFFRPQ1 port map( D => N3354, CK => clk, RB => 
                           resetn, Q => comp_res_57_port);
   comp_res_reg_3_23_inst : DFFRPQ1 port map( D => N3352, CK => clk, RB => 
                           resetn, Q => comp_res_55_port);
   comp_res_reg_3_21_inst : DFFRPQ1 port map( D => N3350, CK => clk, RB => 
                           resetn, Q => comp_res_53_port);
   comp_res_reg_3_19_inst : DFFRPQ1 port map( D => N3348, CK => clk, RB => 
                           resetn, Q => comp_res_51_port);
   comp_res_reg_3_17_inst : DFFRPQ1 port map( D => N3346, CK => clk, RB => 
                           resetn, Q => comp_res_49_port);
   comp_res_reg_3_15_inst : DFFRPQ1 port map( D => N3344, CK => clk, RB => 
                           resetn, Q => comp_res_47_port);
   comp_res_reg_3_13_inst : DFFRPQ1 port map( D => N3342, CK => clk, RB => 
                           resetn, Q => comp_res_45_port);
   comp_res_reg_3_11_inst : DFFRPQ1 port map( D => N3340, CK => clk, RB => 
                           resetn, Q => comp_res_43_port);
   comp_res_reg_3_9_inst : DFFRPQ1 port map( D => N3338, CK => clk, RB => 
                           resetn, Q => comp_res_41_port);
   comp_res_reg_3_7_inst : DFFRPQ1 port map( D => N3336, CK => clk, RB => 
                           resetn, Q => comp_res_39_port);
   comp_res_reg_3_5_inst : DFFRPQ1 port map( D => N3334, CK => clk, RB => 
                           resetn, Q => comp_res_37_port);
   comp_res_reg_3_3_inst : DFFRPQ1 port map( D => N3332, CK => clk, RB => 
                           resetn, Q => comp_res_35_port);
   comp_res_reg_3_1_inst : DFFRPQ1 port map( D => N3330, CK => clk, RB => 
                           resetn, Q => comp_res_33_port);
   comp_res_reg_2_31_inst : DFFRPQ1 port map( D => N3328, CK => clk, RB => 
                           resetn, Q => comp_res_95_port);
   comp_res_reg_2_29_inst : DFFRPQ1 port map( D => N3326, CK => clk, RB => 
                           resetn, Q => comp_res_93_port);
   comp_res_reg_2_27_inst : DFFRPQ1 port map( D => N3324, CK => clk, RB => 
                           resetn, Q => comp_res_91_port);
   comp_res_reg_2_25_inst : DFFRPQ1 port map( D => N3322, CK => clk, RB => 
                           resetn, Q => comp_res_89_port);
   comp_res_reg_2_23_inst : DFFRPQ1 port map( D => N3320, CK => clk, RB => 
                           resetn, Q => comp_res_87_port);
   comp_res_reg_2_21_inst : DFFRPQ1 port map( D => N3318, CK => clk, RB => 
                           resetn, Q => comp_res_85_port);
   comp_res_reg_2_19_inst : DFFRPQ1 port map( D => N3316, CK => clk, RB => 
                           resetn, Q => comp_res_83_port);
   comp_res_reg_2_17_inst : DFFRPQ1 port map( D => N3314, CK => clk, RB => 
                           resetn, Q => comp_res_81_port);
   comp_res_reg_2_15_inst : DFFRPQ1 port map( D => N3312, CK => clk, RB => 
                           resetn, Q => comp_res_79_port);
   comp_res_reg_2_13_inst : DFFRPQ1 port map( D => N3310, CK => clk, RB => 
                           resetn, Q => comp_res_77_port);
   comp_res_reg_2_11_inst : DFFRPQ1 port map( D => N3308, CK => clk, RB => 
                           resetn, Q => comp_res_75_port);
   comp_res_reg_2_9_inst : DFFRPQ1 port map( D => N3306, CK => clk, RB => 
                           resetn, Q => comp_res_73_port);
   comp_res_reg_2_7_inst : DFFRPQ1 port map( D => N3304, CK => clk, RB => 
                           resetn, Q => comp_res_71_port);
   comp_res_reg_2_5_inst : DFFRPQ1 port map( D => N3302, CK => clk, RB => 
                           resetn, Q => comp_res_69_port);
   comp_res_reg_2_3_inst : DFFRPQ1 port map( D => N3300, CK => clk, RB => 
                           resetn, Q => comp_res_67_port);
   comp_res_reg_2_1_inst : DFFRPQ1 port map( D => N3298, CK => clk, RB => 
                           resetn, Q => comp_res_65_port);
   in_buf_reg_3_31_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n168,
                           CK => clk, RB => resetn, Q => in_buf_159_port);
   in_buf_reg_3_29_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n168,
                           CK => clk, RB => resetn, Q => in_buf_157_port);
   in_buf_reg_3_27_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n168,
                           CK => clk, RB => resetn, Q => in_buf_155_port);
   in_buf_reg_3_25_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n168, 
                           CK => clk, RB => resetn, Q => in_buf_153_port);
   in_buf_reg_3_23_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n168, 
                           CK => clk, RB => resetn, Q => in_buf_151_port);
   in_buf_reg_3_21_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n168, 
                           CK => clk, RB => resetn, Q => in_buf_149_port);
   in_buf_reg_3_19_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n168, 
                           CK => clk, RB => resetn, Q => in_buf_147_port);
   in_buf_reg_3_17_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n168, 
                           CK => clk, RB => resetn, Q => in_buf_145_port);
   in_buf_reg_3_15_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n169,
                           CK => clk, RB => resetn, Q => in_buf_143_port);
   in_buf_reg_3_13_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n169,
                           CK => clk, RB => resetn, Q => in_buf_141_port);
   in_buf_reg_3_11_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n169,
                           CK => clk, RB => resetn, Q => in_buf_139_port);
   in_buf_reg_3_9_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n169, 
                           CK => clk, RB => resetn, Q => in_buf_137_port);
   in_buf_reg_3_7_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n169, 
                           CK => clk, RB => resetn, Q => in_buf_135_port);
   in_buf_reg_3_5_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n169, 
                           CK => clk, RB => resetn, Q => in_buf_133_port);
   in_buf_reg_3_3_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n169, 
                           CK => clk, RB => resetn, Q => in_buf_131_port);
   in_buf_reg_3_1_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n169, 
                           CK => clk, RB => resetn, Q => in_buf_129_port);
   in_buf_reg_2_31_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n166,
                           CK => clk, RB => resetn, Q => in_buf_191_port);
   in_buf_reg_2_29_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n166,
                           CK => clk, RB => resetn, Q => in_buf_189_port);
   in_buf_reg_2_27_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n166,
                           CK => clk, RB => resetn, Q => in_buf_187_port);
   in_buf_reg_2_25_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n166, 
                           CK => clk, RB => resetn, Q => in_buf_185_port);
   in_buf_reg_2_23_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n166, 
                           CK => clk, RB => resetn, Q => in_buf_183_port);
   in_buf_reg_2_21_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n166, 
                           CK => clk, RB => resetn, Q => in_buf_181_port);
   in_buf_reg_2_19_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n166, 
                           CK => clk, RB => resetn, Q => in_buf_179_port);
   in_buf_reg_2_17_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n166, 
                           CK => clk, RB => resetn, Q => in_buf_177_port);
   in_buf_reg_6_31_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n174,
                           CK => clk, RB => resetn, Q => in_buf_63_port);
   in_buf_reg_6_29_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n174,
                           CK => clk, RB => resetn, Q => in_buf_61_port);
   in_buf_reg_6_27_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n174,
                           CK => clk, RB => resetn, Q => in_buf_59_port);
   in_buf_reg_6_25_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n174, 
                           CK => clk, RB => resetn, Q => in_buf_57_port);
   in_buf_reg_6_23_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n174, 
                           CK => clk, RB => resetn, Q => in_buf_55_port);
   in_buf_reg_6_21_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n174, 
                           CK => clk, RB => resetn, Q => in_buf_53_port);
   in_buf_reg_6_19_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n174, 
                           CK => clk, RB => resetn, Q => in_buf_51_port);
   in_buf_reg_6_17_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n174, 
                           CK => clk, RB => resetn, Q => in_buf_49_port);
   in_buf_reg_2_15_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n167,
                           CK => clk, RB => resetn, Q => in_buf_175_port);
   in_buf_reg_2_13_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n167,
                           CK => clk, RB => resetn, Q => in_buf_173_port);
   in_buf_reg_2_11_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n167,
                           CK => clk, RB => resetn, Q => in_buf_171_port);
   in_buf_reg_2_9_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n167, 
                           CK => clk, RB => resetn, Q => in_buf_169_port);
   in_buf_reg_2_7_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n167, 
                           CK => clk, RB => resetn, Q => in_buf_167_port);
   in_buf_reg_2_5_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n167, 
                           CK => clk, RB => resetn, Q => in_buf_165_port);
   in_buf_reg_2_3_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n167, 
                           CK => clk, RB => resetn, Q => in_buf_163_port);
   in_buf_reg_2_1_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n167, 
                           CK => clk, RB => resetn, Q => in_buf_161_port);
   in_buf_reg_6_15_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n175,
                           CK => clk, RB => resetn, Q => in_buf_47_port);
   in_buf_reg_6_13_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n175,
                           CK => clk, RB => resetn, Q => in_buf_45_port);
   in_buf_reg_6_11_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n175,
                           CK => clk, RB => resetn, Q => in_buf_43_port);
   in_buf_reg_6_9_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n175, 
                           CK => clk, RB => resetn, Q => in_buf_41_port);
   in_buf_reg_6_7_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n175, 
                           CK => clk, RB => resetn, Q => in_buf_39_port);
   in_buf_reg_6_5_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n175, 
                           CK => clk, RB => resetn, Q => in_buf_37_port);
   in_buf_reg_6_3_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n175, 
                           CK => clk, RB => resetn, Q => in_buf_35_port);
   in_buf_reg_6_1_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n175, 
                           CK => clk, RB => resetn, Q => in_buf_33_port);
   in_buf_reg_5_31_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n172,
                           CK => clk, RB => resetn, Q => in_buf_95_port);
   in_buf_reg_5_29_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n172,
                           CK => clk, RB => resetn, Q => in_buf_93_port);
   in_buf_reg_5_27_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n172,
                           CK => clk, RB => resetn, Q => in_buf_91_port);
   in_buf_reg_5_25_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n172, 
                           CK => clk, RB => resetn, Q => in_buf_89_port);
   in_buf_reg_5_23_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n172, 
                           CK => clk, RB => resetn, Q => in_buf_87_port);
   in_buf_reg_5_21_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n172, 
                           CK => clk, RB => resetn, Q => in_buf_85_port);
   in_buf_reg_5_19_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n172, 
                           CK => clk, RB => resetn, Q => in_buf_83_port);
   in_buf_reg_5_17_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n172, 
                           CK => clk, RB => resetn, Q => in_buf_81_port);
   in_buf_reg_5_15_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n173,
                           CK => clk, RB => resetn, Q => in_buf_79_port);
   in_buf_reg_5_13_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n173,
                           CK => clk, RB => resetn, Q => in_buf_77_port);
   in_buf_reg_5_11_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n173,
                           CK => clk, RB => resetn, Q => in_buf_75_port);
   in_buf_reg_5_9_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n173, 
                           CK => clk, RB => resetn, Q => in_buf_73_port);
   in_buf_reg_5_7_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n173, 
                           CK => clk, RB => resetn, Q => in_buf_71_port);
   in_buf_reg_5_5_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n173, 
                           CK => clk, RB => resetn, Q => in_buf_69_port);
   in_buf_reg_5_3_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n173, 
                           CK => clk, RB => resetn, Q => in_buf_67_port);
   in_buf_reg_5_1_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n173, 
                           CK => clk, RB => resetn, Q => in_buf_65_port);
   comp_res_reg_1_31_inst : DFFRPQ1 port map( D => N3296, CK => clk, RB => 
                           resetn, Q => comp_res_127_port);
   comp_res_reg_1_29_inst : DFFRPQ1 port map( D => N3294, CK => clk, RB => 
                           resetn, Q => comp_res_125_port);
   comp_res_reg_1_27_inst : DFFRPQ1 port map( D => N3292, CK => clk, RB => 
                           resetn, Q => comp_res_123_port);
   comp_res_reg_1_25_inst : DFFRPQ1 port map( D => N3290, CK => clk, RB => 
                           resetn, Q => comp_res_121_port);
   comp_res_reg_1_23_inst : DFFRPQ1 port map( D => N3288, CK => clk, RB => 
                           resetn, Q => comp_res_119_port);
   comp_res_reg_1_21_inst : DFFRPQ1 port map( D => N3286, CK => clk, RB => 
                           resetn, Q => comp_res_117_port);
   comp_res_reg_1_19_inst : DFFRPQ1 port map( D => N3284, CK => clk, RB => 
                           resetn, Q => comp_res_115_port);
   comp_res_reg_1_17_inst : DFFRPQ1 port map( D => N3282, CK => clk, RB => 
                           resetn, Q => comp_res_113_port);
   comp_res_reg_1_15_inst : DFFRPQ1 port map( D => N3280, CK => clk, RB => 
                           resetn, Q => comp_res_111_port);
   comp_res_reg_1_13_inst : DFFRPQ1 port map( D => N3278, CK => clk, RB => 
                           resetn, Q => comp_res_109_port);
   comp_res_reg_1_11_inst : DFFRPQ1 port map( D => N3276, CK => clk, RB => 
                           resetn, Q => comp_res_107_port);
   comp_res_reg_1_9_inst : DFFRPQ1 port map( D => N3274, CK => clk, RB => 
                           resetn, Q => comp_res_105_port);
   comp_res_reg_1_7_inst : DFFRPQ1 port map( D => N3272, CK => clk, RB => 
                           resetn, Q => comp_res_103_port);
   comp_res_reg_1_5_inst : DFFRPQ1 port map( D => N3270, CK => clk, RB => 
                           resetn, Q => comp_res_101_port);
   comp_res_reg_1_3_inst : DFFRPQ1 port map( D => N3268, CK => clk, RB => 
                           resetn, Q => comp_res_99_port);
   comp_res_reg_1_1_inst : DFFRPQ1 port map( D => N3266, CK => clk, RB => 
                           resetn, Q => comp_res_97_port);
   comp_res_reg_0_31_inst : DFFRPQ1 port map( D => N3264, CK => clk, RB => 
                           resetn, Q => comp_res_159_port);
   comp_res_reg_0_29_inst : DFFRPQ1 port map( D => N3262, CK => clk, RB => 
                           resetn, Q => comp_res_157_port);
   comp_res_reg_0_27_inst : DFFRPQ1 port map( D => N3260, CK => clk, RB => 
                           resetn, Q => comp_res_155_port);
   comp_res_reg_0_25_inst : DFFRPQ1 port map( D => N3258, CK => clk, RB => 
                           resetn, Q => comp_res_153_port);
   comp_res_reg_0_23_inst : DFFRPQ1 port map( D => N3256, CK => clk, RB => 
                           resetn, Q => comp_res_151_port);
   comp_res_reg_0_21_inst : DFFRPQ1 port map( D => N3254, CK => clk, RB => 
                           resetn, Q => comp_res_149_port);
   comp_res_reg_0_19_inst : DFFRPQ1 port map( D => N3252, CK => clk, RB => 
                           resetn, Q => comp_res_147_port);
   comp_res_reg_0_17_inst : DFFRPQ1 port map( D => N3250, CK => clk, RB => 
                           resetn, Q => comp_res_145_port);
   comp_res_reg_0_15_inst : DFFRPQ1 port map( D => N3248, CK => clk, RB => 
                           resetn, Q => comp_res_143_port);
   comp_res_reg_0_13_inst : DFFRPQ1 port map( D => N3246, CK => clk, RB => 
                           resetn, Q => comp_res_141_port);
   comp_res_reg_0_11_inst : DFFRPQ1 port map( D => N3244, CK => clk, RB => 
                           resetn, Q => comp_res_139_port);
   comp_res_reg_0_9_inst : DFFRPQ1 port map( D => N3242, CK => clk, RB => 
                           resetn, Q => comp_res_137_port);
   comp_res_reg_0_7_inst : DFFRPQ1 port map( D => N3240, CK => clk, RB => 
                           resetn, Q => comp_res_135_port);
   comp_res_reg_0_5_inst : DFFRPQ1 port map( D => N3238, CK => clk, RB => 
                           resetn, Q => comp_res_133_port);
   comp_res_reg_0_3_inst : DFFRPQ1 port map( D => N3236, CK => clk, RB => 
                           resetn, Q => comp_res_131_port);
   comp_res_reg_0_1_inst : DFFRPQ1 port map( D => N3234, CK => clk, RB => 
                           resetn, Q => comp_res_129_port);
   in_buf_reg_1_31_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n164,
                           CK => clk, RB => resetn, Q => in_buf_223_port);
   in_buf_reg_1_29_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n164,
                           CK => clk, RB => resetn, Q => in_buf_221_port);
   in_buf_reg_1_27_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n164,
                           CK => clk, RB => resetn, Q => in_buf_219_port);
   in_buf_reg_1_25_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n164, 
                           CK => clk, RB => resetn, Q => in_buf_217_port);
   in_buf_reg_1_23_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n164, 
                           CK => clk, RB => resetn, Q => in_buf_215_port);
   in_buf_reg_1_21_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n164, 
                           CK => clk, RB => resetn, Q => in_buf_213_port);
   in_buf_reg_1_19_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n164, 
                           CK => clk, RB => resetn, Q => in_buf_211_port);
   in_buf_reg_1_17_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n164, 
                           CK => clk, RB => resetn, Q => in_buf_209_port);
   in_buf_reg_1_15_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n165,
                           CK => clk, RB => resetn, Q => in_buf_207_port);
   in_buf_reg_1_13_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n165,
                           CK => clk, RB => resetn, Q => in_buf_205_port);
   in_buf_reg_1_11_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n165,
                           CK => clk, RB => resetn, Q => in_buf_203_port);
   in_buf_reg_1_9_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n165, 
                           CK => clk, RB => resetn, Q => in_buf_201_port);
   in_buf_reg_1_7_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n165, 
                           CK => clk, RB => resetn, Q => in_buf_199_port);
   in_buf_reg_1_5_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n165, 
                           CK => clk, RB => resetn, Q => in_buf_197_port);
   in_buf_reg_1_3_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n165, 
                           CK => clk, RB => resetn, Q => in_buf_195_port);
   in_buf_reg_1_1_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n165, 
                           CK => clk, RB => resetn, Q => in_buf_193_port);
   in_buf_reg_4_31_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n170,
                           CK => clk, RB => resetn, Q => in_buf_127_port);
   in_buf_reg_4_29_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n170,
                           CK => clk, RB => resetn, Q => in_buf_125_port);
   in_buf_reg_4_27_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n170,
                           CK => clk, RB => resetn, Q => in_buf_123_port);
   in_buf_reg_4_25_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n170, 
                           CK => clk, RB => resetn, Q => in_buf_121_port);
   in_buf_reg_4_23_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n170, 
                           CK => clk, RB => resetn, Q => in_buf_119_port);
   in_buf_reg_4_21_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n170, 
                           CK => clk, RB => resetn, Q => in_buf_117_port);
   in_buf_reg_4_19_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n170, 
                           CK => clk, RB => resetn, Q => in_buf_115_port);
   in_buf_reg_4_17_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n170, 
                           CK => clk, RB => resetn, Q => in_buf_113_port);
   in_buf_reg_0_31_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n162,
                           CK => clk, RB => resetn, Q => in_buf_255_port);
   in_buf_reg_0_29_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n162,
                           CK => clk, RB => resetn, Q => in_buf_253_port);
   in_buf_reg_0_27_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n162,
                           CK => clk, RB => resetn, Q => in_buf_251_port);
   in_buf_reg_0_25_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n162, 
                           CK => clk, RB => resetn, Q => in_buf_249_port);
   in_buf_reg_0_23_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n162, 
                           CK => clk, RB => resetn, Q => in_buf_247_port);
   in_buf_reg_0_21_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n162, 
                           CK => clk, RB => resetn, Q => in_buf_245_port);
   in_buf_reg_0_19_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n162, 
                           CK => clk, RB => resetn, Q => in_buf_243_port);
   in_buf_reg_0_17_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n162, 
                           CK => clk, RB => resetn, Q => in_buf_241_port);
   in_buf_reg_0_15_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n163,
                           CK => clk, RB => resetn, Q => in_buf_239_port);
   in_buf_reg_0_13_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n163,
                           CK => clk, RB => resetn, Q => in_buf_237_port);
   in_buf_reg_0_11_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n163,
                           CK => clk, RB => resetn, Q => in_buf_235_port);
   in_buf_reg_0_9_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n163, 
                           CK => clk, RB => resetn, Q => in_buf_233_port);
   in_buf_reg_0_7_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n163, 
                           CK => clk, RB => resetn, Q => in_buf_231_port);
   in_buf_reg_0_5_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n163, 
                           CK => clk, RB => resetn, Q => in_buf_229_port);
   in_buf_reg_0_3_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n163, 
                           CK => clk, RB => resetn, Q => in_buf_227_port);
   in_buf_reg_0_1_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n163, 
                           CK => clk, RB => resetn, Q => in_buf_225_port);
   in_buf_reg_4_15_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n171,
                           CK => clk, RB => resetn, Q => in_buf_111_port);
   in_buf_reg_4_13_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n171,
                           CK => clk, RB => resetn, Q => in_buf_109_port);
   in_buf_reg_4_11_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n171,
                           CK => clk, RB => resetn, Q => in_buf_107_port);
   in_buf_reg_4_9_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n171, 
                           CK => clk, RB => resetn, Q => in_buf_105_port);
   in_buf_reg_4_7_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n171, 
                           CK => clk, RB => resetn, Q => in_buf_103_port);
   in_buf_reg_4_5_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n171, 
                           CK => clk, RB => resetn, Q => in_buf_101_port);
   in_buf_reg_4_3_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n171, 
                           CK => clk, RB => resetn, Q => in_buf_99_port);
   in_buf_reg_4_1_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n171, 
                           CK => clk, RB => resetn, Q => in_buf_97_port);
   in_buf_reg_7_30_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n176,
                           CK => clk, RB => resetn, Q => in_buf_30_port);
   in_buf_reg_7_28_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n176,
                           CK => clk, RB => resetn, Q => in_buf_28_port);
   in_buf_reg_7_26_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n176,
                           CK => clk, RB => resetn, Q => in_buf_26_port);
   in_buf_reg_7_24_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n176, 
                           CK => clk, RB => resetn, Q => in_buf_24_port);
   in_buf_reg_7_22_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n176, 
                           CK => clk, RB => resetn, Q => in_buf_22_port);
   in_buf_reg_7_20_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n176, 
                           CK => clk, RB => resetn, Q => in_buf_20_port);
   in_buf_reg_7_18_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n176, 
                           CK => clk, RB => resetn, Q => in_buf_18_port);
   in_buf_reg_7_16_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n176, 
                           CK => clk, RB => resetn, Q => in_buf_16_port);
   in_buf_reg_7_14_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n177,
                           CK => clk, RB => resetn, Q => in_buf_14_port);
   in_buf_reg_7_12_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n177,
                           CK => clk, RB => resetn, Q => in_buf_12_port);
   in_buf_reg_7_10_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n177,
                           CK => clk, RB => resetn, Q => in_buf_10_port);
   in_buf_reg_7_8_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n177, 
                           CK => clk, RB => resetn, Q => in_buf_8_port);
   in_buf_reg_7_6_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n177, 
                           CK => clk, RB => resetn, Q => in_buf_6_port);
   in_buf_reg_7_4_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n177, 
                           CK => clk, RB => resetn, Q => in_buf_4_port);
   in_buf_reg_7_2_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n177, 
                           CK => clk, RB => resetn, Q => in_buf_2_port);
   in_trigger_reg : DFFRPQ1 port map( D => n241, CK => clk, RB => resetn, Q => 
                           in_trigger);
   in_buf_reg_3_30_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n168,
                           CK => clk, RB => resetn, Q => in_buf_158_port);
   in_buf_reg_3_28_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n168,
                           CK => clk, RB => resetn, Q => in_buf_156_port);
   in_buf_reg_3_26_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n168,
                           CK => clk, RB => resetn, Q => in_buf_154_port);
   in_buf_reg_3_24_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n168, 
                           CK => clk, RB => resetn, Q => in_buf_152_port);
   in_buf_reg_3_22_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n168, 
                           CK => clk, RB => resetn, Q => in_buf_150_port);
   in_buf_reg_3_20_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n168, 
                           CK => clk, RB => resetn, Q => in_buf_148_port);
   in_buf_reg_3_18_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n168, 
                           CK => clk, RB => resetn, Q => in_buf_146_port);
   in_buf_reg_3_16_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n168, 
                           CK => clk, RB => resetn, Q => in_buf_144_port);
   in_buf_reg_3_14_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n169,
                           CK => clk, RB => resetn, Q => in_buf_142_port);
   in_buf_reg_3_12_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n169,
                           CK => clk, RB => resetn, Q => in_buf_140_port);
   in_buf_reg_3_10_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n169,
                           CK => clk, RB => resetn, Q => in_buf_138_port);
   in_buf_reg_3_8_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n169, 
                           CK => clk, RB => resetn, Q => in_buf_136_port);
   in_buf_reg_3_6_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n169, 
                           CK => clk, RB => resetn, Q => in_buf_134_port);
   in_buf_reg_3_4_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n169, 
                           CK => clk, RB => resetn, Q => in_buf_132_port);
   in_buf_reg_3_2_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n169, 
                           CK => clk, RB => resetn, Q => in_buf_130_port);
   in_buf_reg_2_30_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n166,
                           CK => clk, RB => resetn, Q => in_buf_190_port);
   in_buf_reg_2_28_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n166,
                           CK => clk, RB => resetn, Q => in_buf_188_port);
   in_buf_reg_2_26_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n166,
                           CK => clk, RB => resetn, Q => in_buf_186_port);
   in_buf_reg_2_24_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n166, 
                           CK => clk, RB => resetn, Q => in_buf_184_port);
   in_buf_reg_2_22_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n166, 
                           CK => clk, RB => resetn, Q => in_buf_182_port);
   in_buf_reg_2_20_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n166, 
                           CK => clk, RB => resetn, Q => in_buf_180_port);
   in_buf_reg_2_18_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n166, 
                           CK => clk, RB => resetn, Q => in_buf_178_port);
   in_buf_reg_2_16_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n166, 
                           CK => clk, RB => resetn, Q => in_buf_176_port);
   in_buf_reg_6_30_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n174,
                           CK => clk, RB => resetn, Q => in_buf_62_port);
   in_buf_reg_6_28_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n174,
                           CK => clk, RB => resetn, Q => in_buf_60_port);
   in_buf_reg_6_26_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n174,
                           CK => clk, RB => resetn, Q => in_buf_58_port);
   in_buf_reg_6_24_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n174, 
                           CK => clk, RB => resetn, Q => in_buf_56_port);
   in_buf_reg_6_22_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n174, 
                           CK => clk, RB => resetn, Q => in_buf_54_port);
   in_buf_reg_6_20_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n174, 
                           CK => clk, RB => resetn, Q => in_buf_52_port);
   in_buf_reg_6_18_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n174, 
                           CK => clk, RB => resetn, Q => in_buf_50_port);
   in_buf_reg_6_16_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n174, 
                           CK => clk, RB => resetn, Q => in_buf_48_port);
   in_buf_reg_2_14_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n167,
                           CK => clk, RB => resetn, Q => in_buf_174_port);
   in_buf_reg_2_12_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n167,
                           CK => clk, RB => resetn, Q => in_buf_172_port);
   in_buf_reg_2_10_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n167,
                           CK => clk, RB => resetn, Q => in_buf_170_port);
   in_buf_reg_2_8_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n167, 
                           CK => clk, RB => resetn, Q => in_buf_168_port);
   in_buf_reg_2_6_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n167, 
                           CK => clk, RB => resetn, Q => in_buf_166_port);
   in_buf_reg_2_4_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n167, 
                           CK => clk, RB => resetn, Q => in_buf_164_port);
   in_buf_reg_2_2_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n167, 
                           CK => clk, RB => resetn, Q => in_buf_162_port);
   in_buf_reg_6_14_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n175,
                           CK => clk, RB => resetn, Q => in_buf_46_port);
   in_buf_reg_6_12_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n175,
                           CK => clk, RB => resetn, Q => in_buf_44_port);
   in_buf_reg_6_10_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n175,
                           CK => clk, RB => resetn, Q => in_buf_42_port);
   in_buf_reg_6_8_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n175, 
                           CK => clk, RB => resetn, Q => in_buf_40_port);
   in_buf_reg_6_6_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n175, 
                           CK => clk, RB => resetn, Q => in_buf_38_port);
   in_buf_reg_6_4_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n175, 
                           CK => clk, RB => resetn, Q => in_buf_36_port);
   in_buf_reg_6_2_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n175, 
                           CK => clk, RB => resetn, Q => in_buf_34_port);
   in_buf_reg_5_30_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n172,
                           CK => clk, RB => resetn, Q => in_buf_94_port);
   in_buf_reg_5_28_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n172,
                           CK => clk, RB => resetn, Q => in_buf_92_port);
   in_buf_reg_5_26_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n172,
                           CK => clk, RB => resetn, Q => in_buf_90_port);
   in_buf_reg_5_24_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n172, 
                           CK => clk, RB => resetn, Q => in_buf_88_port);
   in_buf_reg_5_22_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n172, 
                           CK => clk, RB => resetn, Q => in_buf_86_port);
   in_buf_reg_5_20_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n172, 
                           CK => clk, RB => resetn, Q => in_buf_84_port);
   in_buf_reg_5_18_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n172, 
                           CK => clk, RB => resetn, Q => in_buf_82_port);
   in_buf_reg_5_16_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n172, 
                           CK => clk, RB => resetn, Q => in_buf_80_port);
   in_buf_reg_5_14_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n173,
                           CK => clk, RB => resetn, Q => in_buf_78_port);
   in_buf_reg_5_12_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n173,
                           CK => clk, RB => resetn, Q => in_buf_76_port);
   in_buf_reg_5_10_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n173,
                           CK => clk, RB => resetn, Q => in_buf_74_port);
   in_buf_reg_5_8_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n173, 
                           CK => clk, RB => resetn, Q => in_buf_72_port);
   in_buf_reg_5_6_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n173, 
                           CK => clk, RB => resetn, Q => in_buf_70_port);
   in_buf_reg_5_4_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n173, 
                           CK => clk, RB => resetn, Q => in_buf_68_port);
   in_buf_reg_5_2_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n173, 
                           CK => clk, RB => resetn, Q => in_buf_66_port);
   in_buf_reg_7_0_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n177, 
                           CK => clk, RB => resetn, Q => in_buf_0_port);
   in_buf_reg_1_30_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n164,
                           CK => clk, RB => resetn, Q => in_buf_222_port);
   in_buf_reg_1_28_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n164,
                           CK => clk, RB => resetn, Q => in_buf_220_port);
   in_buf_reg_1_26_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n164,
                           CK => clk, RB => resetn, Q => in_buf_218_port);
   in_buf_reg_1_24_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n164, 
                           CK => clk, RB => resetn, Q => in_buf_216_port);
   in_buf_reg_1_22_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n164, 
                           CK => clk, RB => resetn, Q => in_buf_214_port);
   in_buf_reg_1_20_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n164, 
                           CK => clk, RB => resetn, Q => in_buf_212_port);
   in_buf_reg_1_18_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n164, 
                           CK => clk, RB => resetn, Q => in_buf_210_port);
   in_buf_reg_1_16_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n164, 
                           CK => clk, RB => resetn, Q => in_buf_208_port);
   in_buf_reg_1_14_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n165,
                           CK => clk, RB => resetn, Q => in_buf_206_port);
   in_buf_reg_1_12_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n165,
                           CK => clk, RB => resetn, Q => in_buf_204_port);
   in_buf_reg_1_10_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n165,
                           CK => clk, RB => resetn, Q => in_buf_202_port);
   in_buf_reg_1_8_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n165, 
                           CK => clk, RB => resetn, Q => in_buf_200_port);
   in_buf_reg_1_6_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n165, 
                           CK => clk, RB => resetn, Q => in_buf_198_port);
   in_buf_reg_1_4_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n165, 
                           CK => clk, RB => resetn, Q => in_buf_196_port);
   in_buf_reg_1_2_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n165, 
                           CK => clk, RB => resetn, Q => in_buf_194_port);
   in_buf_reg_4_30_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n170,
                           CK => clk, RB => resetn, Q => in_buf_126_port);
   in_buf_reg_4_28_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n170,
                           CK => clk, RB => resetn, Q => in_buf_124_port);
   in_buf_reg_4_26_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n170,
                           CK => clk, RB => resetn, Q => in_buf_122_port);
   in_buf_reg_4_24_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n170, 
                           CK => clk, RB => resetn, Q => in_buf_120_port);
   in_buf_reg_4_22_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n170, 
                           CK => clk, RB => resetn, Q => in_buf_118_port);
   in_buf_reg_4_20_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n170, 
                           CK => clk, RB => resetn, Q => in_buf_116_port);
   in_buf_reg_4_18_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n170, 
                           CK => clk, RB => resetn, Q => in_buf_114_port);
   in_buf_reg_4_16_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n170, 
                           CK => clk, RB => resetn, Q => in_buf_112_port);
   in_buf_reg_0_30_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n162,
                           CK => clk, RB => resetn, Q => in_buf_254_port);
   in_buf_reg_0_28_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n162,
                           CK => clk, RB => resetn, Q => in_buf_252_port);
   in_buf_reg_0_26_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n162,
                           CK => clk, RB => resetn, Q => in_buf_250_port);
   in_buf_reg_0_24_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n162, 
                           CK => clk, RB => resetn, Q => in_buf_248_port);
   in_buf_reg_0_22_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n162, 
                           CK => clk, RB => resetn, Q => in_buf_246_port);
   in_buf_reg_0_20_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n162, 
                           CK => clk, RB => resetn, Q => in_buf_244_port);
   in_buf_reg_0_18_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n162, 
                           CK => clk, RB => resetn, Q => in_buf_242_port);
   in_buf_reg_0_16_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n162, 
                           CK => clk, RB => resetn, Q => in_buf_240_port);
   in_buf_reg_0_14_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n163,
                           CK => clk, RB => resetn, Q => in_buf_238_port);
   in_buf_reg_0_12_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n163,
                           CK => clk, RB => resetn, Q => in_buf_236_port);
   in_buf_reg_0_10_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n163,
                           CK => clk, RB => resetn, Q => in_buf_234_port);
   in_buf_reg_0_8_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n163, 
                           CK => clk, RB => resetn, Q => in_buf_232_port);
   in_buf_reg_0_6_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n163, 
                           CK => clk, RB => resetn, Q => in_buf_230_port);
   in_buf_reg_0_4_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n163, 
                           CK => clk, RB => resetn, Q => in_buf_228_port);
   in_buf_reg_0_2_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n163, 
                           CK => clk, RB => resetn, Q => in_buf_226_port);
   in_buf_reg_4_14_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n171,
                           CK => clk, RB => resetn, Q => in_buf_110_port);
   in_buf_reg_4_12_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n171,
                           CK => clk, RB => resetn, Q => in_buf_108_port);
   in_buf_reg_4_10_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n171,
                           CK => clk, RB => resetn, Q => in_buf_106_port);
   in_buf_reg_4_8_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n171, 
                           CK => clk, RB => resetn, Q => in_buf_104_port);
   in_buf_reg_4_6_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n171, 
                           CK => clk, RB => resetn, Q => in_buf_102_port);
   in_buf_reg_4_4_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n171, 
                           CK => clk, RB => resetn, Q => in_buf_100_port);
   in_buf_reg_4_2_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n171, 
                           CK => clk, RB => resetn, Q => in_buf_98_port);
   in_buf_reg_3_0_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n169, 
                           CK => clk, RB => resetn, Q => in_buf_128_port);
   in_buf_reg_2_0_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n167, 
                           CK => clk, RB => resetn, Q => in_buf_160_port);
   in_buf_reg_6_0_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n175, 
                           CK => clk, RB => resetn, Q => in_buf_32_port);
   in_buf_reg_5_0_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n173, 
                           CK => clk, RB => resetn, Q => in_buf_64_port);
   out_buf_reg_7_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n245, CK => clk, RB => resetn, Q => out_buf_15_port)
                           ;
   out_buf_reg_7_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n245, CK => clk, RB => resetn, Q => out_buf_14_port)
                           ;
   out_buf_reg_7_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n245, CK => clk, RB => resetn, Q => out_buf_13_port)
                           ;
   out_buf_reg_7_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n245, CK => clk, RB => resetn, Q => out_buf_12_port)
                           ;
   out_buf_reg_7_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n245, CK => clk, RB => resetn, Q => out_buf_11_port)
                           ;
   out_buf_reg_7_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n245, CK => clk, RB => resetn, Q => out_buf_10_port)
                           ;
   out_buf_reg_7_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => n245,
                           CK => clk, RB => resetn, Q => out_buf_9_port);
   out_buf_reg_7_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => n245,
                           CK => clk, RB => resetn, Q => out_buf_8_port);
   out_buf_reg_7_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => n245,
                           CK => clk, RB => resetn, Q => out_buf_7_port);
   out_buf_reg_7_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => n245,
                           CK => clk, RB => resetn, Q => out_buf_6_port);
   out_buf_reg_7_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => n245,
                           CK => clk, RB => resetn, Q => out_buf_5_port);
   out_buf_reg_7_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => n245,
                           CK => clk, RB => resetn, Q => out_buf_4_port);
   out_buf_reg_7_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => n245,
                           CK => clk, RB => resetn, Q => out_buf_3_port);
   out_buf_reg_7_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => n245,
                           CK => clk, RB => resetn, Q => out_buf_2_port);
   out_buf_reg_7_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => n245,
                           CK => clk, RB => resetn, Q => out_buf_1_port);
   out_buf_reg_7_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => n245,
                           CK => clk, RB => resetn, Q => out_buf_0_port);
   in_buf_reg_1_0_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n165, 
                           CK => clk, RB => resetn, Q => in_buf_192_port);
   out_buf_reg_3_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_143_port
                           );
   out_buf_reg_3_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_142_port
                           );
   out_buf_reg_3_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_141_port
                           );
   out_buf_reg_3_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_140_port
                           );
   out_buf_reg_3_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_139_port
                           );
   out_buf_reg_3_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_138_port
                           );
   out_buf_reg_3_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => n252,
                           CK => clk, RB => resetn, Q => out_buf_137_port);
   out_buf_reg_3_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => n252,
                           CK => clk, RB => resetn, Q => out_buf_136_port);
   out_buf_reg_3_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => n252,
                           CK => clk, RB => resetn, Q => out_buf_135_port);
   out_buf_reg_3_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => n252,
                           CK => clk, RB => resetn, Q => out_buf_134_port);
   out_buf_reg_3_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => n252,
                           CK => clk, RB => resetn, Q => out_buf_133_port);
   out_buf_reg_3_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => n252,
                           CK => clk, RB => resetn, Q => out_buf_132_port);
   out_buf_reg_3_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => n252,
                           CK => clk, RB => resetn, Q => out_buf_131_port);
   out_buf_reg_3_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => n252,
                           CK => clk, RB => resetn, Q => out_buf_130_port);
   out_buf_reg_3_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => n252,
                           CK => clk, RB => resetn, Q => out_buf_129_port);
   out_buf_reg_3_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => n252,
                           CK => clk, RB => resetn, Q => out_buf_128_port);
   in_buf_reg_0_0_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n163, 
                           CK => clk, RB => resetn, Q => in_buf_224_port);
   in_buf_reg_4_0_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n171, 
                           CK => clk, RB => resetn, Q => in_buf_96_port);
   out_buf_reg_2_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_175_port
                           );
   out_buf_reg_2_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_174_port
                           );
   out_buf_reg_2_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_173_port
                           );
   out_buf_reg_2_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_172_port
                           );
   out_buf_reg_2_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_171_port
                           );
   out_buf_reg_2_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_170_port
                           );
   out_buf_reg_2_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => n251,
                           CK => clk, RB => resetn, Q => out_buf_169_port);
   out_buf_reg_2_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => n251,
                           CK => clk, RB => resetn, Q => out_buf_168_port);
   out_buf_reg_2_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => n251,
                           CK => clk, RB => resetn, Q => out_buf_167_port);
   out_buf_reg_2_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => n251,
                           CK => clk, RB => resetn, Q => out_buf_166_port);
   out_buf_reg_2_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => n251,
                           CK => clk, RB => resetn, Q => out_buf_165_port);
   out_buf_reg_2_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => n251,
                           CK => clk, RB => resetn, Q => out_buf_164_port);
   out_buf_reg_2_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => n251,
                           CK => clk, RB => resetn, Q => out_buf_163_port);
   out_buf_reg_2_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => n251,
                           CK => clk, RB => resetn, Q => out_buf_162_port);
   out_buf_reg_2_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => n251,
                           CK => clk, RB => resetn, Q => out_buf_161_port);
   out_buf_reg_2_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => n251,
                           CK => clk, RB => resetn, Q => out_buf_160_port);
   out_buf_reg_6_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_47_port)
                           ;
   out_buf_reg_6_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_46_port)
                           ;
   out_buf_reg_6_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_45_port)
                           ;
   out_buf_reg_6_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_44_port)
                           ;
   out_buf_reg_6_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_43_port)
                           ;
   out_buf_reg_6_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_42_port)
                           ;
   out_buf_reg_6_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => n250,
                           CK => clk, RB => resetn, Q => out_buf_41_port);
   out_buf_reg_6_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => n250,
                           CK => clk, RB => resetn, Q => out_buf_40_port);
   out_buf_reg_6_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => n250,
                           CK => clk, RB => resetn, Q => out_buf_39_port);
   out_buf_reg_6_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => n250,
                           CK => clk, RB => resetn, Q => out_buf_38_port);
   out_buf_reg_6_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => n250,
                           CK => clk, RB => resetn, Q => out_buf_37_port);
   out_buf_reg_6_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => n250,
                           CK => clk, RB => resetn, Q => out_buf_36_port);
   out_buf_reg_6_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => n250,
                           CK => clk, RB => resetn, Q => out_buf_35_port);
   out_buf_reg_6_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => n250,
                           CK => clk, RB => resetn, Q => out_buf_34_port);
   out_buf_reg_6_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => n250,
                           CK => clk, RB => resetn, Q => out_buf_33_port);
   out_buf_reg_6_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => n250,
                           CK => clk, RB => resetn, Q => out_buf_32_port);
   out_buf_reg_7_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n245, CK => clk, RB => resetn, Q => out_buf_31_port)
                           ;
   out_buf_reg_7_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n245, CK => clk, RB => resetn, Q => out_buf_30_port)
                           ;
   out_buf_reg_7_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n245, CK => clk, RB => resetn, Q => out_buf_29_port)
                           ;
   out_buf_reg_7_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n245, CK => clk, RB => resetn, Q => out_buf_28_port)
                           ;
   out_buf_reg_7_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n245, CK => clk, RB => resetn, Q => out_buf_27_port)
                           ;
   out_buf_reg_7_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n245, CK => clk, RB => resetn, Q => out_buf_26_port)
                           ;
   out_buf_reg_7_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n245, CK => clk, RB => resetn, Q => out_buf_25_port)
                           ;
   out_buf_reg_7_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n245, CK => clk, RB => resetn, Q => out_buf_24_port)
                           ;
   out_buf_reg_7_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n245, CK => clk, RB => resetn, Q => out_buf_23_port)
                           ;
   out_buf_reg_7_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n245, CK => clk, RB => resetn, Q => out_buf_22_port)
                           ;
   out_buf_reg_7_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n245, CK => clk, RB => resetn, Q => out_buf_21_port)
                           ;
   out_buf_reg_7_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n245, CK => clk, RB => resetn, Q => out_buf_20_port)
                           ;
   out_buf_reg_7_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n245, CK => clk, RB => resetn, Q => out_buf_19_port)
                           ;
   out_buf_reg_7_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n245, CK => clk, RB => resetn, Q => out_buf_18_port)
                           ;
   out_buf_reg_7_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n245, CK => clk, RB => resetn, Q => out_buf_17_port)
                           ;
   out_buf_reg_7_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n245, CK => clk, RB => resetn, Q => out_buf_16_port)
                           ;
   out_buf_reg_5_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_79_port)
                           ;
   out_buf_reg_5_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_78_port)
                           ;
   out_buf_reg_5_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_77_port)
                           ;
   out_buf_reg_5_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_76_port)
                           ;
   out_buf_reg_5_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_75_port)
                           ;
   out_buf_reg_5_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_74_port)
                           ;
   out_buf_reg_5_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => n249,
                           CK => clk, RB => resetn, Q => out_buf_73_port);
   out_buf_reg_5_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => n249,
                           CK => clk, RB => resetn, Q => out_buf_72_port);
   out_buf_reg_5_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => n249,
                           CK => clk, RB => resetn, Q => out_buf_71_port);
   out_buf_reg_5_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => n249,
                           CK => clk, RB => resetn, Q => out_buf_70_port);
   out_buf_reg_5_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => n249,
                           CK => clk, RB => resetn, Q => out_buf_69_port);
   out_buf_reg_5_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => n249,
                           CK => clk, RB => resetn, Q => out_buf_68_port);
   out_buf_reg_5_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => n249,
                           CK => clk, RB => resetn, Q => out_buf_67_port);
   out_buf_reg_5_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => n249,
                           CK => clk, RB => resetn, Q => out_buf_66_port);
   out_buf_reg_5_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => n249,
                           CK => clk, RB => resetn, Q => out_buf_65_port);
   out_buf_reg_5_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => n249,
                           CK => clk, RB => resetn, Q => out_buf_64_port);
   out_buf_reg_3_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_159_port
                           );
   out_buf_reg_3_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_158_port
                           );
   out_buf_reg_3_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_157_port
                           );
   out_buf_reg_3_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_156_port
                           );
   out_buf_reg_3_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_155_port
                           );
   out_buf_reg_3_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_154_port
                           );
   out_buf_reg_3_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_153_port
                           );
   out_buf_reg_3_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_152_port
                           );
   out_buf_reg_3_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_151_port
                           );
   out_buf_reg_3_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_150_port
                           );
   out_buf_reg_3_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_149_port
                           );
   out_buf_reg_3_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_148_port
                           );
   out_buf_reg_3_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_147_port
                           );
   out_buf_reg_3_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_146_port
                           );
   out_buf_reg_3_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_145_port
                           );
   out_buf_reg_3_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_144_port
                           );
   out_buf_reg_1_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_207_port
                           );
   out_buf_reg_1_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_206_port
                           );
   out_buf_reg_1_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_205_port
                           );
   out_buf_reg_1_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_204_port
                           );
   out_buf_reg_1_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_203_port
                           );
   out_buf_reg_1_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_202_port
                           );
   out_buf_reg_1_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => n248,
                           CK => clk, RB => resetn, Q => out_buf_201_port);
   out_buf_reg_1_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => n248,
                           CK => clk, RB => resetn, Q => out_buf_200_port);
   out_buf_reg_1_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => n248,
                           CK => clk, RB => resetn, Q => out_buf_199_port);
   out_buf_reg_1_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => n248,
                           CK => clk, RB => resetn, Q => out_buf_198_port);
   out_buf_reg_1_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => n248,
                           CK => clk, RB => resetn, Q => out_buf_197_port);
   out_buf_reg_1_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => n248,
                           CK => clk, RB => resetn, Q => out_buf_196_port);
   out_buf_reg_1_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => n248,
                           CK => clk, RB => resetn, Q => out_buf_195_port);
   out_buf_reg_1_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => n248,
                           CK => clk, RB => resetn, Q => out_buf_194_port);
   out_buf_reg_1_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => n248,
                           CK => clk, RB => resetn, Q => out_buf_193_port);
   out_buf_reg_1_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => n248,
                           CK => clk, RB => resetn, Q => out_buf_192_port);
   out_buf_reg_2_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_191_port
                           );
   out_buf_reg_2_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_190_port
                           );
   out_buf_reg_2_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_189_port
                           );
   out_buf_reg_2_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_188_port
                           );
   out_buf_reg_2_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_187_port
                           );
   out_buf_reg_2_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_186_port
                           );
   out_buf_reg_2_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_185_port
                           );
   out_buf_reg_2_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_184_port
                           );
   out_buf_reg_2_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_183_port
                           );
   out_buf_reg_2_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_182_port
                           );
   out_buf_reg_2_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_181_port
                           );
   out_buf_reg_2_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_180_port
                           );
   out_buf_reg_2_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_179_port
                           );
   out_buf_reg_2_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_178_port
                           );
   out_buf_reg_2_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_177_port
                           );
   out_buf_reg_2_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_176_port
                           );
   out_buf_reg_6_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_63_port)
                           ;
   out_buf_reg_6_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_62_port)
                           ;
   out_buf_reg_6_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_61_port)
                           ;
   out_buf_reg_6_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_60_port)
                           ;
   out_buf_reg_6_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_59_port)
                           ;
   out_buf_reg_6_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_58_port)
                           ;
   out_buf_reg_6_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_57_port)
                           ;
   out_buf_reg_6_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_56_port)
                           ;
   out_buf_reg_6_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_55_port)
                           ;
   out_buf_reg_6_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_54_port)
                           ;
   out_buf_reg_6_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_53_port)
                           ;
   out_buf_reg_6_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_52_port)
                           ;
   out_buf_reg_6_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_51_port)
                           ;
   out_buf_reg_6_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_50_port)
                           ;
   out_buf_reg_6_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_49_port)
                           ;
   out_buf_reg_6_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_48_port)
                           ;
   out_buf_reg_0_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_239_port
                           );
   out_buf_reg_0_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_238_port
                           );
   out_buf_reg_0_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_237_port
                           );
   out_buf_reg_0_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_236_port
                           );
   out_buf_reg_0_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_235_port
                           );
   out_buf_reg_0_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_234_port
                           );
   out_buf_reg_0_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => n247,
                           CK => clk, RB => resetn, Q => out_buf_233_port);
   out_buf_reg_0_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => n247,
                           CK => clk, RB => resetn, Q => out_buf_232_port);
   out_buf_reg_0_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => n247,
                           CK => clk, RB => resetn, Q => out_buf_231_port);
   out_buf_reg_0_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => n247,
                           CK => clk, RB => resetn, Q => out_buf_230_port);
   out_buf_reg_0_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => n247,
                           CK => clk, RB => resetn, Q => out_buf_229_port);
   out_buf_reg_0_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => n247,
                           CK => clk, RB => resetn, Q => out_buf_228_port);
   out_buf_reg_0_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => n247,
                           CK => clk, RB => resetn, Q => out_buf_227_port);
   out_buf_reg_0_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => n247,
                           CK => clk, RB => resetn, Q => out_buf_226_port);
   out_buf_reg_0_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => n247,
                           CK => clk, RB => resetn, Q => out_buf_225_port);
   out_buf_reg_0_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => n247,
                           CK => clk, RB => resetn, Q => out_buf_224_port);
   out_buf_reg_4_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_111_port
                           );
   out_buf_reg_4_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_110_port
                           );
   out_buf_reg_4_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_109_port
                           );
   out_buf_reg_4_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_108_port
                           );
   out_buf_reg_4_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_107_port
                           );
   out_buf_reg_4_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_106_port
                           );
   out_buf_reg_4_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => n246,
                           CK => clk, RB => resetn, Q => out_buf_105_port);
   out_buf_reg_4_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => n246,
                           CK => clk, RB => resetn, Q => out_buf_104_port);
   out_buf_reg_4_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => n246,
                           CK => clk, RB => resetn, Q => out_buf_103_port);
   out_buf_reg_4_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => n246,
                           CK => clk, RB => resetn, Q => out_buf_102_port);
   out_buf_reg_4_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => n246,
                           CK => clk, RB => resetn, Q => out_buf_101_port);
   out_buf_reg_4_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => n246,
                           CK => clk, RB => resetn, Q => out_buf_100_port);
   out_buf_reg_4_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => n246,
                           CK => clk, RB => resetn, Q => out_buf_99_port);
   out_buf_reg_4_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => n246,
                           CK => clk, RB => resetn, Q => out_buf_98_port);
   out_buf_reg_4_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => n246,
                           CK => clk, RB => resetn, Q => out_buf_97_port);
   out_buf_reg_4_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => n246,
                           CK => clk, RB => resetn, Q => out_buf_96_port);
   out_buf_reg_5_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_95_port)
                           ;
   out_buf_reg_5_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_94_port)
                           ;
   out_buf_reg_5_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_93_port)
                           ;
   out_buf_reg_5_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_92_port)
                           ;
   out_buf_reg_5_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_91_port)
                           ;
   out_buf_reg_5_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_90_port)
                           ;
   out_buf_reg_5_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_89_port)
                           ;
   out_buf_reg_5_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_88_port)
                           ;
   out_buf_reg_5_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_87_port)
                           ;
   out_buf_reg_5_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_86_port)
                           ;
   out_buf_reg_5_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_85_port)
                           ;
   out_buf_reg_5_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_84_port)
                           ;
   out_buf_reg_5_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_83_port)
                           ;
   out_buf_reg_5_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_82_port)
                           ;
   out_buf_reg_5_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_81_port)
                           ;
   out_buf_reg_5_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_80_port)
                           ;
   out_buf_reg_1_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_223_port
                           );
   out_buf_reg_1_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_222_port
                           );
   out_buf_reg_1_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_221_port
                           );
   out_buf_reg_1_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_220_port
                           );
   out_buf_reg_1_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_219_port
                           );
   out_buf_reg_1_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_218_port
                           );
   out_buf_reg_1_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_217_port
                           );
   out_buf_reg_1_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_216_port
                           );
   out_buf_reg_1_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_215_port
                           );
   out_buf_reg_1_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_214_port
                           );
   out_buf_reg_1_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_213_port
                           );
   out_buf_reg_1_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_212_port
                           );
   out_buf_reg_1_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_211_port
                           );
   out_buf_reg_1_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_210_port
                           );
   out_buf_reg_1_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_209_port
                           );
   out_buf_reg_1_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_208_port
                           );
   out_buf_reg_0_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_255_port
                           );
   out_buf_reg_0_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_254_port
                           );
   out_buf_reg_0_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_253_port
                           );
   out_buf_reg_0_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_252_port
                           );
   out_buf_reg_0_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_251_port
                           );
   out_buf_reg_0_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_250_port
                           );
   out_buf_reg_0_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_249_port
                           );
   out_buf_reg_0_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_248_port
                           );
   out_buf_reg_0_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_247_port
                           );
   out_buf_reg_0_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_246_port
                           );
   out_buf_reg_0_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_245_port
                           );
   out_buf_reg_0_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_244_port
                           );
   out_buf_reg_0_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_243_port
                           );
   out_buf_reg_0_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_242_port
                           );
   out_buf_reg_0_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_241_port
                           );
   out_buf_reg_0_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_240_port
                           );
   out_buf_reg_4_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_127_port
                           );
   out_buf_reg_4_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_126_port
                           );
   out_buf_reg_4_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_125_port
                           );
   out_buf_reg_4_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_124_port
                           );
   out_buf_reg_4_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_123_port
                           );
   out_buf_reg_4_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_122_port
                           );
   out_buf_reg_4_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_121_port
                           );
   out_buf_reg_4_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_120_port
                           );
   out_buf_reg_4_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_119_port
                           );
   out_buf_reg_4_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_118_port
                           );
   out_buf_reg_4_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_117_port
                           );
   out_buf_reg_4_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_116_port
                           );
   out_buf_reg_4_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_115_port
                           );
   out_buf_reg_4_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_114_port
                           );
   out_buf_reg_4_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_113_port
                           );
   out_buf_reg_4_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_112_port
                           );
   out_trigger_reg : DFFRPQ1 port map( D => n240, CK => clk, RB => resetn, Q =>
                           out_trigger);
   read_comp_res_reg : DFERPQ1 port map( D => avs_writedata(2), CEB => n179, CK
                           => clk, RB => resetn, Q => read_comp_res);
   in_counter_reg_0_inst : DFERPQ1 port map( D => n155, CEB => n683, CK => clk,
                           RB => resetn, Q => in_counter_0_port);
   in_counter_reg_2_inst : DFFRPQ1 port map( D => n238, CK => clk, RB => resetn
                           , Q => in_counter_2_port);
   in_counter_reg_1_inst : DFFRPQ1 port map( D => n237, CK => clk, RB => resetn
                           , Q => in_counter_1_port);
   in_busy_reg : DFFRPQ1 port map( D => n239, CK => clk, RB => resetn, Q => 
                           in_busy);
   odd_reg : DFFRPQ1 port map( D => n156, CK => clk, RB => resetn, Q => odd);
   out_busy_reg : DFFRPQ1 port map( D => n234, CK => clk, RB => resetn, Q => 
                           out_busy);
   odd_reg2 : DFFRPQ1 port map( D => n154, CK => clk, RB => resetn, Q => odd1);
   operand_load_reg : DFERPQ1 port map( D => avs_writedata(1), CEB => n179, CK 
                           => clk, RB => resetn, Q => operand_load);
   coeff_load_reg : DFERPQ1 port map( D => avs_writedata(0), CEB => n179, CK =>
                           clk, RB => resetn, Q => coeff_load);
   out_counter_reg_0_inst : DFFRPQ1 port map( D => n236, CK => clk, RB => 
                           resetn, Q => N62);
   out_counter_reg_2_inst : DFFRPQ1 port map( D => n235, CK => clk, RB => 
                           resetn, Q => N64);
   out_counter_reg_1_inst : DFFRPQ1 port map( D => n201, CK => clk, RB => 
                           resetn, Q => N63);
   operand_regs_reg_3_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_159_port);
   operand_regs_reg_5_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_95_port);
   operand_regs_reg_1_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_223_port);
   coeff_memory_reg_1_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_31_port);
   coeff_memory_reg_2_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB 
                           => n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_31_port);
   coeff_memory_reg_3_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_31_port);
   coeff_memory_reg_0_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_31_port);
   coeff_memory_reg_4_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_31_port);
   operand_regs_reg_2_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB 
                           => n254, CK => clk, RB => resetn, Q => 
                           operand_regs_191_port);
   operand_regs_reg_4_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_127_port);
   operand_regs_reg_6_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_63_port);
   operand_regs_reg_7_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB 
                           => n253, CK => clk, RB => resetn, Q => 
                           operand_regs_31_port);
   operand_regs_reg_3_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_158_port);
   operand_regs_reg_5_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_94_port);
   operand_regs_reg_0_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_255_port);
   operand_regs_reg_3_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_157_port);
   operand_regs_reg_5_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_93_port);
   coeff_memory_reg_1_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_30_port);
   coeff_memory_reg_2_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB 
                           => n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_30_port);
   coeff_memory_reg_3_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_30_port);
   coeff_memory_reg_0_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_30_port);
   coeff_memory_reg_4_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_30_port);
   operand_regs_reg_2_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB 
                           => n254, CK => clk, RB => resetn, Q => 
                           operand_regs_190_port);
   operand_regs_reg_4_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_126_port);
   operand_regs_reg_6_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_62_port);
   operand_regs_reg_1_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_222_port);
   operand_regs_reg_7_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB 
                           => n253, CK => clk, RB => resetn, Q => 
                           operand_regs_30_port);
   operand_regs_reg_0_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_254_port);
   operand_regs_reg_1_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_221_port);
   operand_regs_reg_3_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_156_port);
   operand_regs_reg_5_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_92_port);
   operand_regs_reg_1_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_220_port);
   coeff_memory_reg_1_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_29_port);
   coeff_memory_reg_2_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB 
                           => n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_29_port);
   coeff_memory_reg_3_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_29_port);
   operand_regs_reg_3_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_155_port);
   operand_regs_reg_5_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_91_port);
   coeff_memory_reg_0_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_29_port);
   coeff_memory_reg_4_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_29_port);
   operand_regs_reg_2_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB 
                           => n254, CK => clk, RB => resetn, Q => 
                           operand_regs_189_port);
   operand_regs_reg_4_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_125_port);
   operand_regs_reg_6_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_61_port);
   operand_regs_reg_7_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB 
                           => n253, CK => clk, RB => resetn, Q => 
                           operand_regs_29_port);
   operand_regs_reg_0_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_253_port);
   coeff_memory_reg_1_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_28_port);
   coeff_memory_reg_2_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB 
                           => n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_28_port);
   coeff_memory_reg_3_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_28_port);
   coeff_memory_reg_0_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_28_port);
   coeff_memory_reg_4_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_28_port);
   operand_regs_reg_2_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB 
                           => n254, CK => clk, RB => resetn, Q => 
                           operand_regs_188_port);
   operand_regs_reg_4_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_124_port);
   operand_regs_reg_6_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_60_port);
   operand_regs_reg_7_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB 
                           => n253, CK => clk, RB => resetn, Q => 
                           operand_regs_28_port);
   operand_regs_reg_0_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_252_port);
   operand_regs_reg_1_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_219_port);
   coeff_memory_reg_1_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_27_port);
   coeff_memory_reg_2_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB 
                           => n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_27_port);
   coeff_memory_reg_3_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_27_port);
   operand_regs_reg_3_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_154_port);
   operand_regs_reg_5_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_90_port);
   coeff_memory_reg_0_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_27_port);
   coeff_memory_reg_4_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_27_port);
   operand_regs_reg_2_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB 
                           => n254, CK => clk, RB => resetn, Q => 
                           operand_regs_187_port);
   operand_regs_reg_4_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_123_port);
   operand_regs_reg_6_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_59_port);
   operand_regs_reg_7_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB 
                           => n253, CK => clk, RB => resetn, Q => 
                           operand_regs_27_port);
   operand_regs_reg_0_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_251_port);
   coeff_memory_reg_1_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_26_port);
   coeff_memory_reg_2_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB 
                           => n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_26_port);
   coeff_memory_reg_3_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_26_port);
   coeff_memory_reg_0_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_26_port);
   coeff_memory_reg_4_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_26_port);
   operand_regs_reg_2_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB 
                           => n254, CK => clk, RB => resetn, Q => 
                           operand_regs_186_port);
   operand_regs_reg_4_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_122_port);
   operand_regs_reg_6_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_58_port);
   operand_regs_reg_7_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB 
                           => n253, CK => clk, RB => resetn, Q => 
                           operand_regs_26_port);
   operand_regs_reg_1_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_218_port);
   operand_regs_reg_0_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_250_port);
   operand_regs_reg_3_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_153_port);
   operand_regs_reg_5_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_89_port);
   operand_regs_reg_1_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_217_port);
   coeff_memory_reg_1_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_25_port);
   coeff_memory_reg_2_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB 
                           => n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_25_port);
   coeff_memory_reg_3_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_25_port);
   coeff_memory_reg_0_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_25_port);
   coeff_memory_reg_4_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_25_port);
   operand_regs_reg_2_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB 
                           => n254, CK => clk, RB => resetn, Q => 
                           operand_regs_185_port);
   operand_regs_reg_4_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_121_port);
   operand_regs_reg_6_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_57_port);
   operand_regs_reg_7_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB 
                           => n253, CK => clk, RB => resetn, Q => 
                           operand_regs_25_port);
   operand_regs_reg_0_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_249_port);
   operand_regs_reg_3_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_152_port);
   operand_regs_reg_5_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_88_port);
   coeff_memory_reg_1_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_24_port);
   coeff_memory_reg_2_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB 
                           => n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_24_port);
   coeff_memory_reg_3_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_24_port);
   coeff_memory_reg_0_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_24_port);
   coeff_memory_reg_4_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_24_port);
   operand_regs_reg_2_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB 
                           => n254, CK => clk, RB => resetn, Q => 
                           operand_regs_184_port);
   operand_regs_reg_4_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_120_port);
   operand_regs_reg_6_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_56_port);
   operand_regs_reg_0_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_248_port);
   operand_regs_reg_7_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB 
                           => n253, CK => clk, RB => resetn, Q => 
                           operand_regs_24_port);
   operand_regs_reg_1_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_216_port);
   operand_regs_reg_3_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_151_port);
   operand_regs_reg_5_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_87_port);
   operand_regs_reg_1_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_215_port);
   coeff_memory_reg_1_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_23_port);
   coeff_memory_reg_2_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB 
                           => n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_23_port);
   coeff_memory_reg_3_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_23_port);
   coeff_memory_reg_0_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_23_port);
   coeff_memory_reg_4_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_23_port);
   operand_regs_reg_2_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB 
                           => n254, CK => clk, RB => resetn, Q => 
                           operand_regs_183_port);
   operand_regs_reg_4_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_119_port);
   operand_regs_reg_6_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_55_port);
   operand_regs_reg_7_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB 
                           => n253, CK => clk, RB => resetn, Q => 
                           operand_regs_23_port);
   operand_regs_reg_0_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_247_port);
   operand_regs_reg_3_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_150_port);
   operand_regs_reg_5_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_86_port);
   operand_regs_reg_3_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_149_port);
   operand_regs_reg_5_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_85_port);
   coeff_memory_reg_1_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_22_port);
   coeff_memory_reg_2_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB 
                           => n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_22_port);
   coeff_memory_reg_3_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_22_port);
   coeff_memory_reg_0_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_22_port);
   coeff_memory_reg_4_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_22_port);
   operand_regs_reg_2_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB 
                           => n254, CK => clk, RB => resetn, Q => 
                           operand_regs_182_port);
   operand_regs_reg_4_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_118_port);
   operand_regs_reg_6_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_54_port);
   operand_regs_reg_0_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_246_port);
   operand_regs_reg_7_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB 
                           => n253, CK => clk, RB => resetn, Q => 
                           operand_regs_22_port);
   operand_regs_reg_1_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_214_port);
   operand_regs_reg_1_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_213_port);
   coeff_memory_reg_1_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_21_port);
   coeff_memory_reg_2_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB 
                           => n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_21_port);
   coeff_memory_reg_3_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_21_port);
   operand_regs_reg_3_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_148_port);
   operand_regs_reg_5_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_84_port);
   operand_regs_reg_3_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_147_port);
   operand_regs_reg_5_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_83_port);
   coeff_memory_reg_0_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_21_port);
   coeff_memory_reg_4_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_21_port);
   operand_regs_reg_2_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB 
                           => n254, CK => clk, RB => resetn, Q => 
                           operand_regs_181_port);
   operand_regs_reg_4_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_117_port);
   operand_regs_reg_6_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_53_port);
   operand_regs_reg_7_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB 
                           => n253, CK => clk, RB => resetn, Q => 
                           operand_regs_21_port);
   operand_regs_reg_0_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_245_port);
   coeff_memory_reg_1_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_20_port);
   coeff_memory_reg_2_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB 
                           => n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_20_port);
   coeff_memory_reg_3_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_20_port);
   coeff_memory_reg_0_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_20_port);
   coeff_memory_reg_4_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_20_port);
   operand_regs_reg_2_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB 
                           => n254, CK => clk, RB => resetn, Q => 
                           operand_regs_180_port);
   operand_regs_reg_4_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_116_port);
   operand_regs_reg_6_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_52_port);
   operand_regs_reg_0_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_244_port);
   operand_regs_reg_7_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB 
                           => n253, CK => clk, RB => resetn, Q => 
                           operand_regs_20_port);
   operand_regs_reg_1_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_212_port);
   operand_regs_reg_1_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_211_port);
   operand_regs_reg_5_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_82_port);
   operand_regs_reg_3_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_146_port);
   operand_regs_reg_3_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_145_port);
   operand_regs_reg_5_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_81_port);
   operand_regs_reg_1_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_210_port);
   coeff_memory_reg_1_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_19_port);
   coeff_memory_reg_2_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB 
                           => n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_19_port);
   coeff_memory_reg_3_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_19_port);
   coeff_memory_reg_0_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_19_port);
   coeff_memory_reg_4_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_19_port);
   operand_regs_reg_2_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB 
                           => n254, CK => clk, RB => resetn, Q => 
                           operand_regs_179_port);
   operand_regs_reg_4_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_115_port);
   operand_regs_reg_6_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_51_port);
   operand_regs_reg_7_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB 
                           => n253, CK => clk, RB => resetn, Q => 
                           operand_regs_19_port);
   operand_regs_reg_0_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_243_port);
   operand_regs_reg_1_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_209_port);
   coeff_memory_reg_1_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_18_port);
   coeff_memory_reg_2_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB 
                           => n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_18_port);
   coeff_memory_reg_3_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_18_port);
   coeff_memory_reg_0_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_18_port);
   coeff_memory_reg_4_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_18_port);
   operand_regs_reg_2_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB 
                           => n254, CK => clk, RB => resetn, Q => 
                           operand_regs_178_port);
   operand_regs_reg_4_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_114_port);
   operand_regs_reg_6_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_50_port);
   operand_regs_reg_7_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB 
                           => n253, CK => clk, RB => resetn, Q => 
                           operand_regs_18_port);
   operand_regs_reg_0_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_242_port);
   operand_regs_reg_3_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_144_port);
   operand_regs_reg_5_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_80_port);
   coeff_memory_reg_1_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_17_port);
   coeff_memory_reg_2_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB 
                           => n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_17_port);
   coeff_memory_reg_3_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_17_port);
   coeff_memory_reg_0_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_17_port);
   coeff_memory_reg_4_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_17_port);
   operand_regs_reg_2_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB 
                           => n254, CK => clk, RB => resetn, Q => 
                           operand_regs_177_port);
   operand_regs_reg_4_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_113_port);
   operand_regs_reg_6_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_49_port);
   operand_regs_reg_7_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB 
                           => n253, CK => clk, RB => resetn, Q => 
                           operand_regs_17_port);
   operand_regs_reg_0_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_241_port);
   coeff_memory_reg_1_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_16_port);
   coeff_memory_reg_2_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB 
                           => n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_16_port);
   coeff_memory_reg_3_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_16_port);
   coeff_memory_reg_0_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_16_port);
   coeff_memory_reg_4_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_16_port);
   operand_regs_reg_2_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB 
                           => n254, CK => clk, RB => resetn, Q => 
                           operand_regs_176_port);
   operand_regs_reg_4_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_112_port);
   operand_regs_reg_6_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_48_port);
   operand_regs_reg_7_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB 
                           => n253, CK => clk, RB => resetn, Q => 
                           operand_regs_16_port);
   operand_regs_reg_0_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_240_port);
   operand_regs_reg_1_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_208_port);
   operand_regs_reg_3_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_143_port);
   operand_regs_reg_5_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_79_port);
   coeff_memory_reg_1_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_15_port);
   coeff_memory_reg_2_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB 
                           => n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_15_port);
   coeff_memory_reg_3_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_15_port);
   coeff_memory_reg_0_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_15_port);
   coeff_memory_reg_4_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_15_port);
   operand_regs_reg_2_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB 
                           => n254, CK => clk, RB => resetn, Q => 
                           operand_regs_175_port);
   operand_regs_reg_4_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_111_port);
   operand_regs_reg_6_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_47_port);
   operand_regs_reg_0_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_239_port);
   operand_regs_reg_3_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_142_port);
   operand_regs_reg_5_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_78_port);
   operand_regs_reg_7_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB 
                           => n253, CK => clk, RB => resetn, Q => 
                           operand_regs_15_port);
   operand_regs_reg_3_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_141_port);
   operand_regs_reg_5_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_77_port);
   operand_regs_reg_1_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_207_port);
   coeff_memory_reg_1_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_14_port);
   coeff_memory_reg_2_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB 
                           => n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_14_port);
   coeff_memory_reg_3_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_14_port);
   coeff_memory_reg_0_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_14_port);
   coeff_memory_reg_4_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_14_port);
   operand_regs_reg_2_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB 
                           => n254, CK => clk, RB => resetn, Q => 
                           operand_regs_174_port);
   operand_regs_reg_4_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_110_port);
   operand_regs_reg_6_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_46_port);
   operand_regs_reg_0_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_238_port);
   operand_regs_reg_7_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB 
                           => n253, CK => clk, RB => resetn, Q => 
                           operand_regs_14_port);
   operand_regs_reg_1_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_206_port);
   operand_regs_reg_1_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_205_port);
   coeff_memory_reg_1_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_13_port);
   coeff_memory_reg_2_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB 
                           => n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_13_port);
   coeff_memory_reg_3_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_13_port);
   coeff_memory_reg_0_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_13_port);
   coeff_memory_reg_4_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_13_port);
   operand_regs_reg_2_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB 
                           => n254, CK => clk, RB => resetn, Q => 
                           operand_regs_173_port);
   operand_regs_reg_4_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_109_port);
   operand_regs_reg_6_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_45_port);
   operand_regs_reg_7_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB 
                           => n253, CK => clk, RB => resetn, Q => 
                           operand_regs_13_port);
   operand_regs_reg_0_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_237_port);
   operand_regs_reg_3_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_140_port);
   operand_regs_reg_5_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_76_port);
   operand_regs_reg_3_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_139_port);
   operand_regs_reg_5_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_75_port);
   coeff_memory_reg_1_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_12_port);
   coeff_memory_reg_2_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB 
                           => n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_12_port);
   coeff_memory_reg_3_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_12_port);
   coeff_memory_reg_0_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_12_port);
   coeff_memory_reg_4_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_12_port);
   operand_regs_reg_2_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB 
                           => n254, CK => clk, RB => resetn, Q => 
                           operand_regs_172_port);
   operand_regs_reg_4_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_108_port);
   operand_regs_reg_6_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_44_port);
   operand_regs_reg_0_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_236_port);
   operand_regs_reg_3_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_138_port);
   operand_regs_reg_5_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_74_port);
   operand_regs_reg_7_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB 
                           => n253, CK => clk, RB => resetn, Q => 
                           operand_regs_12_port);
   operand_regs_reg_1_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_203_port);
   operand_regs_reg_1_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_204_port);
   coeff_memory_reg_1_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_11_port);
   coeff_memory_reg_2_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB 
                           => n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_11_port);
   coeff_memory_reg_3_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_11_port);
   coeff_memory_reg_0_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_11_port);
   coeff_memory_reg_4_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_11_port);
   operand_regs_reg_2_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB 
                           => n254, CK => clk, RB => resetn, Q => 
                           operand_regs_171_port);
   operand_regs_reg_4_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_107_port);
   operand_regs_reg_6_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_43_port);
   operand_regs_reg_7_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB 
                           => n253, CK => clk, RB => resetn, Q => 
                           operand_regs_11_port);
   operand_regs_reg_0_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_235_port);
   operand_regs_reg_3_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_137_port);
   operand_regs_reg_5_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_73_port);
   coeff_memory_reg_1_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_10_port);
   coeff_memory_reg_2_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB 
                           => n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_10_port);
   coeff_memory_reg_3_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_10_port);
   coeff_memory_reg_0_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_10_port);
   coeff_memory_reg_4_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_10_port);
   operand_regs_reg_2_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB 
                           => n254, CK => clk, RB => resetn, Q => 
                           operand_regs_170_port);
   operand_regs_reg_4_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_106_port);
   operand_regs_reg_6_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_42_port);
   operand_regs_reg_7_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB 
                           => n253, CK => clk, RB => resetn, Q => 
                           operand_regs_10_port);
   operand_regs_reg_1_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_202_port);
   operand_regs_reg_0_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_234_port);
   coeff_memory_reg_1_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_9_port);
   coeff_memory_reg_2_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_9_port);
   coeff_memory_reg_3_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_9_port);
   operand_regs_reg_1_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_201_port);
   coeff_memory_reg_0_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_9_port);
   coeff_memory_reg_4_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_9_port);
   operand_regs_reg_2_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_169_port);
   operand_regs_reg_4_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_105_port);
   operand_regs_reg_6_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_41_port);
   operand_regs_reg_7_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_9_port);
   operand_regs_reg_0_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_233_port);
   operand_regs_reg_3_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_135_port);
   operand_regs_reg_5_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_71_port);
   operand_regs_reg_3_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_136_port);
   operand_regs_reg_5_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_72_port);
   coeff_memory_reg_1_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_8_port);
   coeff_memory_reg_2_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_8_port);
   coeff_memory_reg_3_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_8_port);
   coeff_memory_reg_0_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_8_port);
   coeff_memory_reg_4_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_8_port);
   operand_regs_reg_2_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_168_port);
   operand_regs_reg_4_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_104_port);
   operand_regs_reg_6_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_40_port);
   operand_regs_reg_0_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_232_port);
   operand_regs_reg_7_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_8_port);
   operand_regs_reg_3_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_134_port);
   operand_regs_reg_5_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_70_port);
   operand_regs_reg_1_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_199_port);
   operand_regs_reg_1_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_200_port);
   operand_regs_reg_1_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_198_port);
   coeff_memory_reg_1_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_7_port);
   coeff_memory_reg_2_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_7_port);
   coeff_memory_reg_3_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_7_port);
   operand_regs_reg_3_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_133_port);
   operand_regs_reg_5_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_69_port);
   coeff_memory_reg_0_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_7_port);
   coeff_memory_reg_4_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_7_port);
   operand_regs_reg_2_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_167_port);
   operand_regs_reg_4_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_103_port);
   operand_regs_reg_6_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_39_port);
   operand_regs_reg_7_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_7_port);
   operand_regs_reg_0_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_231_port);
   operand_regs_reg_1_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_197_port);
   coeff_memory_reg_1_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_6_port);
   coeff_memory_reg_2_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_6_port);
   coeff_memory_reg_3_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_6_port);
   coeff_memory_reg_0_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_6_port);
   coeff_memory_reg_4_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_6_port);
   operand_regs_reg_2_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_166_port);
   operand_regs_reg_4_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_102_port);
   operand_regs_reg_6_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_38_port);
   operand_regs_reg_7_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_6_port);
   operand_regs_reg_0_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_230_port);
   coeff_memory_reg_1_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_5_port);
   coeff_memory_reg_2_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_5_port);
   coeff_memory_reg_3_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_5_port);
   coeff_memory_reg_0_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_5_port);
   coeff_memory_reg_4_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_5_port);
   operand_regs_reg_2_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_165_port);
   operand_regs_reg_4_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_101_port);
   operand_regs_reg_6_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_37_port);
   operand_regs_reg_7_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_5_port);
   operand_regs_reg_0_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_229_port);
   operand_regs_reg_3_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_132_port);
   operand_regs_reg_5_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_68_port);
   operand_regs_reg_3_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_131_port);
   operand_regs_reg_5_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_67_port);
   coeff_memory_reg_1_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_4_port);
   coeff_memory_reg_2_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_4_port);
   coeff_memory_reg_3_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_4_port);
   coeff_memory_reg_0_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_4_port);
   coeff_memory_reg_4_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_4_port);
   operand_regs_reg_2_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_164_port);
   operand_regs_reg_4_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_100_port);
   operand_regs_reg_6_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_36_port);
   operand_regs_reg_7_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_4_port);
   operand_regs_reg_0_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_228_port);
   operand_regs_reg_1_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_196_port);
   operand_regs_reg_1_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_195_port);
   coeff_memory_reg_1_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_3_port);
   coeff_memory_reg_2_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_3_port);
   coeff_memory_reg_3_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_3_port);
   coeff_memory_reg_0_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_3_port);
   coeff_memory_reg_4_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_3_port);
   operand_regs_reg_2_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_163_port);
   operand_regs_reg_4_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_99_port);
   operand_regs_reg_6_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_35_port);
   operand_regs_reg_7_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_3_port);
   operand_regs_reg_3_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_128_port);
   operand_regs_reg_5_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_64_port);
   operand_regs_reg_0_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_227_port);
   coeff_memory_reg_1_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_2_port);
   coeff_memory_reg_2_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_2_port);
   coeff_memory_reg_3_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_2_port);
   coeff_memory_reg_0_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_2_port);
   coeff_memory_reg_4_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_2_port);
   operand_regs_reg_2_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_162_port);
   operand_regs_reg_4_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_98_port);
   operand_regs_reg_6_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_34_port);
   operand_regs_reg_3_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_129_port);
   operand_regs_reg_5_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_65_port);
   operand_regs_reg_3_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_130_port);
   operand_regs_reg_5_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_66_port);
   operand_regs_reg_1_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_192_port);
   operand_regs_reg_0_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_226_port);
   operand_regs_reg_7_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_2_port);
   operand_regs_reg_1_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_193_port);
   operand_regs_reg_1_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_194_port);
   coeff_memory_reg_1_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_1_port);
   coeff_memory_reg_2_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_1_port);
   coeff_memory_reg_3_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_1_port);
   coeff_memory_reg_0_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_1_port);
   coeff_memory_reg_4_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_1_port);
   operand_regs_reg_2_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_161_port);
   operand_regs_reg_4_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_97_port);
   operand_regs_reg_6_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_33_port);
   operand_regs_reg_7_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_1_port);
   operand_regs_reg_0_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_225_port);
   coeff_memory_reg_1_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_0_port);
   coeff_memory_reg_2_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_0_port);
   coeff_memory_reg_3_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_0_port);
   coeff_memory_reg_0_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_0_port);
   coeff_memory_reg_4_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_0_port);
   operand_regs_reg_2_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_160_port);
   operand_regs_reg_4_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_96_port);
   operand_regs_reg_6_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_32_port);
   operand_regs_reg_7_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_0_port);
   operand_regs_reg_0_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_224_port);
   filt_mult_inputs_reg : DFERPQ1 port map( D => avs_writedata(0), CEB => n178,
                           CK => clk, RB => resetn, Q => filt_mult_inputs);
   avs_readdata_reg_30_inst : DFFSPQ1 port map( D => n203, CK => clk, SB => 
                           resetn, Q => avs_readdata_30_port);
   avs_readdata_reg_28_inst : DFFSPQ1 port map( D => n205, CK => clk, SB => 
                           resetn, Q => avs_readdata_28_port);
   avs_readdata_reg_26_inst : DFFSPQ1 port map( D => n207, CK => clk, SB => 
                           resetn, Q => avs_readdata_26_port);
   avs_readdata_reg_24_inst : DFFSPQ1 port map( D => n209, CK => clk, SB => 
                           resetn, Q => avs_readdata_24_port);
   avs_readdata_reg_22_inst : DFFSPQ1 port map( D => n211, CK => clk, SB => 
                           resetn, Q => avs_readdata_22_port);
   avs_readdata_reg_20_inst : DFFSPQ1 port map( D => n213, CK => clk, SB => 
                           resetn, Q => avs_readdata_20_port);
   avs_readdata_reg_18_inst : DFFSPQ1 port map( D => n215, CK => clk, SB => 
                           resetn, Q => avs_readdata_18_port);
   avs_readdata_reg_16_inst : DFFSPQ1 port map( D => n217, CK => clk, SB => 
                           resetn, Q => avs_readdata_16_port);
   avs_readdata_reg_14_inst : DFFSPQ1 port map( D => n219, CK => clk, SB => 
                           resetn, Q => avs_readdata_14_port);
   avs_readdata_reg_12_inst : DFFSPQ1 port map( D => n221, CK => clk, SB => 
                           resetn, Q => avs_readdata_12_port);
   avs_readdata_reg_10_inst : DFFSPQ1 port map( D => n223, CK => clk, SB => 
                           resetn, Q => avs_readdata_10_port);
   avs_readdata_reg_8_inst : DFFSPQ1 port map( D => n225, CK => clk, SB => 
                           resetn, Q => avs_readdata_8_port);
   avs_readdata_reg_6_inst : DFFSPQ1 port map( D => n227, CK => clk, SB => 
                           resetn, Q => avs_readdata_6_port);
   avs_readdata_reg_4_inst : DFFSPQ1 port map( D => n229, CK => clk, SB => 
                           resetn, Q => avs_readdata_4_port);
   avs_readdata_reg_2_inst : DFFSPQ1 port map( D => n231, CK => clk, SB => 
                           resetn, Q => avs_readdata_2_port);
   avs_readdata_reg_0_inst : DFFSPQ1 port map( D => n233, CK => clk, SB => 
                           resetn, Q => avs_readdata_0_port);
   avs_readdata_reg_31_inst : DFFRPQ1 port map( D => n202, CK => clk, RB => 
                           resetn, Q => avs_readdata_31_port);
   avs_readdata_reg_29_inst : DFFRPQ1 port map( D => n204, CK => clk, RB => 
                           resetn, Q => avs_readdata_29_port);
   avs_readdata_reg_27_inst : DFFRPQ1 port map( D => n206, CK => clk, RB => 
                           resetn, Q => avs_readdata_27_port);
   avs_readdata_reg_25_inst : DFFRPQ1 port map( D => n208, CK => clk, RB => 
                           resetn, Q => avs_readdata_25_port);
   avs_readdata_reg_23_inst : DFFRPQ1 port map( D => n210, CK => clk, RB => 
                           resetn, Q => avs_readdata_23_port);
   avs_readdata_reg_21_inst : DFFRPQ1 port map( D => n212, CK => clk, RB => 
                           resetn, Q => avs_readdata_21_port);
   avs_readdata_reg_19_inst : DFFRPQ1 port map( D => n214, CK => clk, RB => 
                           resetn, Q => avs_readdata_19_port);
   avs_readdata_reg_17_inst : DFFRPQ1 port map( D => n216, CK => clk, RB => 
                           resetn, Q => avs_readdata_17_port);
   avs_readdata_reg_15_inst : DFFRPQ1 port map( D => n218, CK => clk, RB => 
                           resetn, Q => avs_readdata_15_port);
   avs_readdata_reg_13_inst : DFFRPQ1 port map( D => n220, CK => clk, RB => 
                           resetn, Q => avs_readdata_13_port);
   avs_readdata_reg_11_inst : DFFRPQ1 port map( D => n222, CK => clk, RB => 
                           resetn, Q => avs_readdata_11_port);
   avs_readdata_reg_9_inst : DFFRPQ1 port map( D => n224, CK => clk, RB => 
                           resetn, Q => avs_readdata_9_port);
   avs_readdata_reg_7_inst : DFFRPQ1 port map( D => n226, CK => clk, RB => 
                           resetn, Q => avs_readdata_7_port);
   avs_readdata_reg_5_inst : DFFRPQ1 port map( D => n228, CK => clk, RB => 
                           resetn, Q => avs_readdata_5_port);
   avs_readdata_reg_3_inst : DFFRPQ1 port map( D => n230, CK => clk, RB => 
                           resetn, Q => avs_readdata_3_port);
   avs_readdata_reg_1_inst : DFFRPQ1 port map( D => n232, CK => clk, RB => 
                           resetn, Q => avs_readdata_1_port);
   stop_sim_reg : DFFRPQ1 port map( D => n157, CK => clk, RB => resetn, Q => 
                           stop_sim_port);
   siso_req_reg : DFERPQ1 port map( D => n690, CEB => n161, CK => clk, RB => 
                           resetn, Q => siso_req);
   siso_data_out_reg_0_inst : DFERPQ1 port map( D => N2888, CEB => n695, CK => 
                           clk, RB => resetn, Q => siso_data_out(0));
   siso_data_out_reg_15_inst : DFERPQ1 port map( D => N2903, CEB => n695, CK =>
                           clk, RB => resetn, Q => siso_data_out(15));
   siso_data_out_reg_14_inst : DFERPQ1 port map( D => N2902, CEB => n695, CK =>
                           clk, RB => resetn, Q => siso_data_out(14));
   siso_data_out_reg_13_inst : DFERPQ1 port map( D => N2901, CEB => n695, CK =>
                           clk, RB => resetn, Q => siso_data_out(13));
   siso_data_out_reg_12_inst : DFERPQ1 port map( D => N2900, CEB => n695, CK =>
                           clk, RB => resetn, Q => siso_data_out(12));
   siso_data_out_reg_11_inst : DFERPQ1 port map( D => N2899, CEB => n695, CK =>
                           clk, RB => resetn, Q => siso_data_out(11));
   siso_data_out_reg_10_inst : DFERPQ1 port map( D => N2898, CEB => n695, CK =>
                           clk, RB => resetn, Q => siso_data_out(10));
   siso_data_out_reg_9_inst : DFERPQ1 port map( D => N2897, CEB => n695, CK => 
                           clk, RB => resetn, Q => siso_data_out(9));
   siso_data_out_reg_8_inst : DFERPQ1 port map( D => N2896, CEB => n695, CK => 
                           clk, RB => resetn, Q => siso_data_out(8));
   siso_data_out_reg_7_inst : DFERPQ1 port map( D => N2895, CEB => n695, CK => 
                           clk, RB => resetn, Q => siso_data_out(7));
   siso_data_out_reg_6_inst : DFERPQ1 port map( D => N2894, CEB => n695, CK => 
                           clk, RB => resetn, Q => siso_data_out(6));
   siso_data_out_reg_5_inst : DFERPQ1 port map( D => N2893, CEB => n695, CK => 
                           clk, RB => resetn, Q => siso_data_out(5));
   siso_data_out_reg_4_inst : DFERPQ1 port map( D => N2892, CEB => n695, CK => 
                           clk, RB => resetn, Q => siso_data_out(4));
   siso_data_out_reg_3_inst : DFERPQ1 port map( D => N2891, CEB => n695, CK => 
                           clk, RB => resetn, Q => siso_data_out(3));
   siso_data_out_reg_2_inst : DFERPQ1 port map( D => N2890, CEB => n695, CK => 
                           clk, RB => resetn, Q => siso_data_out(2));
   siso_data_out_reg_1_inst : DFERPQ1 port map( D => N2889, CEB => n695, CK => 
                           clk, RB => resetn, Q => siso_data_out(1));
   siso_ready_reg : DFFRPQ1 port map( D => out_busy, CK => clk, RB => resetn, Q
                           => siso_ready);
   U642 : AND2D1 port map( A1 => n289, A2 => avs_addr(0), Z => n242);
   U643 : AND2D1 port map( A1 => n536, A2 => N62, Z => n243);
   U644 : AND2D1 port map( A1 => n538, A2 => N62, Z => n244);
   U645 : NAN3D1 port map( A1 => n106, A2 => avs_addr(0), A3 => n110, Z => n245
                           );
   U646 : NAN2D1 port map( A1 => n110, A2 => n99, Z => n246);
   U647 : NAN2D1 port map( A1 => n110, A2 => n97, Z => n247);
   U648 : NAN2D1 port map( A1 => n110, A2 => n93, Z => n248);
   U649 : NAN2D1 port map( A1 => n110, A2 => n109, Z => n249);
   U650 : NAN2D1 port map( A1 => n110, A2 => n108, Z => n250);
   U651 : NAN2D1 port map( A1 => n110, A2 => n69, Z => n251);
   U652 : NAN2D1 port map( A1 => n110, A2 => n68, Z => n252);
   U653 : NAN3D1 port map( A1 => n106, A2 => avs_addr(0), A3 => n107, Z => n253
                           );
   U654 : NAN2D1 port map( A1 => n107, A2 => n69, Z => n254);
   U655 : NAN2D1 port map( A1 => n107, A2 => n68, Z => n255);
   U656 : NAN2D1 port map( A1 => n107, A2 => n97, Z => n256);
   U657 : NAN2D1 port map( A1 => n107, A2 => n93, Z => n257);
   U658 : NAN2D1 port map( A1 => n107, A2 => n99, Z => n258);
   U659 : NAN2D1 port map( A1 => n108, A2 => n107, Z => n259);
   U660 : NAN2D1 port map( A1 => n109, A2 => n107, Z => n260);
   U661 : NAN2D1 port map( A1 => n103, A2 => n68, Z => n261);
   U662 : NAN2D1 port map( A1 => n103, A2 => n69, Z => n262);
   U663 : NAN2D1 port map( A1 => n103, A2 => n97, Z => n263);
   U664 : NAN2D1 port map( A1 => n103, A2 => n93, Z => n264);
   U665 : NAN2D1 port map( A1 => n103, A2 => n99, Z => n265);
   U666 : AND2D1 port map( A1 => n288, A2 => avs_addr(0), Z => n266);
   U667 : AND3D1 port map( A1 => N66, A2 => n270, A3 => read_comp_res, Z => 
                           n267);
   U668 : AND2D1 port map( A1 => n535, A2 => N62, Z => n268);
   U669 : AND2D1 port map( A1 => n537, A2 => N62, Z => n269);
   U670 : BUFBD2 port map( A => filt_mult_inputs, Z => n673);
   U671 : INVD1 port map( A => n528, Z => n529);
   U672 : INVD1 port map( A => n533, Z => n534);
   U673 : INVD1 port map( A => n530, Z => n532);
   U674 : INVD1 port map( A => n530, Z => n531);
   U675 : INVD1 port map( A => n526, Z => n527);
   U676 : INVD1 port map( A => n523, Z => n524);
   U677 : INVD1 port map( A => n523, Z => n525);
   U678 : INVD1 port map( A => n74, Z => n677);
   U679 : INVD1 port map( A => n96, Z => n678);
   U680 : NAN2D1 port map( A1 => n118, A2 => n691, Z => n176);
   U681 : NAN2D1 port map( A1 => n689, A2 => n118, Z => n174);
   U682 : NOR2M1D1 port map( A1 => n104, A2 => n686, Z => n103);
   U683 : INVD1 port map( A => n270, Z => n676);
   U684 : INVD1 port map( A => n516, Z => n528);
   U685 : INVD1 port map( A => n518, Z => n533);
   U686 : INVD1 port map( A => n517, Z => n530);
   U687 : INVD1 port map( A => n675, Z => n674);
   U688 : INVD1 port map( A => n513, Z => n523);
   U689 : INVD1 port map( A => n514, Z => n526);
   U690 : NAN2D1 port map( A1 => n93, A2 => n679, Z => n74);
   U691 : OAI211D1 port map( A1 => n6300, A2 => n6400, B => n270, C => n65, Z 
                           => n14);
   U692 : NOR2D1 port map( A1 => n68, A2 => n69, Z => n6300);
   U693 : NOR3D1 port map( A1 => n677, A2 => N66, A3 => n678, Z => n65);
   U694 : AND2D1 port map( A1 => n111, A2 => n681, Z => n99);
   U695 : INVD1 port map( A => n6400, Z => n679);
   U696 : NAN2D1 port map( A1 => n97, A2 => n679, Z => n96);
   U697 : AND2D1 port map( A1 => n106, A2 => n681, Z => n108);
   U698 : INVD1 port map( A => n673, Z => n276);
   U699 : INVD1 port map( A => n673, Z => n278);
   U700 : INVD1 port map( A => n673, Z => n279);
   U701 : INVD1 port map( A => n673, Z => n275);
   U702 : INVD1 port map( A => n673, Z => n281);
   U703 : INVD1 port map( A => n673, Z => n272);
   U704 : INVD1 port map( A => n673, Z => n285);
   U705 : INVD1 port map( A => n673, Z => n284);
   U706 : INVD1 port map( A => n673, Z => n280);
   U707 : INVD1 port map( A => n673, Z => n286);
   U708 : INVD1 port map( A => n673, Z => n271);
   U709 : INVD1 port map( A => n673, Z => n273);
   U710 : INVD1 port map( A => n673, Z => n274);
   U711 : INVD1 port map( A => n673, Z => n282);
   U712 : INVD1 port map( A => n673, Z => n277);
   U713 : INVD1 port map( A => n673, Z => n283);
   U714 : INVD1 port map( A => n673, Z => n287);
   U715 : NOR3D1 port map( A1 => n697, A2 => n694, A3 => n671, Z => n78);
   U716 : INVD1 port map( A => n81, Z => n684);
   U717 : INVD1 port map( A => n672, Z => n696);
   U718 : NOR2D1 port map( A1 => n693, A2 => n687, Z => n118);
   U719 : INVD1 port map( A => n88, Z => n691);
   U720 : NOR2D1 port map( A1 => n683, A2 => n91, Z => n89);
   U721 : INVD1 port map( A => n84, Z => n683);
   U722 : INVD1 port map( A => n155, Z => n688);
   U723 : NAN2D1 port map( A1 => n119, A2 => n115, Z => n171);
   U724 : NAN2D1 port map( A1 => n119, A2 => n101, Z => n162);
   U725 : NAN2D1 port map( A1 => n119, A2 => n118, Z => n170);
   U726 : NAN2D1 port map( A1 => n120, A2 => n119, Z => n163);
   U727 : NAN2D1 port map( A1 => n87, A2 => n84, Z => n86);
   U728 : NAN2D1 port map( A1 => n689, A2 => n115, Z => n175);
   U729 : NAN2D1 port map( A1 => n120, A2 => n689, Z => n167);
   U730 : NAN2D1 port map( A1 => n689, A2 => n101, Z => n166);
   U731 : INVD1 port map( A => n85, Z => n689);
   U732 : NAN2D1 port map( A1 => n87, A2 => n101, Z => n164);
   U733 : NAN2D1 port map( A1 => n115, A2 => n87, Z => n173);
   U734 : NAN2D1 port map( A1 => n120, A2 => n87, Z => n165);
   U735 : NAN2D1 port map( A1 => n118, A2 => n87, Z => n172);
   U736 : NAN2D1 port map( A1 => n691, A2 => n101, Z => n168);
   U737 : NAN2D1 port map( A1 => n115, A2 => n691, Z => n177);
   U738 : NAN2D1 port map( A1 => n120, A2 => n691, Z => n169);
   U739 : NOR3M1D1 port map( A1 => n104, A2 => coeff_load, A3 => operand_load, 
                           Z => n110);
   U740 : AND2D1 port map( A1 => N66, A2 => avs_write, Z => n104);
   U741 : AND3D1 port map( A1 => n686, A2 => n104, A3 => operand_load, Z => 
                           n107);
   U742 : NAN4D1 port map( A1 => n5900, A2 => n14, A3 => n6000, A4 => n6100, Z 
                           => n233);
   U743 : NAN2M1D1 port map( A1 => n70, A2 => n270, Z => n5900);
   U744 : NAN2D1 port map( A1 => N2009, A2 => n267, Z => n6000);
   U745 : INVD1 port map( A => n12, Z => n675);
   U746 : NOR3M1D1 port map( A1 => N66, A2 => n676, A3 => read_comp_res, Z => 
                           n12);
   U747 : INVD1 port map( A => avs_write, Z => n682);
   U748 : AND2D1 port map( A1 => avs_read, A2 => n682, Z => n270);
   U749 : NAN3D1 port map( A1 => n56, A2 => n14, A3 => n57, Z => n231);
   U750 : NAN2D1 port map( A1 => N2007, A2 => n267, Z => n56);
   U751 : NAN3D1 port map( A1 => n427, A2 => n426, A3 => n428, Z => N2007);
   U752 : NAN3D1 port map( A1 => n53, A2 => n14, A3 => n54, Z => n229);
   U753 : NAN2D1 port map( A1 => N2005, A2 => n267, Z => n53);
   U754 : NAN3D1 port map( A1 => n433, A2 => n432, A3 => n434, Z => N2005);
   U755 : NAN3D1 port map( A1 => n50, A2 => n14, A3 => n51, Z => n227);
   U756 : NAN2D1 port map( A1 => N2003, A2 => n267, Z => n50);
   U757 : NAN3D1 port map( A1 => n439, A2 => n438, A3 => n440, Z => N2003);
   U758 : NAN3D1 port map( A1 => n47, A2 => n14, A3 => n48, Z => n225);
   U759 : NAN2D1 port map( A1 => N2001, A2 => n267, Z => n47);
   U760 : NAN3D1 port map( A1 => n445, A2 => n444, A3 => n446, Z => N2001);
   U761 : NAN3D1 port map( A1 => n44, A2 => n14, A3 => n45, Z => n223);
   U762 : NAN2D1 port map( A1 => N1999, A2 => n267, Z => n44);
   U763 : NAN3D1 port map( A1 => n451, A2 => n450, A3 => n452, Z => N1999);
   U764 : NAN3D1 port map( A1 => n41, A2 => n14, A3 => n42, Z => n221);
   U765 : NAN2D1 port map( A1 => N1997, A2 => n267, Z => n41);
   U766 : NAN3D1 port map( A1 => n457, A2 => n456, A3 => n458, Z => N1997);
   U767 : NAN3D1 port map( A1 => n38, A2 => n14, A3 => n39, Z => n219);
   U768 : NAN2D1 port map( A1 => N1995, A2 => n267, Z => n38);
   U769 : NAN3D1 port map( A1 => n463, A2 => n462, A3 => n464, Z => N1995);
   U770 : NAN3D1 port map( A1 => n35, A2 => n14, A3 => n36, Z => n217);
   U771 : NAN2D1 port map( A1 => N1993, A2 => n267, Z => n35);
   U772 : NAN3D1 port map( A1 => n469, A2 => n468, A3 => n470, Z => N1993);
   U773 : NAN3D1 port map( A1 => n13, A2 => n14, A3 => n15, Z => n203);
   U774 : NAN2D1 port map( A1 => N1979, A2 => n267, Z => n13);
   U775 : NAN3D1 port map( A1 => n511, A2 => n510, A3 => n512, Z => N1979);
   U776 : INVD1 port map( A => avs_addr(2), Z => n522);
   U777 : NAN3D1 port map( A1 => n32, A2 => n14, A3 => n33, Z => n215);
   U778 : NAN2D1 port map( A1 => N1991, A2 => n267, Z => n32);
   U779 : NAN3D1 port map( A1 => n475, A2 => n474, A3 => n476, Z => N1991);
   U780 : NAN3D1 port map( A1 => n29, A2 => n14, A3 => n30, Z => n213);
   U781 : NAN2D1 port map( A1 => N1989, A2 => n267, Z => n29);
   U782 : NAN3D1 port map( A1 => n481, A2 => n480, A3 => n482, Z => N1989);
   U783 : NAN3D1 port map( A1 => n26, A2 => n14, A3 => n27, Z => n211);
   U784 : NAN2D1 port map( A1 => N1987, A2 => n267, Z => n26);
   U785 : NAN3D1 port map( A1 => n487, A2 => n486, A3 => n488, Z => N1987);
   U786 : NAN3D1 port map( A1 => n23, A2 => n14, A3 => n24, Z => n209);
   U787 : NAN2D1 port map( A1 => N1985, A2 => n267, Z => n23);
   U788 : NAN3D1 port map( A1 => n493, A2 => n492, A3 => n494, Z => N1985);
   U789 : NAN3D1 port map( A1 => n20, A2 => n14, A3 => n21, Z => n207);
   U790 : NAN2D1 port map( A1 => N1983, A2 => n267, Z => n20);
   U791 : NAN3D1 port map( A1 => n499, A2 => n498, A3 => n500, Z => N1983);
   U792 : NAN3D1 port map( A1 => n17, A2 => n14, A3 => n18, Z => n205);
   U793 : NAN2D1 port map( A1 => N1981, A2 => n267, Z => n17);
   U794 : NAN3D1 port map( A1 => n505, A2 => n504, A3 => n506, Z => N1981);
   U795 : OAI21M20D1 port map( A1 => avs_readdata_1_port, A2 => n676, B => n58,
                           Z => n232);
   U796 : NAN3D1 port map( A1 => n424, A2 => n423, A3 => n425, Z => N2008);
   U797 : OAI21M20D1 port map( A1 => avs_readdata_3_port, A2 => n676, B => n55,
                           Z => n230);
   U798 : NAN3D1 port map( A1 => n430, A2 => n429, A3 => n431, Z => N2006);
   U799 : OAI21M20D1 port map( A1 => avs_readdata_5_port, A2 => n676, B => n52,
                           Z => n228);
   U800 : NAN3D1 port map( A1 => n436, A2 => n435, A3 => n437, Z => N2004);
   U801 : OAI21M20D1 port map( A1 => avs_readdata_7_port, A2 => n676, B => n49,
                           Z => n226);
   U802 : NAN3D1 port map( A1 => n442, A2 => n441, A3 => n443, Z => N2002);
   U803 : OAI21M20D1 port map( A1 => avs_readdata_15_port, A2 => n676, B => n37
                           , Z => n218);
   U804 : NAN3D1 port map( A1 => n466, A2 => n465, A3 => n467, Z => N1994);
   U805 : OAI21M20D1 port map( A1 => avs_readdata_17_port, A2 => n676, B => n34
                           , Z => n216);
   U806 : NAN3D1 port map( A1 => n472, A2 => n471, A3 => n473, Z => N1992);
   U807 : OAI21M20D1 port map( A1 => avs_readdata_19_port, A2 => n676, B => n31
                           , Z => n214);
   U808 : NAN3D1 port map( A1 => n478, A2 => n477, A3 => n479, Z => N1990);
   U809 : OAI21M20D1 port map( A1 => avs_readdata_21_port, A2 => n676, B => n28
                           , Z => n212);
   U810 : NAN3D1 port map( A1 => n484, A2 => n483, A3 => n485, Z => N1988);
   U811 : OAI21M20D1 port map( A1 => avs_readdata_23_port, A2 => n676, B => n25
                           , Z => n210);
   U812 : NAN3D1 port map( A1 => n490, A2 => n489, A3 => n491, Z => N1986);
   U813 : OAI21M20D1 port map( A1 => avs_readdata_25_port, A2 => n676, B => n22
                           , Z => n208);
   U814 : NAN3D1 port map( A1 => n496, A2 => n495, A3 => n497, Z => N1984);
   U815 : OAI21M20D1 port map( A1 => avs_readdata_27_port, A2 => n676, B => n19
                           , Z => n206);
   U816 : NAN3D1 port map( A1 => n502, A2 => n501, A3 => n503, Z => N1982);
   U817 : OAI21M20D1 port map( A1 => avs_readdata_29_port, A2 => n676, B => n16
                           , Z => n204);
   U818 : NAN3D1 port map( A1 => n508, A2 => n507, A3 => n509, Z => N1980);
   U819 : OAI21M20D1 port map( A1 => avs_readdata_31_port, A2 => n676, B => n10
                           , Z => n202);
   U820 : OAI21M20D1 port map( A1 => avs_readdata_9_port, A2 => n676, B => n46,
                           Z => n224);
   U821 : NAN3D1 port map( A1 => n448, A2 => n447, A3 => n449, Z => N2000);
   U822 : OAI21M20D1 port map( A1 => avs_readdata_11_port, A2 => n676, B => n43
                           , Z => n222);
   U823 : NAN3D1 port map( A1 => n454, A2 => n453, A3 => n455, Z => N1998);
   U824 : OAI21M20D1 port map( A1 => avs_readdata_13_port, A2 => n676, B => n40
                           , Z => n220);
   U825 : NAN3D1 port map( A1 => n460, A2 => n459, A3 => n461, Z => N1996);
   U826 : NAN3D1 port map( A1 => n520, A2 => n519, A3 => n521, Z => N1978);
   U827 : NAN2D1 port map( A1 => comp_res_31_port, A2 => n529, Z => n520);
   U828 : AOI22M10D1 port map( B1 => in_buf_63_port, B2 => n515, A1 => n528, A2
                           => in_buf_127_port, Z => n417);
   U829 : NAN3D1 port map( A1 => n421, A2 => n420, A3 => n422, Z => N2009);
   U830 : NAN2D1 port map( A1 => comp_res_0_port, A2 => n529, Z => n421);
   U831 : NAN2D1 port map( A1 => comp_res_25_port, A2 => n529, Z => n496);
   U832 : NAN2D1 port map( A1 => comp_res_27_port, A2 => n529, Z => n502);
   U833 : NAN2D1 port map( A1 => comp_res_29_port, A2 => n529, Z => n508);
   U834 : NAN2D1 port map( A1 => comp_res_1_port, A2 => n529, Z => n424);
   U835 : NAN2D1 port map( A1 => comp_res_3_port, A2 => n529, Z => n430);
   U836 : NAN2D1 port map( A1 => comp_res_5_port, A2 => n529, Z => n436);
   U837 : NAN2D1 port map( A1 => comp_res_7_port, A2 => n529, Z => n442);
   U838 : NAN2D1 port map( A1 => comp_res_9_port, A2 => n529, Z => n448);
   U839 : NAN2D1 port map( A1 => comp_res_11_port, A2 => n529, Z => n454);
   U840 : NAN2D1 port map( A1 => comp_res_13_port, A2 => n529, Z => n460);
   U841 : NAN2D1 port map( A1 => comp_res_15_port, A2 => n529, Z => n466);
   U842 : NAN2D1 port map( A1 => comp_res_17_port, A2 => n516, Z => n472);
   U843 : NAN2D1 port map( A1 => comp_res_19_port, A2 => n529, Z => n478);
   U844 : NAN2D1 port map( A1 => comp_res_21_port, A2 => n516, Z => n484);
   U845 : NAN2D1 port map( A1 => comp_res_23_port, A2 => n516, Z => n490);
   U846 : NAN2D1 port map( A1 => comp_res_24_port, A2 => n529, Z => n493);
   U847 : NAN2D1 port map( A1 => comp_res_26_port, A2 => n529, Z => n499);
   U848 : NAN2D1 port map( A1 => comp_res_28_port, A2 => n529, Z => n505);
   U849 : NAN2D1 port map( A1 => comp_res_30_port, A2 => n529, Z => n511);
   U850 : NAN2D1 port map( A1 => comp_res_2_port, A2 => n516, Z => n427);
   U851 : NAN2D1 port map( A1 => comp_res_4_port, A2 => n516, Z => n433);
   U852 : NAN2D1 port map( A1 => comp_res_6_port, A2 => n516, Z => n439);
   U853 : NAN2D1 port map( A1 => comp_res_8_port, A2 => n516, Z => n445);
   U854 : NAN2D1 port map( A1 => comp_res_10_port, A2 => n516, Z => n451);
   U855 : NAN2D1 port map( A1 => comp_res_12_port, A2 => n516, Z => n457);
   U856 : NAN2D1 port map( A1 => comp_res_14_port, A2 => n516, Z => n463);
   U857 : NAN2D1 port map( A1 => comp_res_16_port, A2 => n516, Z => n469);
   U858 : NAN2D1 port map( A1 => comp_res_18_port, A2 => n516, Z => n475);
   U859 : NAN2D1 port map( A1 => comp_res_20_port, A2 => n516, Z => n481);
   U860 : NAN2D1 port map( A1 => comp_res_22_port, A2 => n516, Z => n487);
   U861 : NOR3D1 port map( A1 => avs_addr(1), A2 => avs_addr(2), A3 => n681, Z 
                           => n93);
   U862 : INVD1 port map( A => avs_addr(0), Z => n681);
   U863 : NOR3D1 port map( A1 => n681, A2 => avs_addr(2), A3 => n680, Z => n68)
                           ;
   U864 : INVD1 port map( A => avs_addr(1), Z => n680);
   U865 : NOR3D1 port map( A1 => avs_addr(0), A2 => avs_addr(2), A3 => n680, Z 
                           => n69);
   U866 : AND2D1 port map( A1 => avs_addr(2), A2 => n680, Z => n111);
   U867 : AND2D1 port map( A1 => n111, A2 => avs_addr(0), Z => n109);
   U868 : NAN2D1 port map( A1 => n114, A2 => avs_addr(3), Z => n6400);
   U869 : NOR2D1 port map( A1 => avs_addr(5), A2 => avs_addr(4), Z => n114);
   U870 : AND2D1 port map( A1 => avs_addr(2), A2 => avs_addr(1), Z => n106);
   U871 : NOR3D1 port map( A1 => avs_addr(1), A2 => avs_addr(2), A3 => 
                           avs_addr(0), Z => n97);
   U872 : NOR2D1 port map( A1 => n92, A2 => n682, Z => n240);
   U873 : NOR2D1 port map( A1 => n95, A2 => n682, Z => n241);
   U874 : NAN3D1 port map( A1 => avs_write, A2 => n679, A3 => n109, Z => n179);
   U875 : AO31D1 port map( A1 => avs_write, A2 => n679, A3 => n99, B => 
                           stop_sim_port, Z => n157);
   U876 : NAN3D1 port map( A1 => avs_write, A2 => n679, A3 => n108, Z => n178);
   U877 : AO22D1 port map( A1 => operand_regs_32_port, A2 => n278, B1 => 
                           coeff_memory_3_0_port, B2 => n673, Z => N3009);
   U878 : AO22D1 port map( A1 => operand_regs_96_port, A2 => n279, B1 => 
                           coeff_memory_2_0_port, B2 => n673, Z => N2977);
   U879 : AO22D1 port map( A1 => operand_regs_160_port, A2 => n276, B1 => 
                           coeff_memory_1_0_port, B2 => n673, Z => N2945);
   U880 : AO22D1 port map( A1 => coeff_memory_4_0_port, A2 => n673, B1 => n275,
                           B2 => operand_regs_0_port, Z => N3041);
   U881 : AO22D1 port map( A1 => coeff_memory_0_0_port, A2 => n673, B1 => n275,
                           B2 => operand_regs_224_port, Z => N2913);
   U882 : AO22D1 port map( A1 => operand_regs_33_port, A2 => n276, B1 => 
                           coeff_memory_3_1_port, B2 => n673, Z => N3010);
   U883 : AO22D1 port map( A1 => operand_regs_97_port, A2 => n278, B1 => 
                           coeff_memory_2_1_port, B2 => n673, Z => N2978);
   U884 : AO22D1 port map( A1 => operand_regs_161_port, A2 => n281, B1 => 
                           coeff_memory_1_1_port, B2 => n673, Z => N2946);
   U885 : AO22D1 port map( A1 => coeff_memory_4_1_port, A2 => n673, B1 => n275,
                           B2 => operand_regs_1_port, Z => N3042);
   U886 : AO22D1 port map( A1 => coeff_memory_0_1_port, A2 => n673, B1 => n272,
                           B2 => operand_regs_225_port, Z => N2914);
   U887 : AO22D1 port map( A1 => n673, A2 => operand_regs_194_port, B1 => n272,
                           B2 => operand_regs_2_port, Z => N3203);
   U888 : AO22D1 port map( A1 => n673, A2 => operand_regs_193_port, B1 => n272,
                           B2 => operand_regs_1_port, Z => N3202);
   U889 : OAI21M20D1 port map( A1 => operand_regs_66_port, A2 => n285, B => 
                           n151, Z => N3139);
   U890 : OAI21M20D1 port map( A1 => operand_regs_130_port, A2 => n285, B => 
                           n151, Z => N3107);
   U891 : OAI21M20D1 port map( A1 => operand_regs_65_port, A2 => n285, B => 
                           n152, Z => N3138);
   U892 : OAI21M20D1 port map( A1 => operand_regs_129_port, A2 => n284, B => 
                           n152, Z => N3106);
   U893 : AO22D1 port map( A1 => operand_regs_34_port, A2 => n278, B1 => 
                           coeff_memory_3_2_port, B2 => n673, Z => N3011);
   U894 : AO22D1 port map( A1 => operand_regs_98_port, A2 => n280, B1 => 
                           coeff_memory_2_2_port, B2 => n673, Z => N2979);
   U895 : AO22D1 port map( A1 => operand_regs_162_port, A2 => n281, B1 => 
                           coeff_memory_1_2_port, B2 => n673, Z => N2947);
   U896 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_194_port, B => 
                           n151, Z => N3075);
   U897 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_193_port, B => 
                           n152, Z => N3074);
   U898 : AO22D1 port map( A1 => n673, A2 => operand_regs_192_port, B1 => n271,
                           B2 => operand_regs_0_port, Z => N3201);
   U899 : AO22D1 port map( A1 => coeff_memory_4_2_port, A2 => n673, B1 => n275,
                           B2 => operand_regs_2_port, Z => N3043);
   U900 : AO22D1 port map( A1 => coeff_memory_0_2_port, A2 => n673, B1 => n271,
                           B2 => operand_regs_226_port, Z => N2915);
   U901 : OAI21M20D1 port map( A1 => operand_regs_64_port, A2 => n285, B => 
                           n153, Z => N3137);
   U902 : OAI21M20D1 port map( A1 => operand_regs_128_port, A2 => n284, B => 
                           n153, Z => N3105);
   U903 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_192_port, B => 
                           n153, Z => N3073);
   U904 : AO22D1 port map( A1 => operand_regs_35_port, A2 => n276, B1 => 
                           coeff_memory_3_3_port, B2 => n673, Z => N3012);
   U905 : AO22D1 port map( A1 => operand_regs_99_port, A2 => n280, B1 => 
                           coeff_memory_2_3_port, B2 => n673, Z => N2980);
   U906 : AO22D1 port map( A1 => operand_regs_163_port, A2 => n281, B1 => 
                           coeff_memory_1_3_port, B2 => n673, Z => N2948);
   U907 : AO22D1 port map( A1 => coeff_memory_4_3_port, A2 => n673, B1 => n275,
                           B2 => operand_regs_3_port, Z => N3044);
   U908 : AO22D1 port map( A1 => coeff_memory_0_3_port, A2 => n673, B1 => n272,
                           B2 => operand_regs_227_port, Z => N2916);
   U909 : AO22D1 port map( A1 => operand_regs_36_port, A2 => n278, B1 => 
                           coeff_memory_3_4_port, B2 => n673, Z => N3013);
   U910 : AO22D1 port map( A1 => operand_regs_100_port, A2 => n280, B1 => 
                           coeff_memory_2_4_port, B2 => n673, Z => N2981);
   U911 : AO22D1 port map( A1 => operand_regs_164_port, A2 => n281, B1 => 
                           coeff_memory_1_4_port, B2 => n673, Z => N2949);
   U912 : AO22D1 port map( A1 => n673, A2 => operand_regs_195_port, B1 => n273,
                           B2 => operand_regs_3_port, Z => N3204);
   U913 : AO22D1 port map( A1 => coeff_memory_4_4_port, A2 => n673, B1 => n275,
                           B2 => operand_regs_4_port, Z => N3045);
   U914 : AO22D1 port map( A1 => coeff_memory_0_4_port, A2 => n673, B1 => n272,
                           B2 => operand_regs_228_port, Z => N2917);
   U915 : AO22D1 port map( A1 => n673, A2 => operand_regs_196_port, B1 => n272,
                           B2 => operand_regs_4_port, Z => N3205);
   U916 : NAN2D1 port map( A1 => operand_regs_226_port, A2 => n673, Z => n151);
   U917 : NAN2D1 port map( A1 => operand_regs_225_port, A2 => n673, Z => n152);
   U918 : OAI21M20D1 port map( A1 => operand_regs_67_port, A2 => n285, B => 
                           n150, Z => N3140);
   U919 : OAI21M20D1 port map( A1 => operand_regs_131_port, A2 => n285, B => 
                           n150, Z => N3108);
   U920 : OAI21M20D1 port map( A1 => operand_regs_68_port, A2 => n285, B => 
                           n149, Z => N3141);
   U921 : OAI21M20D1 port map( A1 => operand_regs_132_port, A2 => n285, B => 
                           n149, Z => N3109);
   U922 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_195_port, B => 
                           n150, Z => N3076);
   U923 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_196_port, B => 
                           n149, Z => N3077);
   U924 : AO22D1 port map( A1 => operand_regs_37_port, A2 => n276, B1 => 
                           coeff_memory_3_5_port, B2 => n673, Z => N3014);
   U925 : AO22D1 port map( A1 => operand_regs_101_port, A2 => n280, B1 => 
                           coeff_memory_2_5_port, B2 => n673, Z => N2982);
   U926 : AO22D1 port map( A1 => operand_regs_165_port, A2 => n281, B1 => 
                           coeff_memory_1_5_port, B2 => n673, Z => N2950);
   U927 : NAN2D1 port map( A1 => operand_regs_224_port, A2 => n673, Z => n153);
   U928 : AO22D1 port map( A1 => coeff_memory_4_5_port, A2 => n673, B1 => n274,
                           B2 => operand_regs_5_port, Z => N3046);
   U929 : AO22D1 port map( A1 => coeff_memory_0_5_port, A2 => n673, B1 => n272,
                           B2 => operand_regs_229_port, Z => N2918);
   U930 : AO22D1 port map( A1 => operand_regs_38_port, A2 => n278, B1 => 
                           coeff_memory_3_6_port, B2 => n673, Z => N3015);
   U931 : AO22D1 port map( A1 => operand_regs_102_port, A2 => n280, B1 => 
                           coeff_memory_2_6_port, B2 => n673, Z => N2983);
   U932 : AO22D1 port map( A1 => operand_regs_166_port, A2 => n281, B1 => 
                           coeff_memory_1_6_port, B2 => n673, Z => N2951);
   U933 : AO22D1 port map( A1 => coeff_memory_4_6_port, A2 => n673, B1 => n274,
                           B2 => operand_regs_6_port, Z => N3047);
   U934 : AO22D1 port map( A1 => coeff_memory_0_6_port, A2 => n673, B1 => n272,
                           B2 => operand_regs_230_port, Z => N2919);
   U935 : NAN2D1 port map( A1 => operand_regs_227_port, A2 => n673, Z => n150);
   U936 : NAN2D1 port map( A1 => operand_regs_228_port, A2 => n673, Z => n149);
   U937 : AO22D1 port map( A1 => n673, A2 => operand_regs_197_port, B1 => n271,
                           B2 => operand_regs_5_port, Z => N3206);
   U938 : AO22D1 port map( A1 => operand_regs_39_port, A2 => n277, B1 => 
                           coeff_memory_3_7_port, B2 => n673, Z => N3016);
   U939 : AO22D1 port map( A1 => operand_regs_103_port, A2 => n280, B1 => 
                           coeff_memory_2_7_port, B2 => n673, Z => N2984);
   U940 : AO22D1 port map( A1 => operand_regs_167_port, A2 => n282, B1 => 
                           coeff_memory_1_7_port, B2 => n673, Z => N2952);
   U941 : OAI21M20D1 port map( A1 => operand_regs_69_port, A2 => n285, B => 
                           n148, Z => N3142);
   U942 : OAI21M20D1 port map( A1 => operand_regs_133_port, A2 => n284, B => 
                           n148, Z => N3110);
   U943 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_197_port, B => 
                           n148, Z => N3078);
   U944 : AO22D1 port map( A1 => coeff_memory_4_7_port, A2 => n673, B1 => n274,
                           B2 => operand_regs_7_port, Z => N3048);
   U945 : AO22D1 port map( A1 => coeff_memory_0_7_port, A2 => n673, B1 => n272,
                           B2 => operand_regs_231_port, Z => N2920);
   U946 : AO22D1 port map( A1 => n673, A2 => operand_regs_198_port, B1 => n272,
                           B2 => operand_regs_6_port, Z => N3207);
   U947 : OAI21M20D1 port map( A1 => operand_regs_134_port, A2 => n283, B => 
                           n147, Z => N3111);
   U948 : OAI21M20D1 port map( A1 => operand_regs_70_port, A2 => n285, B => 
                           n147, Z => N3143);
   U949 : NAN2D1 port map( A1 => operand_regs_229_port, A2 => n673, Z => n148);
   U950 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_198_port, B => 
                           n147, Z => N3079);
   U951 : AO22D1 port map( A1 => n673, A2 => operand_regs_200_port, B1 => n271,
                           B2 => operand_regs_8_port, Z => N3209);
   U952 : AO22D1 port map( A1 => n673, A2 => operand_regs_199_port, B1 => n273,
                           B2 => operand_regs_7_port, Z => N3208);
   U953 : AO22D1 port map( A1 => operand_regs_40_port, A2 => n278, B1 => 
                           coeff_memory_3_8_port, B2 => n673, Z => N3017);
   U954 : AO22D1 port map( A1 => operand_regs_104_port, A2 => n280, B1 => 
                           coeff_memory_2_8_port, B2 => n673, Z => N2985);
   U955 : AO22D1 port map( A1 => operand_regs_168_port, A2 => n282, B1 => 
                           coeff_memory_1_8_port, B2 => n673, Z => N2953);
   U956 : AO22D1 port map( A1 => coeff_memory_4_8_port, A2 => n673, B1 => n274,
                           B2 => operand_regs_8_port, Z => N3049);
   U957 : AO22D1 port map( A1 => coeff_memory_0_8_port, A2 => n673, B1 => n273,
                           B2 => operand_regs_232_port, Z => N2921);
   U958 : OAI21M20D1 port map( A1 => operand_regs_136_port, A2 => n283, B => 
                           n145, Z => N3113);
   U959 : OAI21M20D1 port map( A1 => operand_regs_72_port, A2 => n285, B => 
                           n145, Z => N3145);
   U960 : OAI21M20D1 port map( A1 => operand_regs_71_port, A2 => n285, B => 
                           n146, Z => N3144);
   U961 : OAI21M20D1 port map( A1 => operand_regs_135_port, A2 => n284, B => 
                           n146, Z => N3112);
   U962 : OAI21M20D1 port map( A1 => n283, A2 => operand_regs_199_port, B => 
                           n146, Z => N3080);
   U963 : OAI21M20D1 port map( A1 => n287, A2 => operand_regs_200_port, B => 
                           n145, Z => N3081);
   U964 : NAN2D1 port map( A1 => operand_regs_230_port, A2 => n673, Z => n147);
   U965 : AO22D1 port map( A1 => operand_regs_41_port, A2 => n276, B1 => 
                           coeff_memory_3_9_port, B2 => n673, Z => N3018);
   U966 : AO22D1 port map( A1 => operand_regs_105_port, A2 => n280, B1 => 
                           coeff_memory_2_9_port, B2 => n673, Z => N2986);
   U967 : AO22D1 port map( A1 => operand_regs_169_port, A2 => n282, B1 => 
                           coeff_memory_1_9_port, B2 => n673, Z => N2954);
   U968 : AO22D1 port map( A1 => coeff_memory_4_9_port, A2 => n673, B1 => n274,
                           B2 => operand_regs_9_port, Z => N3050);
   U969 : AO22D1 port map( A1 => coeff_memory_0_9_port, A2 => n673, B1 => n273,
                           B2 => operand_regs_233_port, Z => N2922);
   U970 : NAN2D1 port map( A1 => operand_regs_232_port, A2 => n673, Z => n145);
   U971 : NAN2D1 port map( A1 => operand_regs_231_port, A2 => n673, Z => n146);
   U972 : AO22D1 port map( A1 => n673, A2 => operand_regs_201_port, B1 => n271,
                           B2 => operand_regs_9_port, Z => N3210);
   U973 : AO22D1 port map( A1 => operand_regs_42_port, A2 => n277, B1 => 
                           coeff_memory_3_10_port, B2 => n673, Z => N3019);
   U974 : AO22D1 port map( A1 => operand_regs_106_port, A2 => n280, B1 => 
                           coeff_memory_2_10_port, B2 => n673, Z => N2987);
   U975 : AO22D1 port map( A1 => operand_regs_170_port, A2 => n282, B1 => 
                           coeff_memory_1_10_port, B2 => n673, Z => N2955);
   U976 : AO22D1 port map( A1 => coeff_memory_4_10_port, A2 => n673, B1 => n274
                           , B2 => operand_regs_10_port, Z => N3051);
   U977 : AO22D1 port map( A1 => coeff_memory_0_10_port, A2 => n673, B1 => n273
                           , B2 => operand_regs_234_port, Z => N2923);
   U978 : AO22D1 port map( A1 => n673, A2 => operand_regs_202_port, B1 => n271,
                           B2 => operand_regs_10_port, Z => N3211);
   U979 : OAI21M20D1 port map( A1 => operand_regs_73_port, A2 => n285, B => 
                           n144, Z => N3146);
   U980 : OAI21M20D1 port map( A1 => operand_regs_137_port, A2 => n284, B => 
                           n144, Z => N3114);
   U981 : OAI21M20D1 port map( A1 => n287, A2 => operand_regs_201_port, B => 
                           n144, Z => N3082);
   U982 : AO22D1 port map( A1 => operand_regs_43_port, A2 => n276, B1 => 
                           coeff_memory_3_11_port, B2 => n673, Z => N3020);
   U983 : AO22D1 port map( A1 => operand_regs_107_port, A2 => n280, B1 => 
                           coeff_memory_2_11_port, B2 => n673, Z => N2988);
   U984 : AO22D1 port map( A1 => operand_regs_171_port, A2 => n282, B1 => 
                           coeff_memory_1_11_port, B2 => n673, Z => N2956);
   U985 : AO22D1 port map( A1 => coeff_memory_4_11_port, A2 => n673, B1 => n271
                           , B2 => operand_regs_11_port, Z => N3052);
   U986 : AO22D1 port map( A1 => coeff_memory_0_11_port, A2 => n673, B1 => n273
                           , B2 => operand_regs_235_port, Z => N2924);
   U987 : AO22D1 port map( A1 => n673, A2 => operand_regs_204_port, B1 => n271,
                           B2 => operand_regs_12_port, Z => N3213);
   U988 : AO22D1 port map( A1 => n673, A2 => operand_regs_203_port, B1 => n271,
                           B2 => operand_regs_11_port, Z => N3212);
   U989 : NAN2D1 port map( A1 => operand_regs_233_port, A2 => n673, Z => n144);
   U990 : OAI21M20D1 port map( A1 => operand_regs_74_port, A2 => n285, B => 
                           n143, Z => N3147);
   U991 : OAI21M20D1 port map( A1 => operand_regs_138_port, A2 => n284, B => 
                           n143, Z => N3115);
   U992 : OAI21M20D1 port map( A1 => n287, A2 => operand_regs_202_port, B => 
                           n143, Z => N3083);
   U993 : AO22D1 port map( A1 => operand_regs_44_port, A2 => n281, B1 => 
                           coeff_memory_3_12_port, B2 => n673, Z => N3021);
   U994 : AO22D1 port map( A1 => operand_regs_108_port, A2 => n280, B1 => 
                           coeff_memory_2_12_port, B2 => n673, Z => N2989);
   U995 : AO22D1 port map( A1 => operand_regs_172_port, A2 => n282, B1 => 
                           coeff_memory_1_12_port, B2 => n673, Z => N2957);
   U996 : AO22D1 port map( A1 => coeff_memory_4_12_port, A2 => n673, B1 => n287
                           , B2 => operand_regs_12_port, Z => N3053);
   U997 : AO22D1 port map( A1 => coeff_memory_0_12_port, A2 => n673, B1 => n273
                           , B2 => operand_regs_236_port, Z => N2925);
   U998 : NAN2D1 port map( A1 => operand_regs_234_port, A2 => n673, Z => n143);
   U999 : OAI21M20D1 port map( A1 => operand_regs_75_port, A2 => n287, B => 
                           n142, Z => N3148);
   U1000 : OAI21M20D1 port map( A1 => operand_regs_139_port, A2 => n284, B => 
                           n142, Z => N3116);
   U1001 : OAI21M20D1 port map( A1 => operand_regs_76_port, A2 => n287, B => 
                           n141, Z => N3149);
   U1002 : OAI21M20D1 port map( A1 => operand_regs_140_port, A2 => n284, B => 
                           n141, Z => N3117);
   U1003 : OAI21M20D1 port map( A1 => n287, A2 => operand_regs_203_port, B => 
                           n142, Z => N3084);
   U1004 : OAI21M20D1 port map( A1 => n287, A2 => operand_regs_204_port, B => 
                           n141, Z => N3085);
   U1005 : AO22D1 port map( A1 => operand_regs_45_port, A2 => n276, B1 => 
                           coeff_memory_3_13_port, B2 => n673, Z => N3022);
   U1006 : AO22D1 port map( A1 => operand_regs_109_port, A2 => n280, B1 => 
                           coeff_memory_2_13_port, B2 => n673, Z => N2990);
   U1007 : AO22D1 port map( A1 => operand_regs_173_port, A2 => n282, B1 => 
                           coeff_memory_1_13_port, B2 => n673, Z => N2958);
   U1008 : AO22D1 port map( A1 => coeff_memory_4_13_port, A2 => n673, B1 => 
                           n275, B2 => operand_regs_13_port, Z => N3054);
   U1009 : AO22D1 port map( A1 => coeff_memory_0_13_port, A2 => n673, B1 => 
                           n273, B2 => operand_regs_237_port, Z => N2926);
   U1010 : NAN2D1 port map( A1 => operand_regs_235_port, A2 => n673, Z => n142)
                           ;
   U1011 : NAN2D1 port map( A1 => operand_regs_236_port, A2 => n673, Z => n141)
                           ;
   U1012 : AO22D1 port map( A1 => n673, A2 => operand_regs_205_port, B1 => n287
                           , B2 => operand_regs_13_port, Z => N3214);
   U1013 : AO22D1 port map( A1 => n673, A2 => operand_regs_206_port, B1 => n271
                           , B2 => operand_regs_14_port, Z => N3215);
   U1014 : AO22D1 port map( A1 => operand_regs_46_port, A2 => n278, B1 => 
                           coeff_memory_3_14_port, B2 => n673, Z => N3023);
   U1015 : AO22D1 port map( A1 => operand_regs_110_port, A2 => n279, B1 => 
                           coeff_memory_2_14_port, B2 => n673, Z => N2991);
   U1016 : AO22D1 port map( A1 => operand_regs_174_port, A2 => n282, B1 => 
                           coeff_memory_1_14_port, B2 => n673, Z => N2959);
   U1017 : AO22D1 port map( A1 => coeff_memory_4_14_port, A2 => n673, B1 => 
                           n276, B2 => operand_regs_14_port, Z => N3055);
   U1018 : AO22D1 port map( A1 => coeff_memory_0_14_port, A2 => n673, B1 => 
                           n287, B2 => operand_regs_238_port, Z => N2927);
   U1019 : OAI21M20D1 port map( A1 => operand_regs_77_port, A2 => n287, B => 
                           n140, Z => N3150);
   U1020 : OAI21M20D1 port map( A1 => operand_regs_141_port, A2 => n284, B => 
                           n140, Z => N3118);
   U1021 : OAI21M20D1 port map( A1 => operand_regs_78_port, A2 => n287, B => 
                           n139, Z => N3151);
   U1022 : OAI21M20D1 port map( A1 => operand_regs_142_port, A2 => n284, B => 
                           n139, Z => N3119);
   U1023 : OAI21M20D1 port map( A1 => n287, A2 => operand_regs_205_port, B => 
                           n140, Z => N3086);
   U1024 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_206_port, B => 
                           n139, Z => N3087);
   U1025 : AO22D1 port map( A1 => operand_regs_47_port, A2 => n278, B1 => 
                           coeff_memory_3_15_port, B2 => n673, Z => N3024);
   U1026 : AO22D1 port map( A1 => operand_regs_111_port, A2 => n277, B1 => 
                           coeff_memory_2_15_port, B2 => n673, Z => N2992);
   U1027 : AO22D1 port map( A1 => operand_regs_175_port, A2 => n278, B1 => 
                           coeff_memory_1_15_port, B2 => n673, Z => N2960);
   U1028 : AO22D1 port map( A1 => n673, A2 => operand_regs_207_port, B1 => n272
                           , B2 => operand_regs_15_port, Z => N3216);
   U1029 : AO22D1 port map( A1 => coeff_memory_4_15_port, A2 => n673, B1 => 
                           n275, B2 => operand_regs_15_port, Z => N3056);
   U1030 : AO22D1 port map( A1 => coeff_memory_0_15_port, A2 => n673, B1 => 
                           n287, B2 => operand_regs_239_port, Z => N2928);
   U1031 : NAN2D1 port map( A1 => operand_regs_237_port, A2 => n673, Z => n140)
                           ;
   U1032 : NAN2D1 port map( A1 => operand_regs_238_port, A2 => n673, Z => n139)
                           ;
   U1033 : OAI21M20D1 port map( A1 => operand_regs_79_port, A2 => n287, B => 
                           n138, Z => N3152);
   U1034 : OAI21M20D1 port map( A1 => operand_regs_143_port, A2 => n284, B => 
                           n138, Z => N3120);
   U1035 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_207_port, B => 
                           n138, Z => N3088);
   U1036 : AO22D1 port map( A1 => operand_regs_48_port, A2 => n281, B1 => 
                           coeff_memory_3_16_port, B2 => n673, Z => N3025);
   U1037 : AO22D1 port map( A1 => operand_regs_112_port, A2 => n277, B1 => 
                           coeff_memory_2_16_port, B2 => n673, Z => N2993);
   U1038 : AO22D1 port map( A1 => operand_regs_176_port, A2 => n282, B1 => 
                           coeff_memory_1_16_port, B2 => n673, Z => N2961);
   U1039 : AO22D1 port map( A1 => coeff_memory_4_16_port, A2 => n673, B1 => 
                           n276, B2 => operand_regs_16_port, Z => N3057);
   U1040 : AO22D1 port map( A1 => coeff_memory_0_16_port, A2 => n673, B1 => 
                           n287, B2 => operand_regs_240_port, Z => N2929);
   U1041 : AO22D1 port map( A1 => n673, A2 => operand_regs_208_port, B1 => n271
                           , B2 => operand_regs_16_port, Z => N3217);
   U1042 : NAN2D1 port map( A1 => operand_regs_239_port, A2 => n673, Z => n138)
                           ;
   U1043 : AO22D1 port map( A1 => operand_regs_49_port, A2 => n281, B1 => 
                           coeff_memory_3_17_port, B2 => n673, Z => N3026);
   U1044 : AO22D1 port map( A1 => operand_regs_113_port, A2 => n277, B1 => 
                           coeff_memory_2_17_port, B2 => n673, Z => N2994);
   U1045 : AO22D1 port map( A1 => operand_regs_177_port, A2 => n282, B1 => 
                           coeff_memory_1_17_port, B2 => n673, Z => N2962);
   U1046 : AO22D1 port map( A1 => coeff_memory_4_17_port, A2 => n673, B1 => 
                           n276, B2 => operand_regs_17_port, Z => N3058);
   U1047 : AO22D1 port map( A1 => coeff_memory_0_17_port, A2 => n673, B1 => 
                           n287, B2 => operand_regs_241_port, Z => N2930);
   U1048 : OAI21M20D1 port map( A1 => operand_regs_80_port, A2 => n287, B => 
                           n137, Z => N3153);
   U1049 : OAI21M20D1 port map( A1 => operand_regs_144_port, A2 => n284, B => 
                           n137, Z => N3121);
   U1050 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_208_port, B => 
                           n137, Z => N3089);
   U1051 : AO22D1 port map( A1 => operand_regs_50_port, A2 => n281, B1 => 
                           coeff_memory_3_18_port, B2 => n673, Z => N3027);
   U1052 : AO22D1 port map( A1 => operand_regs_114_port, A2 => n277, B1 => 
                           coeff_memory_2_18_port, B2 => n673, Z => N2995);
   U1053 : AO22D1 port map( A1 => operand_regs_178_port, A2 => n282, B1 => 
                           coeff_memory_1_18_port, B2 => n673, Z => N2963);
   U1054 : AO22D1 port map( A1 => coeff_memory_4_18_port, A2 => n673, B1 => 
                           n275, B2 => operand_regs_18_port, Z => N3059);
   U1055 : AO22D1 port map( A1 => coeff_memory_0_18_port, A2 => n673, B1 => 
                           n283, B2 => operand_regs_242_port, Z => N2931);
   U1056 : AO22D1 port map( A1 => n673, A2 => operand_regs_209_port, B1 => n272
                           , B2 => operand_regs_17_port, Z => N3218);
   U1057 : AO22D1 port map( A1 => operand_regs_51_port, A2 => n281, B1 => 
                           coeff_memory_3_19_port, B2 => n673, Z => N3028);
   U1058 : AO22D1 port map( A1 => operand_regs_115_port, A2 => n277, B1 => 
                           coeff_memory_2_19_port, B2 => n673, Z => N2996);
   U1059 : AO22D1 port map( A1 => operand_regs_179_port, A2 => n282, B1 => 
                           coeff_memory_1_19_port, B2 => n673, Z => N2964);
   U1060 : NAN2D1 port map( A1 => operand_regs_240_port, A2 => n673, Z => n137)
                           ;
   U1061 : AO22D1 port map( A1 => coeff_memory_0_19_port, A2 => n673, B1 => 
                           n274, B2 => operand_regs_243_port, Z => N2932);
   U1062 : AO22D1 port map( A1 => coeff_memory_4_19_port, A2 => n673, B1 => 
                           n276, B2 => operand_regs_19_port, Z => N3060);
   U1063 : OAI21M20D1 port map( A1 => operand_regs_81_port, A2 => n287, B => 
                           n136, Z => N3154);
   U1064 : OAI21M20D1 port map( A1 => operand_regs_145_port, A2 => n284, B => 
                           n136, Z => N3122);
   U1065 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_209_port, B => 
                           n136, Z => N3090);
   U1066 : AO22D1 port map( A1 => n673, A2 => operand_regs_210_port, B1 => n271
                           , B2 => operand_regs_18_port, Z => N3219);
   U1067 : NAN2D1 port map( A1 => operand_regs_241_port, A2 => n673, Z => n136)
                           ;
   U1068 : OAI21M20D1 port map( A1 => operand_regs_82_port, A2 => n282, B => 
                           n135, Z => N3155);
   U1069 : OAI21M20D1 port map( A1 => operand_regs_146_port, A2 => n287, B => 
                           n135, Z => N3123);
   U1070 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_210_port, B => 
                           n135, Z => N3091);
   U1071 : AO22D1 port map( A1 => n673, A2 => operand_regs_211_port, B1 => n277
                           , B2 => operand_regs_19_port, Z => N3220);
   U1072 : AO22D1 port map( A1 => n673, A2 => operand_regs_212_port, B1 => n271
                           , B2 => operand_regs_20_port, Z => N3221);
   U1073 : AO22D1 port map( A1 => operand_regs_52_port, A2 => n281, B1 => 
                           coeff_memory_3_20_port, B2 => n673, Z => N3029);
   U1074 : AO22D1 port map( A1 => operand_regs_116_port, A2 => n277, B1 => 
                           coeff_memory_2_20_port, B2 => n673, Z => N2997);
   U1075 : AO22D1 port map( A1 => operand_regs_180_port, A2 => n282, B1 => 
                           coeff_memory_1_20_port, B2 => n673, Z => N2965);
   U1076 : AO22D1 port map( A1 => coeff_memory_4_20_port, A2 => n673, B1 => 
                           n276, B2 => operand_regs_20_port, Z => N3061);
   U1077 : AO22D1 port map( A1 => coeff_memory_0_20_port, A2 => n673, B1 => 
                           n274, B2 => operand_regs_244_port, Z => N2933);
   U1078 : NAN2D1 port map( A1 => operand_regs_242_port, A2 => n673, Z => n135)
                           ;
   U1079 : OAI21M20D1 port map( A1 => operand_regs_83_port, A2 => n287, B => 
                           n134, Z => N3156);
   U1080 : OAI21M20D1 port map( A1 => operand_regs_147_port, A2 => n287, B => 
                           n134, Z => N3124);
   U1081 : OAI21M20D1 port map( A1 => operand_regs_84_port, A2 => n283, B => 
                           n133, Z => N3157);
   U1082 : OAI21M20D1 port map( A1 => operand_regs_148_port, A2 => n277, B => 
                           n133, Z => N3125);
   U1083 : AO22D1 port map( A1 => operand_regs_53_port, A2 => n281, B1 => 
                           coeff_memory_3_21_port, B2 => n673, Z => N3030);
   U1084 : AO22D1 port map( A1 => operand_regs_117_port, A2 => n277, B1 => 
                           coeff_memory_2_21_port, B2 => n673, Z => N2998);
   U1085 : AO22D1 port map( A1 => operand_regs_181_port, A2 => n279, B1 => 
                           coeff_memory_1_21_port, B2 => n673, Z => N2966);
   U1086 : OAI21M20D1 port map( A1 => n287, A2 => operand_regs_211_port, B => 
                           n134, Z => N3092);
   U1087 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_212_port, B => 
                           n133, Z => N3093);
   U1088 : AO22D1 port map( A1 => coeff_memory_4_21_port, A2 => n673, B1 => 
                           n275, B2 => operand_regs_21_port, Z => N3062);
   U1089 : AO22D1 port map( A1 => coeff_memory_0_21_port, A2 => n673, B1 => 
                           n274, B2 => operand_regs_245_port, Z => N2934);
   U1090 : NAN2D1 port map( A1 => operand_regs_243_port, A2 => n673, Z => n134)
                           ;
   U1091 : NAN2D1 port map( A1 => operand_regs_244_port, A2 => n673, Z => n133)
                           ;
   U1092 : AO22D1 port map( A1 => n673, A2 => operand_regs_213_port, B1 => n273
                           , B2 => operand_regs_21_port, Z => N3222);
   U1093 : AO22D1 port map( A1 => n673, A2 => operand_regs_214_port, B1 => n273
                           , B2 => operand_regs_22_port, Z => N3223);
   U1094 : AO22D1 port map( A1 => operand_regs_54_port, A2 => n283, B1 => 
                           coeff_memory_3_22_port, B2 => n673, Z => N3031);
   U1095 : AO22D1 port map( A1 => operand_regs_118_port, A2 => n277, B1 => 
                           coeff_memory_2_22_port, B2 => n673, Z => N2999);
   U1096 : AO22D1 port map( A1 => operand_regs_182_port, A2 => n279, B1 => 
                           coeff_memory_1_22_port, B2 => n673, Z => N2967);
   U1097 : AO22D1 port map( A1 => coeff_memory_4_22_port, A2 => n673, B1 => 
                           n275, B2 => operand_regs_22_port, Z => N3063);
   U1098 : AO22D1 port map( A1 => coeff_memory_0_22_port, A2 => n673, B1 => 
                           n274, B2 => operand_regs_246_port, Z => N2935);
   U1099 : OAI21M20D1 port map( A1 => operand_regs_85_port, A2 => n282, B => 
                           n132, Z => N3158);
   U1100 : OAI21M20D1 port map( A1 => operand_regs_149_port, A2 => n287, B => 
                           n132, Z => N3126);
   U1101 : OAI21M20D1 port map( A1 => operand_regs_86_port, A2 => n287, B => 
                           n131, Z => N3159);
   U1102 : OAI21M20D1 port map( A1 => operand_regs_150_port, A2 => n283, B => 
                           n131, Z => N3127);
   U1103 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_213_port, B => 
                           n132, Z => N3094);
   U1104 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_214_port, B => 
                           n131, Z => N3095);
   U1105 : AO22D1 port map( A1 => operand_regs_55_port, A2 => n283, B1 => 
                           coeff_memory_3_23_port, B2 => n673, Z => N3032);
   U1106 : AO22D1 port map( A1 => operand_regs_119_port, A2 => n277, B1 => 
                           coeff_memory_2_23_port, B2 => n673, Z => N3000);
   U1107 : AO22D1 port map( A1 => operand_regs_183_port, A2 => n279, B1 => 
                           coeff_memory_1_23_port, B2 => n673, Z => N2968);
   U1108 : AO22D1 port map( A1 => coeff_memory_4_23_port, A2 => n673, B1 => 
                           n275, B2 => operand_regs_23_port, Z => N3064);
   U1109 : AO22D1 port map( A1 => coeff_memory_0_23_port, A2 => n673, B1 => 
                           n274, B2 => operand_regs_247_port, Z => N2936);
   U1110 : AO22D1 port map( A1 => n673, A2 => operand_regs_215_port, B1 => n287
                           , B2 => operand_regs_23_port, Z => N3224);
   U1111 : NAN2D1 port map( A1 => operand_regs_245_port, A2 => n673, Z => n132)
                           ;
   U1112 : NAN2D1 port map( A1 => operand_regs_246_port, A2 => n673, Z => n131)
                           ;
   U1113 : OAI21M20D1 port map( A1 => operand_regs_87_port, A2 => n283, B => 
                           n130, Z => N3160);
   U1114 : OAI21M20D1 port map( A1 => operand_regs_151_port, A2 => n287, B => 
                           n130, Z => N3128);
   U1115 : OAI21M20D1 port map( A1 => n283, A2 => operand_regs_215_port, B => 
                           n130, Z => N3096);
   U1116 : AO22D1 port map( A1 => operand_regs_56_port, A2 => n283, B1 => 
                           coeff_memory_3_24_port, B2 => n673, Z => N3033);
   U1117 : AO22D1 port map( A1 => operand_regs_120_port, A2 => n277, B1 => 
                           coeff_memory_2_24_port, B2 => n673, Z => N3001);
   U1118 : AO22D1 port map( A1 => operand_regs_184_port, A2 => n279, B1 => 
                           coeff_memory_1_24_port, B2 => n673, Z => N2969);
   U1119 : AO22D1 port map( A1 => n673, A2 => operand_regs_216_port, B1 => n273
                           , B2 => operand_regs_24_port, Z => N3225);
   U1120 : AO22D1 port map( A1 => coeff_memory_4_24_port, A2 => n673, B1 => 
                           n287, B2 => operand_regs_24_port, Z => N3065);
   U1121 : AO22D1 port map( A1 => coeff_memory_0_24_port, A2 => n673, B1 => 
                           n274, B2 => operand_regs_248_port, Z => N2937);
   U1122 : NAN2D1 port map( A1 => operand_regs_247_port, A2 => n673, Z => n130)
                           ;
   U1123 : OAI21M20D1 port map( A1 => operand_regs_88_port, A2 => n282, B => 
                           n129, Z => N3161);
   U1124 : OAI21M20D1 port map( A1 => operand_regs_152_port, A2 => n287, B => 
                           n129, Z => N3129);
   U1125 : OAI21M20D1 port map( A1 => n287, A2 => operand_regs_216_port, B => 
                           n129, Z => N3097);
   U1126 : AO22D1 port map( A1 => operand_regs_57_port, A2 => n283, B1 => 
                           coeff_memory_3_25_port, B2 => n673, Z => N3034);
   U1127 : AO22D1 port map( A1 => operand_regs_121_port, A2 => n277, B1 => 
                           coeff_memory_2_25_port, B2 => n673, Z => N3002);
   U1128 : AO22D1 port map( A1 => operand_regs_185_port, A2 => n279, B1 => 
                           coeff_memory_1_25_port, B2 => n673, Z => N2970);
   U1129 : AO22D1 port map( A1 => coeff_memory_4_25_port, A2 => n673, B1 => 
                           n277, B2 => operand_regs_25_port, Z => N3066);
   U1130 : AO22D1 port map( A1 => coeff_memory_0_25_port, A2 => n673, B1 => 
                           n274, B2 => operand_regs_249_port, Z => N2938);
   U1131 : AO22D1 port map( A1 => n673, A2 => operand_regs_217_port, B1 => n283
                           , B2 => operand_regs_25_port, Z => N3226);
   U1132 : NAN2D1 port map( A1 => operand_regs_248_port, A2 => n673, Z => n129)
                           ;
   U1133 : OAI21M20D1 port map( A1 => operand_regs_89_port, A2 => n277, B => 
                           n128, Z => N3162);
   U1134 : OAI21M20D1 port map( A1 => operand_regs_153_port, A2 => n287, B => 
                           n128, Z => N3130);
   U1135 : OAI21M20D1 port map( A1 => n282, A2 => operand_regs_217_port, B => 
                           n128, Z => N3098);
   U1136 : AO22D1 port map( A1 => operand_regs_58_port, A2 => n283, B1 => 
                           coeff_memory_3_26_port, B2 => n673, Z => N3035);
   U1137 : AO22D1 port map( A1 => operand_regs_122_port, A2 => n276, B1 => 
                           coeff_memory_2_26_port, B2 => n673, Z => N3003);
   U1138 : AO22D1 port map( A1 => operand_regs_186_port, A2 => n279, B1 => 
                           coeff_memory_1_26_port, B2 => n673, Z => N2971);
   U1139 : AO22D1 port map( A1 => coeff_memory_4_26_port, A2 => n673, B1 => 
                           n283, B2 => operand_regs_26_port, Z => N3067);
   U1140 : AO22D1 port map( A1 => coeff_memory_0_26_port, A2 => n673, B1 => 
                           n287, B2 => operand_regs_250_port, Z => N2939);
   U1141 : AO22D1 port map( A1 => n673, A2 => operand_regs_218_port, B1 => n273
                           , B2 => operand_regs_26_port, Z => N3227);
   U1142 : NAN2D1 port map( A1 => operand_regs_249_port, A2 => n673, Z => n128)
                           ;
   U1143 : AO22D1 port map( A1 => operand_regs_59_port, A2 => n283, B1 => 
                           coeff_memory_3_27_port, B2 => n673, Z => N3036);
   U1144 : AO22D1 port map( A1 => operand_regs_123_port, A2 => n278, B1 => 
                           coeff_memory_2_27_port, B2 => n673, Z => N3004);
   U1145 : AO22D1 port map( A1 => operand_regs_187_port, A2 => n279, B1 => 
                           coeff_memory_1_27_port, B2 => n673, Z => N2972);
   U1146 : OAI21M20D1 port map( A1 => operand_regs_90_port, A2 => n287, B => 
                           n127, Z => N3163);
   U1147 : OAI21M20D1 port map( A1 => operand_regs_154_port, A2 => n287, B => 
                           n127, Z => N3131);
   U1148 : OAI21M20D1 port map( A1 => n283, A2 => operand_regs_218_port, B => 
                           n127, Z => N3099);
   U1149 : AO22D1 port map( A1 => coeff_memory_4_27_port, A2 => n673, B1 => 
                           n287, B2 => operand_regs_27_port, Z => N3068);
   U1150 : AO22D1 port map( A1 => coeff_memory_0_27_port, A2 => n673, B1 => 
                           n283, B2 => operand_regs_251_port, Z => N2940);
   U1151 : AO22D1 port map( A1 => operand_regs_60_port, A2 => n283, B1 => 
                           coeff_memory_3_28_port, B2 => n673, Z => N3037);
   U1152 : AO22D1 port map( A1 => operand_regs_124_port, A2 => n278, B1 => 
                           coeff_memory_2_28_port, B2 => n673, Z => N3005);
   U1153 : AO22D1 port map( A1 => operand_regs_188_port, A2 => n279, B1 => 
                           coeff_memory_1_28_port, B2 => n673, Z => N2973);
   U1154 : NAN2D1 port map( A1 => operand_regs_250_port, A2 => n673, Z => n127)
                           ;
   U1155 : AO22D1 port map( A1 => n673, A2 => operand_regs_219_port, B1 => n277
                           , B2 => operand_regs_27_port, Z => N3228);
   U1156 : AO22D1 port map( A1 => coeff_memory_4_28_port, A2 => n673, B1 => 
                           n283, B2 => operand_regs_28_port, Z => N3069);
   U1157 : AO22D1 port map( A1 => coeff_memory_0_28_port, A2 => n673, B1 => 
                           n282, B2 => operand_regs_252_port, Z => N2941);
   U1158 : OAI21M20D1 port map( A1 => operand_regs_91_port, A2 => n283, B => 
                           n126, Z => N3164);
   U1159 : OAI21M20D1 port map( A1 => operand_regs_155_port, A2 => n283, B => 
                           n126, Z => N3132);
   U1160 : AO22D1 port map( A1 => operand_regs_61_port, A2 => n283, B1 => 
                           coeff_memory_3_29_port, B2 => n673, Z => N3038);
   U1161 : AO22D1 port map( A1 => operand_regs_125_port, A2 => n278, B1 => 
                           coeff_memory_2_29_port, B2 => n673, Z => N3006);
   U1162 : AO22D1 port map( A1 => operand_regs_189_port, A2 => n279, B1 => 
                           coeff_memory_1_29_port, B2 => n673, Z => N2974);
   U1163 : OAI21M20D1 port map( A1 => n287, A2 => operand_regs_219_port, B => 
                           n126, Z => N3100);
   U1164 : AO22D1 port map( A1 => coeff_memory_4_29_port, A2 => n673, B1 => 
                           n287, B2 => operand_regs_29_port, Z => N3070);
   U1165 : AO22D1 port map( A1 => coeff_memory_0_29_port, A2 => n673, B1 => 
                           n287, B2 => operand_regs_253_port, Z => N2942);
   U1166 : AO22D1 port map( A1 => n673, A2 => operand_regs_220_port, B1 => n273
                           , B2 => operand_regs_28_port, Z => N3229);
   U1167 : NAN2D1 port map( A1 => operand_regs_251_port, A2 => n673, Z => n126)
                           ;
   U1168 : OAI21M20D1 port map( A1 => operand_regs_92_port, A2 => n287, B => 
                           n125, Z => N3165);
   U1169 : OAI21M20D1 port map( A1 => operand_regs_156_port, A2 => n277, B => 
                           n125, Z => N3133);
   U1170 : OAI21M20D1 port map( A1 => n283, A2 => operand_regs_220_port, B => 
                           n125, Z => N3101);
   U1171 : AO22D1 port map( A1 => operand_regs_62_port, A2 => n283, B1 => 
                           coeff_memory_3_30_port, B2 => n673, Z => N3039);
   U1172 : AO22D1 port map( A1 => operand_regs_126_port, A2 => n278, B1 => 
                           coeff_memory_2_30_port, B2 => n673, Z => N3007);
   U1173 : AO22D1 port map( A1 => operand_regs_190_port, A2 => n279, B1 => 
                           coeff_memory_1_30_port, B2 => n673, Z => N2975);
   U1174 : NAN2D1 port map( A1 => operand_regs_252_port, A2 => n673, Z => n125)
                           ;
   U1175 : AO22D1 port map( A1 => coeff_memory_4_30_port, A2 => n673, B1 => 
                           n282, B2 => operand_regs_30_port, Z => N3071);
   U1176 : AO22D1 port map( A1 => coeff_memory_0_30_port, A2 => n673, B1 => 
                           n283, B2 => operand_regs_254_port, Z => N2943);
   U1177 : AO22D1 port map( A1 => n673, A2 => operand_regs_221_port, B1 => n272
                           , B2 => operand_regs_29_port, Z => N3230);
   U1178 : AO22D1 port map( A1 => n673, A2 => operand_regs_222_port, B1 => n283
                           , B2 => operand_regs_30_port, Z => N3231);
   U1179 : OAI21M20D1 port map( A1 => operand_regs_93_port, A2 => n287, B => 
                           n124, Z => N3166);
   U1180 : OAI21M20D1 port map( A1 => operand_regs_157_port, A2 => n287, B => 
                           n124, Z => N3134);
   U1181 : OAI21M20D1 port map( A1 => operand_regs_94_port, A2 => n283, B => 
                           n123, Z => N3167);
   U1182 : OAI21M20D1 port map( A1 => operand_regs_158_port, A2 => n287, B => 
                           n123, Z => N3135);
   U1183 : OAI21M20D1 port map( A1 => n277, A2 => operand_regs_221_port, B => 
                           n124, Z => N3102);
   U1184 : OAI21M20D1 port map( A1 => n283, A2 => operand_regs_222_port, B => 
                           n123, Z => N3103);
   U1185 : AO22D1 port map( A1 => operand_regs_63_port, A2 => n283, B1 => 
                           coeff_memory_3_31_port, B2 => n673, Z => N3040);
   U1186 : AO22D1 port map( A1 => operand_regs_127_port, A2 => n280, B1 => 
                           coeff_memory_2_31_port, B2 => n673, Z => N3008);
   U1187 : AO22D1 port map( A1 => operand_regs_191_port, A2 => n279, B1 => 
                           coeff_memory_1_31_port, B2 => n673, Z => N2976);
   U1188 : AO22D1 port map( A1 => coeff_memory_4_31_port, A2 => n673, B1 => 
                           n287, B2 => operand_regs_31_port, Z => N3072);
   U1189 : AO22D1 port map( A1 => coeff_memory_0_31_port, A2 => n673, B1 => 
                           n282, B2 => operand_regs_255_port, Z => N2944);
   U1190 : NAN2D1 port map( A1 => operand_regs_253_port, A2 => n673, Z => n124)
                           ;
   U1191 : NAN2D1 port map( A1 => operand_regs_254_port, A2 => n673, Z => n123)
                           ;
   U1192 : OAI21M20D1 port map( A1 => operand_regs_95_port, A2 => n284, B => 
                           n122, Z => N3168);
   U1193 : OAI21M20D1 port map( A1 => operand_regs_159_port, A2 => n287, B => 
                           n122, Z => N3136);
   U1194 : OAI21M20D1 port map( A1 => n287, A2 => operand_regs_223_port, B => 
                           n122, Z => N3104);
   U1195 : AO22D1 port map( A1 => n673, A2 => operand_regs_223_port, B1 => n275
                           , B2 => operand_regs_31_port, Z => N3232);
   U1196 : NAN2D1 port map( A1 => operand_regs_255_port, A2 => n673, Z => n122)
                           ;
   U1197 : AO22D1 port map( A1 => N2876, A2 => n672, B1 => N2859, B2 => n696, Z
                           => N2894);
   U1198 : AO22D1 port map( A1 => N2875, A2 => n672, B1 => N2858, B2 => n696, Z
                           => N2895);
   U1199 : AO22D1 port map( A1 => N2874, A2 => n672, B1 => N2857, B2 => n696, Z
                           => N2896);
   U1200 : AO22D1 port map( A1 => N2873, A2 => n672, B1 => N2856, B2 => n696, Z
                           => N2897);
   U1201 : AO22D1 port map( A1 => N2872, A2 => n672, B1 => N2855, B2 => n696, Z
                           => N2898);
   U1202 : AO22D1 port map( A1 => N2871, A2 => n672, B1 => N2854, B2 => n696, Z
                           => N2899);
   U1203 : AO22D1 port map( A1 => N2870, A2 => n672, B1 => N2853, B2 => n696, Z
                           => N2900);
   U1204 : AO22D1 port map( A1 => N2869, A2 => n672, B1 => N2852, B2 => n696, Z
                           => N2901);
   U1205 : AO22D1 port map( A1 => N2868, A2 => n672, B1 => N2851, B2 => n696, Z
                           => N2902);
   U1206 : AO22D1 port map( A1 => N2867, A2 => n672, B1 => N2850, B2 => n696, Z
                           => N2903);
   U1207 : AO22D1 port map( A1 => N2881, A2 => n672, B1 => N2864, B2 => n696, Z
                           => N2889);
   U1208 : AO22D1 port map( A1 => N2880, A2 => n672, B1 => N2863, B2 => n696, Z
                           => N2890);
   U1209 : AO22D1 port map( A1 => N2879, A2 => n672, B1 => N2862, B2 => n696, Z
                           => N2891);
   U1210 : AO22D1 port map( A1 => N2878, A2 => n672, B1 => N2861, B2 => n696, Z
                           => N2892);
   U1211 : AO22D1 port map( A1 => N2877, A2 => n672, B1 => N2860, B2 => n696, Z
                           => N2893);
   U1212 : AO22D1 port map( A1 => N2882, A2 => n672, B1 => N2865, B2 => n696, Z
                           => N2888);
   U1213 : INVD1 port map( A => N64, Z => n671);
   U1214 : INVD1 port map( A => coeff_load, Z => n686);
   U1215 : NOR2D1 port map( A1 => n684, A2 => out_busy, Z => n79);
   U1216 : NAN3D1 port map( A1 => n81, A2 => out_busy, A3 => N62, Z => n4);
   U1217 : INVD1 port map( A => N62, Z => n694);
   U1218 : BUFD1 port map( A => odd1, Z => n672);
   U1219 : INVD1 port map( A => out_busy, Z => n695);
   U1220 : INVD1 port map( A => odd, Z => n687);
   U1221 : NAN3D1 port map( A1 => in_counter_1_port, A2 => in_busy, A3 => 
                           in_counter_0_port, Z => n88);
   U1222 : NOR2D1 port map( A1 => n690, A2 => in_counter_0_port, Z => n155);
   U1223 : OAI21M20D1 port map( A1 => n690, A2 => in_trigger, B => n100, Z => 
                           n84);
   U1224 : INVD1 port map( A => in_busy, Z => n690);
   U1225 : INVD1 port map( A => in_counter_2_port, Z => n693);
   U1226 : INVD1 port map( A => N63, Z => n697);
   U1227 : NOR2D1 port map( A1 => n688, A2 => in_counter_1_port, Z => n119);
   U1228 : NAN2D1 port map( A1 => in_counter_1_port, A2 => n155, Z => n85);
   U1229 : AND3D1 port map( A1 => in_counter_0_port, A2 => in_busy, A3 => n692,
                           Z => n87);
   U1230 : INVD1 port map( A => in_counter_1_port, Z => n692);
   U1231 : NAN2D1 port map( A1 => n78, A2 => n672, Z => n77);
   U1232 : NOR2D1 port map( A1 => n687, A2 => in_counter_2_port, Z => n101);
   U1233 : NOR2D1 port map( A1 => n693, A2 => odd, Z => n115);
   U1234 : NOR2D1 port map( A1 => odd, A2 => in_counter_2_port, Z => n120);
   U1235 : INVD1 port map( A => out_trigger, Z => n685);
   U1236 : NOR2D1 port map( A1 => n522, A2 => avs_addr(1), Z => n288);
   U1237 : NOR2D1 port map( A1 => n522, A2 => n680, Z => n289);
   U1238 : AOI22D1 port map( A1 => in_buf_64_port, A2 => n266, B1 => 
                           in_buf_0_port, B2 => n242, Z => n295);
   U1239 : NOR2D1 port map( A1 => avs_addr(1), A2 => avs_addr(2), Z => n290);
   U1240 : AND2D1 port map( A1 => n290, A2 => avs_addr(0), Z => n514);
   U1241 : NOR2D1 port map( A1 => n680, A2 => avs_addr(2), Z => n291);
   U1242 : AND2D1 port map( A1 => n291, A2 => avs_addr(0), Z => n513);
   U1243 : AOI22D1 port map( A1 => in_buf_192_port, A2 => n527, B1 => 
                           in_buf_128_port, B2 => n525, Z => n294);
   U1244 : NOR2M1D1 port map( A1 => n288, A2 => avs_addr(0), Z => n516);
   U1245 : NOR2M1D1 port map( A1 => n289, A2 => avs_addr(0), Z => n515);
   U1246 : AOI22D1 port map( A1 => in_buf_96_port, A2 => n529, B1 => 
                           in_buf_32_port, B2 => n515, Z => n293);
   U1247 : NOR2M1D1 port map( A1 => n290, A2 => avs_addr(0), Z => n518);
   U1248 : NOR2M1D1 port map( A1 => n291, A2 => avs_addr(0), Z => n517);
   U1249 : AOI22D1 port map( A1 => in_buf_224_port, A2 => n534, B1 => 
                           in_buf_160_port, B2 => n532, Z => n292);
   U1250 : NAN4D1 port map( A1 => n295, A2 => n294, A3 => n293, A4 => n292, Z 
                           => N2041);
   U1251 : AOI22D1 port map( A1 => in_buf_65_port, A2 => n266, B1 => 
                           in_buf_1_port, B2 => n242, Z => n299);
   U1252 : AOI22D1 port map( A1 => in_buf_193_port, A2 => n527, B1 => 
                           in_buf_129_port, B2 => n513, Z => n298);
   U1253 : AOI22D1 port map( A1 => in_buf_97_port, A2 => n529, B1 => 
                           in_buf_33_port, B2 => n515, Z => n297);
   U1254 : AOI22D1 port map( A1 => in_buf_225_port, A2 => n518, B1 => 
                           in_buf_161_port, B2 => n517, Z => n296);
   U1255 : NAN4D1 port map( A1 => n299, A2 => n298, A3 => n297, A4 => n296, Z 
                           => N2040);
   U1256 : AOI22D1 port map( A1 => in_buf_66_port, A2 => n266, B1 => 
                           in_buf_2_port, B2 => n242, Z => n303);
   U1257 : AOI22D1 port map( A1 => in_buf_194_port, A2 => n527, B1 => 
                           in_buf_130_port, B2 => n513, Z => n302);
   U1258 : AOI22D1 port map( A1 => in_buf_98_port, A2 => n529, B1 => 
                           in_buf_34_port, B2 => n515, Z => n301);
   U1259 : AOI22D1 port map( A1 => in_buf_226_port, A2 => n518, B1 => 
                           in_buf_162_port, B2 => n517, Z => n300);
   U1260 : NAN4D1 port map( A1 => n303, A2 => n302, A3 => n301, A4 => n300, Z 
                           => N2039);
   U1261 : AOI22D1 port map( A1 => in_buf_67_port, A2 => n266, B1 => 
                           in_buf_3_port, B2 => n242, Z => n307);
   U1262 : AOI22D1 port map( A1 => in_buf_195_port, A2 => n527, B1 => 
                           in_buf_131_port, B2 => n513, Z => n306);
   U1263 : AOI22D1 port map( A1 => in_buf_99_port, A2 => n529, B1 => 
                           in_buf_35_port, B2 => n515, Z => n305);
   U1264 : AOI22D1 port map( A1 => in_buf_227_port, A2 => n518, B1 => 
                           in_buf_163_port, B2 => n517, Z => n304);
   U1265 : NAN4D1 port map( A1 => n307, A2 => n306, A3 => n305, A4 => n304, Z 
                           => N2038);
   U1266 : AOI22D1 port map( A1 => in_buf_68_port, A2 => n266, B1 => 
                           in_buf_4_port, B2 => n242, Z => n311);
   U1267 : AOI22D1 port map( A1 => in_buf_196_port, A2 => n527, B1 => 
                           in_buf_132_port, B2 => n513, Z => n310);
   U1268 : AOI22D1 port map( A1 => in_buf_100_port, A2 => n529, B1 => 
                           in_buf_36_port, B2 => n515, Z => n309);
   U1269 : AOI22D1 port map( A1 => in_buf_228_port, A2 => n518, B1 => 
                           in_buf_164_port, B2 => n517, Z => n308);
   U1270 : NAN4D1 port map( A1 => n311, A2 => n310, A3 => n309, A4 => n308, Z 
                           => N2037);
   U1271 : AOI22D1 port map( A1 => in_buf_69_port, A2 => n266, B1 => 
                           in_buf_5_port, B2 => n242, Z => n315);
   U1272 : AOI22D1 port map( A1 => in_buf_197_port, A2 => n527, B1 => 
                           in_buf_133_port, B2 => n513, Z => n314);
   U1273 : AOI22D1 port map( A1 => in_buf_101_port, A2 => n529, B1 => 
                           in_buf_37_port, B2 => n515, Z => n313);
   U1274 : AOI22D1 port map( A1 => in_buf_229_port, A2 => n518, B1 => 
                           in_buf_165_port, B2 => n517, Z => n312);
   U1275 : NAN4D1 port map( A1 => n315, A2 => n314, A3 => n313, A4 => n312, Z 
                           => N2036);
   U1276 : AOI22D1 port map( A1 => in_buf_70_port, A2 => n266, B1 => 
                           in_buf_6_port, B2 => n242, Z => n319);
   U1277 : AOI22D1 port map( A1 => in_buf_198_port, A2 => n527, B1 => 
                           in_buf_134_port, B2 => n513, Z => n318);
   U1278 : AOI22D1 port map( A1 => in_buf_102_port, A2 => n529, B1 => 
                           in_buf_38_port, B2 => n515, Z => n317);
   U1279 : AOI22D1 port map( A1 => in_buf_230_port, A2 => n518, B1 => 
                           in_buf_166_port, B2 => n517, Z => n316);
   U1280 : NAN4D1 port map( A1 => n319, A2 => n318, A3 => n317, A4 => n316, Z 
                           => N2035);
   U1281 : AOI22D1 port map( A1 => in_buf_71_port, A2 => n266, B1 => 
                           in_buf_7_port, B2 => n242, Z => n323);
   U1282 : AOI22D1 port map( A1 => in_buf_199_port, A2 => n527, B1 => 
                           in_buf_135_port, B2 => n513, Z => n322);
   U1283 : AOI22D1 port map( A1 => in_buf_103_port, A2 => n529, B1 => 
                           in_buf_39_port, B2 => n515, Z => n321);
   U1284 : AOI22D1 port map( A1 => in_buf_231_port, A2 => n518, B1 => 
                           in_buf_167_port, B2 => n517, Z => n320);
   U1285 : NAN4D1 port map( A1 => n323, A2 => n322, A3 => n321, A4 => n320, Z 
                           => N2034);
   U1286 : AOI22D1 port map( A1 => in_buf_72_port, A2 => n266, B1 => 
                           in_buf_8_port, B2 => n242, Z => n327);
   U1287 : AOI22D1 port map( A1 => in_buf_200_port, A2 => n527, B1 => 
                           in_buf_136_port, B2 => n513, Z => n326);
   U1288 : AOI22D1 port map( A1 => in_buf_104_port, A2 => n516, B1 => 
                           in_buf_40_port, B2 => n515, Z => n325);
   U1289 : AOI22D1 port map( A1 => in_buf_232_port, A2 => n518, B1 => 
                           in_buf_168_port, B2 => n517, Z => n324);
   U1290 : NAN4D1 port map( A1 => n327, A2 => n326, A3 => n325, A4 => n324, Z 
                           => N2033);
   U1291 : AOI22D1 port map( A1 => in_buf_73_port, A2 => n266, B1 => 
                           in_buf_9_port, B2 => n242, Z => n331);
   U1292 : AOI22D1 port map( A1 => in_buf_201_port, A2 => n527, B1 => 
                           in_buf_137_port, B2 => n513, Z => n330);
   U1293 : AOI22D1 port map( A1 => in_buf_105_port, A2 => n516, B1 => 
                           in_buf_41_port, B2 => n515, Z => n329);
   U1294 : AOI22D1 port map( A1 => in_buf_233_port, A2 => n518, B1 => 
                           in_buf_169_port, B2 => n517, Z => n328);
   U1295 : NAN4D1 port map( A1 => n331, A2 => n330, A3 => n329, A4 => n328, Z 
                           => N2032);
   U1296 : AOI22D1 port map( A1 => in_buf_74_port, A2 => n266, B1 => 
                           in_buf_10_port, B2 => n242, Z => n335);
   U1297 : AOI22D1 port map( A1 => in_buf_202_port, A2 => n527, B1 => 
                           in_buf_138_port, B2 => n513, Z => n334);
   U1298 : AOI22D1 port map( A1 => in_buf_106_port, A2 => n516, B1 => 
                           in_buf_42_port, B2 => n515, Z => n333);
   U1299 : AOI22D1 port map( A1 => in_buf_234_port, A2 => n534, B1 => 
                           in_buf_170_port, B2 => n517, Z => n332);
   U1300 : NAN4D1 port map( A1 => n335, A2 => n334, A3 => n333, A4 => n332, Z 
                           => N2031);
   U1301 : AOI22D1 port map( A1 => in_buf_75_port, A2 => n266, B1 => 
                           in_buf_11_port, B2 => n242, Z => n339);
   U1302 : AOI22D1 port map( A1 => in_buf_203_port, A2 => n527, B1 => 
                           in_buf_139_port, B2 => n513, Z => n338);
   U1303 : AOI22D1 port map( A1 => in_buf_107_port, A2 => n516, B1 => 
                           in_buf_43_port, B2 => n515, Z => n337);
   U1304 : AOI22D1 port map( A1 => in_buf_235_port, A2 => n518, B1 => 
                           in_buf_171_port, B2 => n517, Z => n336);
   U1305 : NAN4D1 port map( A1 => n339, A2 => n338, A3 => n337, A4 => n336, Z 
                           => N2030);
   U1306 : AOI22D1 port map( A1 => in_buf_76_port, A2 => n266, B1 => 
                           in_buf_12_port, B2 => n242, Z => n343);
   U1307 : AOI22D1 port map( A1 => in_buf_204_port, A2 => n527, B1 => 
                           in_buf_140_port, B2 => n513, Z => n342);
   U1308 : AOI22D1 port map( A1 => in_buf_108_port, A2 => n529, B1 => 
                           in_buf_44_port, B2 => n515, Z => n341);
   U1309 : AOI22D1 port map( A1 => in_buf_236_port, A2 => n534, B1 => 
                           in_buf_172_port, B2 => n532, Z => n340);
   U1310 : NAN4D1 port map( A1 => n343, A2 => n342, A3 => n341, A4 => n340, Z 
                           => N2029);
   U1311 : AOI22D1 port map( A1 => in_buf_77_port, A2 => n266, B1 => 
                           in_buf_13_port, B2 => n242, Z => n347);
   U1312 : AOI22D1 port map( A1 => in_buf_205_port, A2 => n514, B1 => 
                           in_buf_141_port, B2 => n525, Z => n346);
   U1313 : AOI22D1 port map( A1 => in_buf_109_port, A2 => n516, B1 => 
                           in_buf_45_port, B2 => n515, Z => n345);
   U1314 : AOI22D1 port map( A1 => in_buf_237_port, A2 => n534, B1 => 
                           in_buf_173_port, B2 => n531, Z => n344);
   U1315 : NAN4D1 port map( A1 => n347, A2 => n346, A3 => n345, A4 => n344, Z 
                           => N2028);
   U1316 : AOI22D1 port map( A1 => in_buf_78_port, A2 => n266, B1 => 
                           in_buf_14_port, B2 => n242, Z => n351);
   U1317 : AOI22D1 port map( A1 => in_buf_206_port, A2 => n514, B1 => 
                           in_buf_142_port, B2 => n525, Z => n350);
   U1318 : AOI22D1 port map( A1 => in_buf_110_port, A2 => n516, B1 => 
                           in_buf_46_port, B2 => n515, Z => n349);
   U1319 : AOI22D1 port map( A1 => in_buf_238_port, A2 => n534, B1 => 
                           in_buf_174_port, B2 => n517, Z => n348);
   U1320 : NAN4D1 port map( A1 => n351, A2 => n350, A3 => n349, A4 => n348, Z 
                           => N2027);
   U1321 : AOI22D1 port map( A1 => in_buf_79_port, A2 => n266, B1 => 
                           in_buf_15_port, B2 => n242, Z => n355);
   U1322 : AOI22D1 port map( A1 => in_buf_207_port, A2 => n514, B1 => 
                           in_buf_143_port, B2 => n525, Z => n354);
   U1323 : AOI22D1 port map( A1 => in_buf_111_port, A2 => n516, B1 => 
                           in_buf_47_port, B2 => n515, Z => n353);
   U1324 : AOI22D1 port map( A1 => in_buf_239_port, A2 => n534, B1 => 
                           in_buf_175_port, B2 => n517, Z => n352);
   U1325 : NAN4D1 port map( A1 => n355, A2 => n354, A3 => n353, A4 => n352, Z 
                           => N2026);
   U1326 : AOI22D1 port map( A1 => in_buf_80_port, A2 => n266, B1 => 
                           in_buf_16_port, B2 => n242, Z => n359);
   U1327 : AOI22D1 port map( A1 => in_buf_208_port, A2 => n514, B1 => 
                           in_buf_144_port, B2 => n525, Z => n358);
   U1328 : AOI22D1 port map( A1 => in_buf_112_port, A2 => n516, B1 => 
                           in_buf_48_port, B2 => n515, Z => n357);
   U1329 : AOI22D1 port map( A1 => in_buf_240_port, A2 => n534, B1 => 
                           in_buf_176_port, B2 => n517, Z => n356);
   U1330 : NAN4D1 port map( A1 => n359, A2 => n358, A3 => n357, A4 => n356, Z 
                           => N2025);
   U1331 : AOI22D1 port map( A1 => in_buf_81_port, A2 => n266, B1 => 
                           in_buf_17_port, B2 => n242, Z => n363);
   U1332 : AOI22D1 port map( A1 => in_buf_209_port, A2 => n514, B1 => 
                           in_buf_145_port, B2 => n525, Z => n362);
   U1333 : AOI22D1 port map( A1 => in_buf_113_port, A2 => n516, B1 => 
                           in_buf_49_port, B2 => n515, Z => n361);
   U1334 : AOI22D1 port map( A1 => in_buf_241_port, A2 => n534, B1 => 
                           in_buf_177_port, B2 => n517, Z => n360);
   U1335 : NAN4D1 port map( A1 => n363, A2 => n362, A3 => n361, A4 => n360, Z 
                           => N2024);
   U1336 : AOI22D1 port map( A1 => in_buf_82_port, A2 => n266, B1 => 
                           in_buf_18_port, B2 => n242, Z => n367);
   U1337 : AOI22D1 port map( A1 => in_buf_210_port, A2 => n514, B1 => 
                           in_buf_146_port, B2 => n525, Z => n366);
   U1338 : AOI22D1 port map( A1 => in_buf_114_port, A2 => n516, B1 => 
                           in_buf_50_port, B2 => n515, Z => n365);
   U1339 : AOI22D1 port map( A1 => in_buf_242_port, A2 => n534, B1 => 
                           in_buf_178_port, B2 => n517, Z => n364);
   U1340 : NAN4D1 port map( A1 => n367, A2 => n366, A3 => n365, A4 => n364, Z 
                           => N2023);
   U1341 : AOI22D1 port map( A1 => in_buf_83_port, A2 => n266, B1 => 
                           in_buf_19_port, B2 => n242, Z => n371);
   U1342 : AOI22D1 port map( A1 => in_buf_211_port, A2 => n514, B1 => 
                           in_buf_147_port, B2 => n525, Z => n370);
   U1343 : AOI22D1 port map( A1 => in_buf_115_port, A2 => n516, B1 => 
                           in_buf_51_port, B2 => n515, Z => n369);
   U1344 : AOI22D1 port map( A1 => in_buf_243_port, A2 => n534, B1 => 
                           in_buf_179_port, B2 => n517, Z => n368);
   U1345 : NAN4D1 port map( A1 => n371, A2 => n370, A3 => n369, A4 => n368, Z 
                           => N2022);
   U1346 : AOI22D1 port map( A1 => in_buf_84_port, A2 => n266, B1 => 
                           in_buf_20_port, B2 => n242, Z => n375);
   U1347 : AOI22D1 port map( A1 => in_buf_212_port, A2 => n514, B1 => 
                           in_buf_148_port, B2 => n525, Z => n374);
   U1348 : AOI22D1 port map( A1 => in_buf_116_port, A2 => n516, B1 => 
                           in_buf_52_port, B2 => n515, Z => n373);
   U1349 : AOI22D1 port map( A1 => in_buf_244_port, A2 => n534, B1 => 
                           in_buf_180_port, B2 => n517, Z => n372);
   U1350 : NAN4D1 port map( A1 => n375, A2 => n374, A3 => n373, A4 => n372, Z 
                           => N2021);
   U1351 : AOI22D1 port map( A1 => in_buf_85_port, A2 => n266, B1 => 
                           in_buf_21_port, B2 => n242, Z => n379);
   U1352 : AOI22D1 port map( A1 => in_buf_213_port, A2 => n514, B1 => 
                           in_buf_149_port, B2 => n525, Z => n378);
   U1353 : AOI22D1 port map( A1 => in_buf_117_port, A2 => n516, B1 => 
                           in_buf_53_port, B2 => n515, Z => n377);
   U1354 : AOI22D1 port map( A1 => in_buf_245_port, A2 => n534, B1 => 
                           in_buf_181_port, B2 => n517, Z => n376);
   U1355 : NAN4D1 port map( A1 => n379, A2 => n378, A3 => n377, A4 => n376, Z 
                           => N2020);
   U1356 : AOI22D1 port map( A1 => in_buf_86_port, A2 => n266, B1 => 
                           in_buf_22_port, B2 => n242, Z => n383);
   U1357 : AOI22D1 port map( A1 => in_buf_214_port, A2 => n514, B1 => 
                           in_buf_150_port, B2 => n525, Z => n382);
   U1358 : AOI22D1 port map( A1 => in_buf_118_port, A2 => n516, B1 => 
                           in_buf_54_port, B2 => n515, Z => n381);
   U1359 : AOI22D1 port map( A1 => in_buf_246_port, A2 => n534, B1 => 
                           in_buf_182_port, B2 => n517, Z => n380);
   U1360 : NAN4D1 port map( A1 => n383, A2 => n382, A3 => n381, A4 => n380, Z 
                           => N2019);
   U1361 : AOI22D1 port map( A1 => in_buf_87_port, A2 => n266, B1 => 
                           in_buf_23_port, B2 => n242, Z => n387);
   U1362 : AOI22D1 port map( A1 => in_buf_215_port, A2 => n514, B1 => 
                           in_buf_151_port, B2 => n525, Z => n386);
   U1363 : AOI22D1 port map( A1 => in_buf_119_port, A2 => n516, B1 => 
                           in_buf_55_port, B2 => n515, Z => n385);
   U1364 : AOI22D1 port map( A1 => in_buf_247_port, A2 => n534, B1 => 
                           in_buf_183_port, B2 => n517, Z => n384);
   U1365 : NAN4D1 port map( A1 => n387, A2 => n386, A3 => n385, A4 => n384, Z 
                           => N2018);
   U1366 : AOI22D1 port map( A1 => in_buf_88_port, A2 => n266, B1 => 
                           in_buf_24_port, B2 => n242, Z => n391);
   U1367 : AOI22D1 port map( A1 => in_buf_216_port, A2 => n514, B1 => 
                           in_buf_152_port, B2 => n525, Z => n390);
   U1368 : AOI22D1 port map( A1 => in_buf_120_port, A2 => n516, B1 => 
                           in_buf_56_port, B2 => n515, Z => n389);
   U1369 : AOI22D1 port map( A1 => in_buf_248_port, A2 => n534, B1 => 
                           in_buf_184_port, B2 => n517, Z => n388);
   U1370 : NAN4D1 port map( A1 => n391, A2 => n390, A3 => n389, A4 => n388, Z 
                           => N2017);
   U1371 : AOI22D1 port map( A1 => in_buf_89_port, A2 => n266, B1 => 
                           in_buf_25_port, B2 => n242, Z => n395);
   U1372 : AOI22D1 port map( A1 => in_buf_217_port, A2 => n514, B1 => 
                           in_buf_153_port, B2 => n525, Z => n394);
   U1373 : AOI22D1 port map( A1 => in_buf_121_port, A2 => n516, B1 => 
                           in_buf_57_port, B2 => n515, Z => n393);
   U1374 : AOI22D1 port map( A1 => in_buf_249_port, A2 => n534, B1 => 
                           in_buf_185_port, B2 => n531, Z => n392);
   U1375 : NAN4D1 port map( A1 => n395, A2 => n394, A3 => n393, A4 => n392, Z 
                           => N2016);
   U1376 : AOI22D1 port map( A1 => in_buf_90_port, A2 => n266, B1 => 
                           in_buf_26_port, B2 => n242, Z => n399);
   U1377 : AOI22D1 port map( A1 => in_buf_218_port, A2 => n514, B1 => 
                           in_buf_154_port, B2 => n524, Z => n398);
   U1378 : AOI22D1 port map( A1 => in_buf_122_port, A2 => n516, B1 => 
                           in_buf_58_port, B2 => n515, Z => n397);
   U1379 : AOI22D1 port map( A1 => in_buf_250_port, A2 => n518, B1 => 
                           in_buf_186_port, B2 => n532, Z => n396);
   U1380 : NAN4D1 port map( A1 => n399, A2 => n398, A3 => n397, A4 => n396, Z 
                           => N2015);
   U1381 : AOI22D1 port map( A1 => in_buf_91_port, A2 => n266, B1 => 
                           in_buf_27_port, B2 => n242, Z => n403);
   U1382 : AOI22D1 port map( A1 => in_buf_219_port, A2 => n514, B1 => 
                           in_buf_155_port, B2 => n524, Z => n402);
   U1383 : AOI22D1 port map( A1 => in_buf_123_port, A2 => n516, B1 => 
                           in_buf_59_port, B2 => n515, Z => n401);
   U1384 : AOI22D1 port map( A1 => in_buf_251_port, A2 => n518, B1 => 
                           in_buf_187_port, B2 => n532, Z => n400);
   U1385 : NAN4D1 port map( A1 => n403, A2 => n402, A3 => n401, A4 => n400, Z 
                           => N2014);
   U1386 : AOI22D1 port map( A1 => in_buf_92_port, A2 => n266, B1 => 
                           in_buf_28_port, B2 => n242, Z => n407);
   U1387 : AOI22D1 port map( A1 => in_buf_220_port, A2 => n527, B1 => 
                           in_buf_156_port, B2 => n524, Z => n406);
   U1388 : AOI22D1 port map( A1 => in_buf_124_port, A2 => n516, B1 => 
                           in_buf_60_port, B2 => n515, Z => n405);
   U1389 : AOI22D1 port map( A1 => in_buf_252_port, A2 => n518, B1 => 
                           in_buf_188_port, B2 => n532, Z => n404);
   U1390 : NAN4D1 port map( A1 => n407, A2 => n406, A3 => n405, A4 => n404, Z 
                           => N2013);
   U1391 : AOI22D1 port map( A1 => in_buf_93_port, A2 => n266, B1 => 
                           in_buf_29_port, B2 => n242, Z => n411);
   U1392 : AOI22D1 port map( A1 => in_buf_221_port, A2 => n514, B1 => 
                           in_buf_157_port, B2 => n524, Z => n410);
   U1393 : AOI22D1 port map( A1 => in_buf_125_port, A2 => n516, B1 => 
                           in_buf_61_port, B2 => n515, Z => n409);
   U1394 : AOI22D1 port map( A1 => in_buf_253_port, A2 => n518, B1 => 
                           in_buf_189_port, B2 => n532, Z => n408);
   U1395 : NAN4D1 port map( A1 => n411, A2 => n410, A3 => n409, A4 => n408, Z 
                           => N2012);
   U1396 : AOI22D1 port map( A1 => in_buf_94_port, A2 => n266, B1 => 
                           in_buf_30_port, B2 => n242, Z => n415);
   U1397 : AOI22D1 port map( A1 => in_buf_222_port, A2 => n527, B1 => 
                           in_buf_158_port, B2 => n524, Z => n414);
   U1398 : AOI22D1 port map( A1 => in_buf_126_port, A2 => n516, B1 => 
                           in_buf_62_port, B2 => n515, Z => n413);
   U1399 : AOI22D1 port map( A1 => in_buf_254_port, A2 => n534, B1 => 
                           in_buf_190_port, B2 => n532, Z => n412);
   U1400 : NAN4D1 port map( A1 => n415, A2 => n414, A3 => n413, A4 => n412, Z 
                           => N2011);
   U1401 : AOI22D1 port map( A1 => in_buf_95_port, A2 => n266, B1 => 
                           in_buf_31_port, B2 => n242, Z => n419);
   U1402 : AOI22D1 port map( A1 => in_buf_223_port, A2 => n514, B1 => 
                           in_buf_159_port, B2 => n524, Z => n418);
   U1403 : AOI22D1 port map( A1 => in_buf_255_port, A2 => n518, B1 => 
                           in_buf_191_port, B2 => n532, Z => n416);
   U1404 : NAN4D1 port map( A1 => n419, A2 => n418, A3 => n417, A4 => n416, Z 
                           => N2010);
   U1405 : AOI22D1 port map( A1 => comp_res_96_port, A2 => n514, B1 => 
                           comp_res_32_port, B2 => n524, Z => n422);
   U1406 : AOI22D1 port map( A1 => comp_res_128_port, A2 => n518, B1 => 
                           comp_res_64_port, B2 => n532, Z => n420);
   U1407 : AOI22D1 port map( A1 => comp_res_97_port, A2 => n514, B1 => 
                           comp_res_33_port, B2 => n524, Z => n425);
   U1408 : AOI22D1 port map( A1 => comp_res_129_port, A2 => n518, B1 => 
                           comp_res_65_port, B2 => n532, Z => n423);
   U1409 : AOI22D1 port map( A1 => comp_res_98_port, A2 => n514, B1 => 
                           comp_res_34_port, B2 => n524, Z => n428);
   U1410 : AOI22D1 port map( A1 => comp_res_130_port, A2 => n518, B1 => 
                           comp_res_66_port, B2 => n532, Z => n426);
   U1411 : AOI22D1 port map( A1 => comp_res_99_port, A2 => n514, B1 => 
                           comp_res_35_port, B2 => n524, Z => n431);
   U1412 : AOI22D1 port map( A1 => comp_res_131_port, A2 => n518, B1 => 
                           comp_res_67_port, B2 => n532, Z => n429);
   U1413 : AOI22D1 port map( A1 => comp_res_100_port, A2 => n514, B1 => 
                           comp_res_36_port, B2 => n524, Z => n434);
   U1414 : AOI22D1 port map( A1 => comp_res_132_port, A2 => n518, B1 => 
                           comp_res_68_port, B2 => n532, Z => n432);
   U1415 : AOI22D1 port map( A1 => comp_res_101_port, A2 => n514, B1 => 
                           comp_res_37_port, B2 => n524, Z => n437);
   U1416 : AOI22D1 port map( A1 => comp_res_133_port, A2 => n518, B1 => 
                           comp_res_69_port, B2 => n532, Z => n435);
   U1417 : AOI22D1 port map( A1 => comp_res_102_port, A2 => n514, B1 => 
                           comp_res_38_port, B2 => n524, Z => n440);
   U1418 : AOI22D1 port map( A1 => comp_res_134_port, A2 => n518, B1 => 
                           comp_res_70_port, B2 => n532, Z => n438);
   U1419 : AOI22D1 port map( A1 => comp_res_103_port, A2 => n514, B1 => 
                           comp_res_39_port, B2 => n525, Z => n443);
   U1420 : AOI22D1 port map( A1 => comp_res_135_port, A2 => n518, B1 => 
                           comp_res_71_port, B2 => n531, Z => n441);
   U1421 : AOI22D1 port map( A1 => comp_res_104_port, A2 => n514, B1 => 
                           comp_res_40_port, B2 => n513, Z => n446);
   U1422 : AOI22D1 port map( A1 => comp_res_136_port, A2 => n534, B1 => 
                           comp_res_72_port, B2 => n517, Z => n444);
   U1423 : AOI22D1 port map( A1 => comp_res_105_port, A2 => n514, B1 => 
                           comp_res_41_port, B2 => n525, Z => n449);
   U1424 : AOI22D1 port map( A1 => comp_res_137_port, A2 => n518, B1 => 
                           comp_res_73_port, B2 => n517, Z => n447);
   U1425 : AOI22D1 port map( A1 => comp_res_106_port, A2 => n514, B1 => 
                           comp_res_42_port, B2 => n524, Z => n452);
   U1426 : AOI22D1 port map( A1 => comp_res_138_port, A2 => n534, B1 => 
                           comp_res_74_port, B2 => n517, Z => n450);
   U1427 : AOI22D1 port map( A1 => comp_res_107_port, A2 => n527, B1 => 
                           comp_res_43_port, B2 => n513, Z => n455);
   U1428 : AOI22D1 port map( A1 => comp_res_139_port, A2 => n518, B1 => 
                           comp_res_75_port, B2 => n532, Z => n453);
   U1429 : AOI22D1 port map( A1 => comp_res_108_port, A2 => n514, B1 => 
                           comp_res_44_port, B2 => n525, Z => n458);
   U1430 : AOI22D1 port map( A1 => comp_res_140_port, A2 => n534, B1 => 
                           comp_res_76_port, B2 => n517, Z => n456);
   U1431 : AOI22D1 port map( A1 => comp_res_109_port, A2 => n514, B1 => 
                           comp_res_45_port, B2 => n524, Z => n461);
   U1432 : AOI22D1 port map( A1 => comp_res_141_port, A2 => n518, B1 => 
                           comp_res_77_port, B2 => n517, Z => n459);
   U1433 : AOI22D1 port map( A1 => comp_res_110_port, A2 => n514, B1 => 
                           comp_res_46_port, B2 => n513, Z => n464);
   U1434 : AOI22D1 port map( A1 => comp_res_142_port, A2 => n534, B1 => 
                           comp_res_78_port, B2 => n532, Z => n462);
   U1435 : AOI22D1 port map( A1 => comp_res_111_port, A2 => n514, B1 => 
                           comp_res_47_port, B2 => n524, Z => n467);
   U1436 : AOI22D1 port map( A1 => comp_res_143_port, A2 => n518, B1 => 
                           comp_res_79_port, B2 => n531, Z => n465);
   U1437 : AOI22D1 port map( A1 => comp_res_112_port, A2 => n514, B1 => 
                           comp_res_48_port, B2 => n513, Z => n470);
   U1438 : AOI22D1 port map( A1 => comp_res_144_port, A2 => n518, B1 => 
                           comp_res_80_port, B2 => n517, Z => n468);
   U1439 : AOI22D1 port map( A1 => comp_res_113_port, A2 => n514, B1 => 
                           comp_res_49_port, B2 => n513, Z => n473);
   U1440 : AOI22D1 port map( A1 => comp_res_145_port, A2 => n518, B1 => 
                           comp_res_81_port, B2 => n531, Z => n471);
   U1441 : AOI22D1 port map( A1 => comp_res_114_port, A2 => n514, B1 => 
                           comp_res_50_port, B2 => n524, Z => n476);
   U1442 : AOI22D1 port map( A1 => comp_res_146_port, A2 => n534, B1 => 
                           comp_res_82_port, B2 => n531, Z => n474);
   U1443 : AOI22D1 port map( A1 => comp_res_115_port, A2 => n514, B1 => 
                           comp_res_51_port, B2 => n524, Z => n479);
   U1444 : AOI22D1 port map( A1 => comp_res_147_port, A2 => n518, B1 => 
                           comp_res_83_port, B2 => n531, Z => n477);
   U1445 : AOI22D1 port map( A1 => comp_res_116_port, A2 => n514, B1 => 
                           comp_res_52_port, B2 => n513, Z => n482);
   U1446 : AOI22D1 port map( A1 => comp_res_148_port, A2 => n518, B1 => 
                           comp_res_84_port, B2 => n531, Z => n480);
   U1447 : AOI22D1 port map( A1 => comp_res_117_port, A2 => n514, B1 => 
                           comp_res_53_port, B2 => n513, Z => n485);
   U1448 : AOI22D1 port map( A1 => comp_res_149_port, A2 => n518, B1 => 
                           comp_res_85_port, B2 => n531, Z => n483);
   U1449 : AOI22D1 port map( A1 => comp_res_118_port, A2 => n514, B1 => 
                           comp_res_54_port, B2 => n513, Z => n488);
   U1450 : AOI22D1 port map( A1 => comp_res_150_port, A2 => n518, B1 => 
                           comp_res_86_port, B2 => n531, Z => n486);
   U1451 : AOI22D1 port map( A1 => comp_res_119_port, A2 => n527, B1 => 
                           comp_res_55_port, B2 => n513, Z => n491);
   U1452 : AOI22D1 port map( A1 => comp_res_151_port, A2 => n518, B1 => 
                           comp_res_87_port, B2 => n531, Z => n489);
   U1453 : AOI22D1 port map( A1 => comp_res_120_port, A2 => n514, B1 => 
                           comp_res_56_port, B2 => n513, Z => n494);
   U1454 : AOI22D1 port map( A1 => comp_res_152_port, A2 => n518, B1 => 
                           comp_res_88_port, B2 => n531, Z => n492);
   U1455 : AOI22D1 port map( A1 => comp_res_121_port, A2 => n514, B1 => 
                           comp_res_57_port, B2 => n513, Z => n497);
   U1456 : AOI22D1 port map( A1 => comp_res_153_port, A2 => n534, B1 => 
                           comp_res_89_port, B2 => n531, Z => n495);
   U1457 : AOI22D1 port map( A1 => comp_res_122_port, A2 => n514, B1 => 
                           comp_res_58_port, B2 => n513, Z => n500);
   U1458 : AOI22D1 port map( A1 => comp_res_154_port, A2 => n518, B1 => 
                           comp_res_90_port, B2 => n531, Z => n498);
   U1459 : AOI22D1 port map( A1 => comp_res_123_port, A2 => n514, B1 => 
                           comp_res_59_port, B2 => n513, Z => n503);
   U1460 : AOI22D1 port map( A1 => comp_res_155_port, A2 => n518, B1 => 
                           comp_res_91_port, B2 => n531, Z => n501);
   U1461 : AOI22D1 port map( A1 => comp_res_124_port, A2 => n514, B1 => 
                           comp_res_60_port, B2 => n513, Z => n506);
   U1462 : AOI22D1 port map( A1 => comp_res_156_port, A2 => n534, B1 => 
                           comp_res_92_port, B2 => n531, Z => n504);
   U1463 : AOI22D1 port map( A1 => comp_res_125_port, A2 => n514, B1 => 
                           comp_res_61_port, B2 => n513, Z => n509);
   U1464 : AOI22D1 port map( A1 => comp_res_157_port, A2 => n518, B1 => 
                           comp_res_93_port, B2 => n531, Z => n507);
   U1465 : AOI22D1 port map( A1 => comp_res_126_port, A2 => n514, B1 => 
                           comp_res_62_port, B2 => n513, Z => n512);
   U1466 : AOI22D1 port map( A1 => comp_res_158_port, A2 => n534, B1 => 
                           comp_res_94_port, B2 => n531, Z => n510);
   U1467 : AOI22D1 port map( A1 => comp_res_127_port, A2 => n514, B1 => 
                           comp_res_63_port, B2 => n525, Z => n521);
   U1468 : AOI22D1 port map( A1 => comp_res_159_port, A2 => n518, B1 => 
                           comp_res_95_port, B2 => n531, Z => n519);
   U1469 : NOR2D1 port map( A1 => n671, A2 => N63, Z => n535);
   U1470 : NOR2D1 port map( A1 => n671, A2 => n697, Z => n536);
   U1471 : AOI22D1 port map( A1 => out_buf_80_port, A2 => n268, B1 => 
                           out_buf_16_port, B2 => n243, Z => n542);
   U1472 : NOR2D1 port map( A1 => N63, A2 => N64, Z => n537);
   U1473 : NOR2D1 port map( A1 => n697, A2 => N64, Z => n538);
   U1474 : AOI22D1 port map( A1 => out_buf_208_port, A2 => n269, B1 => 
                           out_buf_144_port, B2 => n244, Z => n541);
   U1475 : NOR2M1D1 port map( A1 => n535, A2 => N62, Z => n664);
   U1476 : NOR2M1D1 port map( A1 => n536, A2 => N62, Z => n663);
   U1477 : AOI22D1 port map( A1 => out_buf_112_port, A2 => n664, B1 => 
                           out_buf_48_port, B2 => n663, Z => n540);
   U1478 : NOR2M1D1 port map( A1 => n537, A2 => N62, Z => n666);
   U1479 : NOR2M1D1 port map( A1 => n538, A2 => N62, Z => n665);
   U1480 : AOI22D1 port map( A1 => out_buf_240_port, A2 => n666, B1 => 
                           out_buf_176_port, B2 => n665, Z => n539);
   U1481 : NAN4D1 port map( A1 => n542, A2 => n541, A3 => n540, A4 => n539, Z 
                           => N2882);
   U1482 : AOI22D1 port map( A1 => out_buf_81_port, A2 => n268, B1 => 
                           out_buf_17_port, B2 => n243, Z => n546);
   U1483 : AOI22D1 port map( A1 => out_buf_209_port, A2 => n269, B1 => 
                           out_buf_145_port, B2 => n244, Z => n545);
   U1484 : AOI22D1 port map( A1 => out_buf_113_port, A2 => n664, B1 => 
                           out_buf_49_port, B2 => n663, Z => n544);
   U1485 : AOI22D1 port map( A1 => out_buf_241_port, A2 => n666, B1 => 
                           out_buf_177_port, B2 => n665, Z => n543);
   U1486 : NAN4D1 port map( A1 => n546, A2 => n545, A3 => n544, A4 => n543, Z 
                           => N2881);
   U1487 : AOI22D1 port map( A1 => out_buf_82_port, A2 => n268, B1 => 
                           out_buf_18_port, B2 => n243, Z => n550);
   U1488 : AOI22D1 port map( A1 => out_buf_210_port, A2 => n269, B1 => 
                           out_buf_146_port, B2 => n244, Z => n549);
   U1489 : AOI22D1 port map( A1 => out_buf_114_port, A2 => n664, B1 => 
                           out_buf_50_port, B2 => n663, Z => n548);
   U1490 : AOI22D1 port map( A1 => out_buf_242_port, A2 => n666, B1 => 
                           out_buf_178_port, B2 => n665, Z => n547);
   U1491 : NAN4D1 port map( A1 => n550, A2 => n549, A3 => n548, A4 => n547, Z 
                           => N2880);
   U1492 : AOI22D1 port map( A1 => out_buf_83_port, A2 => n268, B1 => 
                           out_buf_19_port, B2 => n243, Z => n554);
   U1493 : AOI22D1 port map( A1 => out_buf_211_port, A2 => n269, B1 => 
                           out_buf_147_port, B2 => n244, Z => n553);
   U1494 : AOI22D1 port map( A1 => out_buf_115_port, A2 => n664, B1 => 
                           out_buf_51_port, B2 => n663, Z => n552);
   U1495 : AOI22D1 port map( A1 => out_buf_243_port, A2 => n666, B1 => 
                           out_buf_179_port, B2 => n665, Z => n551);
   U1496 : NAN4D1 port map( A1 => n554, A2 => n553, A3 => n552, A4 => n551, Z 
                           => N2879);
   U1497 : AOI22D1 port map( A1 => out_buf_84_port, A2 => n268, B1 => 
                           out_buf_20_port, B2 => n243, Z => n558);
   U1498 : AOI22D1 port map( A1 => out_buf_212_port, A2 => n269, B1 => 
                           out_buf_148_port, B2 => n244, Z => n557);
   U1499 : AOI22D1 port map( A1 => out_buf_116_port, A2 => n664, B1 => 
                           out_buf_52_port, B2 => n663, Z => n556);
   U1500 : AOI22D1 port map( A1 => out_buf_244_port, A2 => n666, B1 => 
                           out_buf_180_port, B2 => n665, Z => n555);
   U1501 : NAN4D1 port map( A1 => n558, A2 => n557, A3 => n556, A4 => n555, Z 
                           => N2878);
   U1502 : AOI22D1 port map( A1 => out_buf_85_port, A2 => n268, B1 => 
                           out_buf_21_port, B2 => n243, Z => n562);
   U1503 : AOI22D1 port map( A1 => out_buf_213_port, A2 => n269, B1 => 
                           out_buf_149_port, B2 => n244, Z => n561);
   U1504 : AOI22D1 port map( A1 => out_buf_117_port, A2 => n664, B1 => 
                           out_buf_53_port, B2 => n663, Z => n560);
   U1505 : AOI22D1 port map( A1 => out_buf_245_port, A2 => n666, B1 => 
                           out_buf_181_port, B2 => n665, Z => n559);
   U1506 : NAN4D1 port map( A1 => n562, A2 => n561, A3 => n560, A4 => n559, Z 
                           => N2877);
   U1507 : AOI22D1 port map( A1 => out_buf_86_port, A2 => n268, B1 => 
                           out_buf_22_port, B2 => n243, Z => n566);
   U1508 : AOI22D1 port map( A1 => out_buf_214_port, A2 => n269, B1 => 
                           out_buf_150_port, B2 => n244, Z => n565);
   U1509 : AOI22D1 port map( A1 => out_buf_118_port, A2 => n664, B1 => 
                           out_buf_54_port, B2 => n663, Z => n564);
   U1510 : AOI22D1 port map( A1 => out_buf_246_port, A2 => n666, B1 => 
                           out_buf_182_port, B2 => n665, Z => n563);
   U1511 : NAN4D1 port map( A1 => n566, A2 => n565, A3 => n564, A4 => n563, Z 
                           => N2876);
   U1512 : AOI22D1 port map( A1 => out_buf_87_port, A2 => n268, B1 => 
                           out_buf_23_port, B2 => n243, Z => n570);
   U1513 : AOI22D1 port map( A1 => out_buf_215_port, A2 => n269, B1 => 
                           out_buf_151_port, B2 => n244, Z => n569);
   U1514 : AOI22D1 port map( A1 => out_buf_119_port, A2 => n664, B1 => 
                           out_buf_55_port, B2 => n663, Z => n568);
   U1515 : AOI22D1 port map( A1 => out_buf_247_port, A2 => n666, B1 => 
                           out_buf_183_port, B2 => n665, Z => n567);
   U1516 : NAN4D1 port map( A1 => n570, A2 => n569, A3 => n568, A4 => n567, Z 
                           => N2875);
   U1517 : AOI22D1 port map( A1 => out_buf_88_port, A2 => n268, B1 => 
                           out_buf_24_port, B2 => n243, Z => n574);
   U1518 : AOI22D1 port map( A1 => out_buf_216_port, A2 => n269, B1 => 
                           out_buf_152_port, B2 => n244, Z => n573);
   U1519 : AOI22D1 port map( A1 => out_buf_120_port, A2 => n664, B1 => 
                           out_buf_56_port, B2 => n663, Z => n572);
   U1520 : AOI22D1 port map( A1 => out_buf_248_port, A2 => n666, B1 => 
                           out_buf_184_port, B2 => n665, Z => n571);
   U1521 : NAN4D1 port map( A1 => n574, A2 => n573, A3 => n572, A4 => n571, Z 
                           => N2874);
   U1522 : AOI22D1 port map( A1 => out_buf_89_port, A2 => n268, B1 => 
                           out_buf_25_port, B2 => n243, Z => n578);
   U1523 : AOI22D1 port map( A1 => out_buf_217_port, A2 => n269, B1 => 
                           out_buf_153_port, B2 => n244, Z => n577);
   U1524 : AOI22D1 port map( A1 => out_buf_121_port, A2 => n664, B1 => 
                           out_buf_57_port, B2 => n663, Z => n576);
   U1525 : AOI22D1 port map( A1 => out_buf_249_port, A2 => n666, B1 => 
                           out_buf_185_port, B2 => n665, Z => n575);
   U1526 : NAN4D1 port map( A1 => n578, A2 => n577, A3 => n576, A4 => n575, Z 
                           => N2873);
   U1527 : AOI22D1 port map( A1 => out_buf_90_port, A2 => n268, B1 => 
                           out_buf_26_port, B2 => n243, Z => n582);
   U1528 : AOI22D1 port map( A1 => out_buf_218_port, A2 => n269, B1 => 
                           out_buf_154_port, B2 => n244, Z => n581);
   U1529 : AOI22D1 port map( A1 => out_buf_122_port, A2 => n664, B1 => 
                           out_buf_58_port, B2 => n663, Z => n580);
   U1530 : AOI22D1 port map( A1 => out_buf_250_port, A2 => n666, B1 => 
                           out_buf_186_port, B2 => n665, Z => n579);
   U1531 : NAN4D1 port map( A1 => n582, A2 => n581, A3 => n580, A4 => n579, Z 
                           => N2872);
   U1532 : AOI22D1 port map( A1 => out_buf_91_port, A2 => n268, B1 => 
                           out_buf_27_port, B2 => n243, Z => n586);
   U1533 : AOI22D1 port map( A1 => out_buf_219_port, A2 => n269, B1 => 
                           out_buf_155_port, B2 => n244, Z => n585);
   U1534 : AOI22D1 port map( A1 => out_buf_123_port, A2 => n664, B1 => 
                           out_buf_59_port, B2 => n663, Z => n584);
   U1535 : AOI22D1 port map( A1 => out_buf_251_port, A2 => n666, B1 => 
                           out_buf_187_port, B2 => n665, Z => n583);
   U1536 : NAN4D1 port map( A1 => n586, A2 => n585, A3 => n584, A4 => n583, Z 
                           => N2871);
   U1537 : AOI22D1 port map( A1 => out_buf_92_port, A2 => n268, B1 => 
                           out_buf_28_port, B2 => n243, Z => n5901);
   U1538 : AOI22D1 port map( A1 => out_buf_220_port, A2 => n269, B1 => 
                           out_buf_156_port, B2 => n244, Z => n589);
   U1539 : AOI22D1 port map( A1 => out_buf_124_port, A2 => n664, B1 => 
                           out_buf_60_port, B2 => n663, Z => n588);
   U1540 : AOI22D1 port map( A1 => out_buf_252_port, A2 => n666, B1 => 
                           out_buf_188_port, B2 => n665, Z => n587);
   U1541 : NAN4D1 port map( A1 => n5901, A2 => n589, A3 => n588, A4 => n587, Z 
                           => N2870);
   U1542 : AOI22D1 port map( A1 => out_buf_93_port, A2 => n268, B1 => 
                           out_buf_29_port, B2 => n243, Z => n594);
   U1543 : AOI22D1 port map( A1 => out_buf_221_port, A2 => n269, B1 => 
                           out_buf_157_port, B2 => n244, Z => n593);
   U1544 : AOI22D1 port map( A1 => out_buf_125_port, A2 => n664, B1 => 
                           out_buf_61_port, B2 => n663, Z => n592);
   U1545 : AOI22D1 port map( A1 => out_buf_253_port, A2 => n666, B1 => 
                           out_buf_189_port, B2 => n665, Z => n591);
   U1546 : NAN4D1 port map( A1 => n594, A2 => n593, A3 => n592, A4 => n591, Z 
                           => N2869);
   U1547 : AOI22D1 port map( A1 => out_buf_94_port, A2 => n268, B1 => 
                           out_buf_30_port, B2 => n243, Z => n598);
   U1548 : AOI22D1 port map( A1 => out_buf_222_port, A2 => n269, B1 => 
                           out_buf_158_port, B2 => n244, Z => n597);
   U1549 : AOI22D1 port map( A1 => out_buf_126_port, A2 => n664, B1 => 
                           out_buf_62_port, B2 => n663, Z => n596);
   U1550 : AOI22D1 port map( A1 => out_buf_254_port, A2 => n666, B1 => 
                           out_buf_190_port, B2 => n665, Z => n595);
   U1551 : NAN4D1 port map( A1 => n598, A2 => n597, A3 => n596, A4 => n595, Z 
                           => N2868);
   U1552 : AOI22D1 port map( A1 => out_buf_95_port, A2 => n268, B1 => 
                           out_buf_31_port, B2 => n243, Z => n602);
   U1553 : AOI22D1 port map( A1 => out_buf_223_port, A2 => n269, B1 => 
                           out_buf_159_port, B2 => n244, Z => n601);
   U1554 : AOI22D1 port map( A1 => out_buf_127_port, A2 => n664, B1 => 
                           out_buf_63_port, B2 => n663, Z => n6001);
   U1555 : AOI22D1 port map( A1 => out_buf_255_port, A2 => n666, B1 => 
                           out_buf_191_port, B2 => n665, Z => n599);
   U1556 : NAN4D1 port map( A1 => n602, A2 => n601, A3 => n6001, A4 => n599, Z 
                           => N2867);
   U1557 : AOI22D1 port map( A1 => out_buf_64_port, A2 => n268, B1 => 
                           out_buf_0_port, B2 => n243, Z => n606);
   U1558 : AOI22D1 port map( A1 => out_buf_192_port, A2 => n269, B1 => 
                           out_buf_128_port, B2 => n244, Z => n605);
   U1559 : AOI22D1 port map( A1 => out_buf_96_port, A2 => n664, B1 => 
                           out_buf_32_port, B2 => n663, Z => n604);
   U1560 : AOI22D1 port map( A1 => out_buf_224_port, A2 => n666, B1 => 
                           out_buf_160_port, B2 => n665, Z => n603);
   U1561 : NAN4D1 port map( A1 => n606, A2 => n605, A3 => n604, A4 => n603, Z 
                           => N2865);
   U1562 : AOI22D1 port map( A1 => out_buf_65_port, A2 => n268, B1 => 
                           out_buf_1_port, B2 => n243, Z => n6101);
   U1563 : AOI22D1 port map( A1 => out_buf_193_port, A2 => n269, B1 => 
                           out_buf_129_port, B2 => n244, Z => n609);
   U1564 : AOI22D1 port map( A1 => out_buf_97_port, A2 => n664, B1 => 
                           out_buf_33_port, B2 => n663, Z => n608);
   U1565 : AOI22D1 port map( A1 => out_buf_225_port, A2 => n666, B1 => 
                           out_buf_161_port, B2 => n665, Z => n607);
   U1566 : NAN4D1 port map( A1 => n6101, A2 => n609, A3 => n608, A4 => n607, Z 
                           => N2864);
   U1567 : AOI22D1 port map( A1 => out_buf_66_port, A2 => n268, B1 => 
                           out_buf_2_port, B2 => n243, Z => n614);
   U1568 : AOI22D1 port map( A1 => out_buf_194_port, A2 => n269, B1 => 
                           out_buf_130_port, B2 => n244, Z => n613);
   U1569 : AOI22D1 port map( A1 => out_buf_98_port, A2 => n664, B1 => 
                           out_buf_34_port, B2 => n663, Z => n612);
   U1570 : AOI22D1 port map( A1 => out_buf_226_port, A2 => n666, B1 => 
                           out_buf_162_port, B2 => n665, Z => n611);
   U1571 : NAN4D1 port map( A1 => n614, A2 => n613, A3 => n612, A4 => n611, Z 
                           => N2863);
   U1572 : AOI22D1 port map( A1 => out_buf_67_port, A2 => n268, B1 => 
                           out_buf_3_port, B2 => n243, Z => n618);
   U1573 : AOI22D1 port map( A1 => out_buf_195_port, A2 => n269, B1 => 
                           out_buf_131_port, B2 => n244, Z => n617);
   U1574 : AOI22D1 port map( A1 => out_buf_99_port, A2 => n664, B1 => 
                           out_buf_35_port, B2 => n663, Z => n616);
   U1575 : AOI22D1 port map( A1 => out_buf_227_port, A2 => n666, B1 => 
                           out_buf_163_port, B2 => n665, Z => n615);
   U1576 : NAN4D1 port map( A1 => n618, A2 => n617, A3 => n616, A4 => n615, Z 
                           => N2862);
   U1577 : AOI22D1 port map( A1 => out_buf_68_port, A2 => n268, B1 => 
                           out_buf_4_port, B2 => n243, Z => n622);
   U1578 : AOI22D1 port map( A1 => out_buf_196_port, A2 => n269, B1 => 
                           out_buf_132_port, B2 => n244, Z => n621);
   U1579 : AOI22D1 port map( A1 => out_buf_100_port, A2 => n664, B1 => 
                           out_buf_36_port, B2 => n663, Z => n620);
   U1580 : AOI22D1 port map( A1 => out_buf_228_port, A2 => n666, B1 => 
                           out_buf_164_port, B2 => n665, Z => n619);
   U1581 : NAN4D1 port map( A1 => n622, A2 => n621, A3 => n620, A4 => n619, Z 
                           => N2861);
   U1582 : AOI22D1 port map( A1 => out_buf_69_port, A2 => n268, B1 => 
                           out_buf_5_port, B2 => n243, Z => n626);
   U1583 : AOI22D1 port map( A1 => out_buf_197_port, A2 => n269, B1 => 
                           out_buf_133_port, B2 => n244, Z => n625);
   U1584 : AOI22D1 port map( A1 => out_buf_101_port, A2 => n664, B1 => 
                           out_buf_37_port, B2 => n663, Z => n624);
   U1585 : AOI22D1 port map( A1 => out_buf_229_port, A2 => n666, B1 => 
                           out_buf_165_port, B2 => n665, Z => n623);
   U1586 : NAN4D1 port map( A1 => n626, A2 => n625, A3 => n624, A4 => n623, Z 
                           => N2860);
   U1587 : AOI22D1 port map( A1 => out_buf_70_port, A2 => n268, B1 => 
                           out_buf_6_port, B2 => n243, Z => n6301);
   U1588 : AOI22D1 port map( A1 => out_buf_198_port, A2 => n269, B1 => 
                           out_buf_134_port, B2 => n244, Z => n629);
   U1589 : AOI22D1 port map( A1 => out_buf_102_port, A2 => n664, B1 => 
                           out_buf_38_port, B2 => n663, Z => n628);
   U1590 : AOI22D1 port map( A1 => out_buf_230_port, A2 => n666, B1 => 
                           out_buf_166_port, B2 => n665, Z => n627);
   U1591 : NAN4D1 port map( A1 => n6301, A2 => n629, A3 => n628, A4 => n627, Z 
                           => N2859);
   U1592 : AOI22D1 port map( A1 => out_buf_71_port, A2 => n268, B1 => 
                           out_buf_7_port, B2 => n243, Z => n634);
   U1593 : AOI22D1 port map( A1 => out_buf_199_port, A2 => n269, B1 => 
                           out_buf_135_port, B2 => n244, Z => n633);
   U1594 : AOI22D1 port map( A1 => out_buf_103_port, A2 => n664, B1 => 
                           out_buf_39_port, B2 => n663, Z => n632);
   U1595 : AOI22D1 port map( A1 => out_buf_231_port, A2 => n666, B1 => 
                           out_buf_167_port, B2 => n665, Z => n631);
   U1596 : NAN4D1 port map( A1 => n634, A2 => n633, A3 => n632, A4 => n631, Z 
                           => N2858);
   U1597 : AOI22D1 port map( A1 => out_buf_72_port, A2 => n268, B1 => 
                           out_buf_8_port, B2 => n243, Z => n638);
   U1598 : AOI22D1 port map( A1 => out_buf_200_port, A2 => n269, B1 => 
                           out_buf_136_port, B2 => n244, Z => n637);
   U1599 : AOI22D1 port map( A1 => out_buf_104_port, A2 => n664, B1 => 
                           out_buf_40_port, B2 => n663, Z => n636);
   U1600 : AOI22D1 port map( A1 => out_buf_232_port, A2 => n666, B1 => 
                           out_buf_168_port, B2 => n665, Z => n635);
   U1601 : NAN4D1 port map( A1 => n638, A2 => n637, A3 => n636, A4 => n635, Z 
                           => N2857);
   U1602 : AOI22D1 port map( A1 => out_buf_73_port, A2 => n268, B1 => 
                           out_buf_9_port, B2 => n243, Z => n642);
   U1603 : AOI22D1 port map( A1 => out_buf_201_port, A2 => n269, B1 => 
                           out_buf_137_port, B2 => n244, Z => n641);
   U1604 : AOI22D1 port map( A1 => out_buf_105_port, A2 => n664, B1 => 
                           out_buf_41_port, B2 => n663, Z => n6401);
   U1605 : AOI22D1 port map( A1 => out_buf_233_port, A2 => n666, B1 => 
                           out_buf_169_port, B2 => n665, Z => n639);
   U1606 : NAN4D1 port map( A1 => n642, A2 => n641, A3 => n6401, A4 => n639, Z 
                           => N2856);
   U1607 : AOI22D1 port map( A1 => out_buf_74_port, A2 => n268, B1 => 
                           out_buf_10_port, B2 => n243, Z => n646);
   U1608 : AOI22D1 port map( A1 => out_buf_202_port, A2 => n269, B1 => 
                           out_buf_138_port, B2 => n244, Z => n645);
   U1609 : AOI22D1 port map( A1 => out_buf_106_port, A2 => n664, B1 => 
                           out_buf_42_port, B2 => n663, Z => n644);
   U1610 : AOI22D1 port map( A1 => out_buf_234_port, A2 => n666, B1 => 
                           out_buf_170_port, B2 => n665, Z => n643);
   U1611 : NAN4D1 port map( A1 => n646, A2 => n645, A3 => n644, A4 => n643, Z 
                           => N2855);
   U1612 : AOI22D1 port map( A1 => out_buf_75_port, A2 => n268, B1 => 
                           out_buf_11_port, B2 => n243, Z => n650);
   U1613 : AOI22D1 port map( A1 => out_buf_203_port, A2 => n269, B1 => 
                           out_buf_139_port, B2 => n244, Z => n649);
   U1614 : AOI22D1 port map( A1 => out_buf_107_port, A2 => n664, B1 => 
                           out_buf_43_port, B2 => n663, Z => n648);
   U1615 : AOI22D1 port map( A1 => out_buf_235_port, A2 => n666, B1 => 
                           out_buf_171_port, B2 => n665, Z => n647);
   U1616 : NAN4D1 port map( A1 => n650, A2 => n649, A3 => n648, A4 => n647, Z 
                           => N2854);
   U1617 : AOI22D1 port map( A1 => out_buf_76_port, A2 => n268, B1 => 
                           out_buf_12_port, B2 => n243, Z => n654);
   U1618 : AOI22D1 port map( A1 => out_buf_204_port, A2 => n269, B1 => 
                           out_buf_140_port, B2 => n244, Z => n653);
   U1619 : AOI22D1 port map( A1 => out_buf_108_port, A2 => n664, B1 => 
                           out_buf_44_port, B2 => n663, Z => n652);
   U1620 : AOI22D1 port map( A1 => out_buf_236_port, A2 => n666, B1 => 
                           out_buf_172_port, B2 => n665, Z => n651);
   U1621 : NAN4D1 port map( A1 => n654, A2 => n653, A3 => n652, A4 => n651, Z 
                           => N2853);
   U1622 : AOI22D1 port map( A1 => out_buf_77_port, A2 => n268, B1 => 
                           out_buf_13_port, B2 => n243, Z => n658);
   U1623 : AOI22D1 port map( A1 => out_buf_205_port, A2 => n269, B1 => 
                           out_buf_141_port, B2 => n244, Z => n657);
   U1624 : AOI22D1 port map( A1 => out_buf_109_port, A2 => n664, B1 => 
                           out_buf_45_port, B2 => n663, Z => n656);
   U1625 : AOI22D1 port map( A1 => out_buf_237_port, A2 => n666, B1 => 
                           out_buf_173_port, B2 => n665, Z => n655);
   U1626 : NAN4D1 port map( A1 => n658, A2 => n657, A3 => n656, A4 => n655, Z 
                           => N2852);
   U1627 : AOI22D1 port map( A1 => out_buf_78_port, A2 => n268, B1 => 
                           out_buf_14_port, B2 => n243, Z => n662);
   U1628 : AOI22D1 port map( A1 => out_buf_206_port, A2 => n269, B1 => 
                           out_buf_142_port, B2 => n244, Z => n661);
   U1629 : AOI22D1 port map( A1 => out_buf_110_port, A2 => n664, B1 => 
                           out_buf_46_port, B2 => n663, Z => n660);
   U1630 : AOI22D1 port map( A1 => out_buf_238_port, A2 => n666, B1 => 
                           out_buf_174_port, B2 => n665, Z => n659);
   U1631 : NAN4D1 port map( A1 => n662, A2 => n661, A3 => n660, A4 => n659, Z 
                           => N2851);
   U1632 : AOI22D1 port map( A1 => out_buf_79_port, A2 => n268, B1 => 
                           out_buf_15_port, B2 => n243, Z => n670);
   U1633 : AOI22D1 port map( A1 => out_buf_207_port, A2 => n269, B1 => 
                           out_buf_143_port, B2 => n244, Z => n669);
   U1634 : AOI22D1 port map( A1 => out_buf_111_port, A2 => n664, B1 => 
                           out_buf_47_port, B2 => n663, Z => n668);
   U1635 : AOI22D1 port map( A1 => out_buf_239_port, A2 => n666, B1 => 
                           out_buf_175_port, B2 => n665, Z => n667);
   U1636 : NAN4D1 port map( A1 => n670, A2 => n669, A3 => n668, A4 => n667, Z 
                           => N2850);
   U1637 : NOR3D1 port map( A1 => avs_addr(3), A2 => avs_addr(5), A3 => 
                           avs_addr(4), Z => N66);

end hier_filter_none_20;
