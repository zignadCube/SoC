
library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

package CONV_PACK_siso_gen is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_siso_gen;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_siso_gen.all;

architecture flat_gcd_16_1p5 of siso_gen is

   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFDL
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVDL
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M10DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22DL
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M20DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component TIELO
      port( Z : out std_logic);
   end component;
   
   component NAN4D1
      port( A1, A2, A3, A4 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN4DL
      port( A1, A2, A3, A4 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22M10DL
      port( B1, B2, A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22M10D1
      port( B1, B2, A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AO21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22M20DL
      port( B1, B2, A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN4M2D1
      port( A1, A2, A3, A4 : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFRPQ1
      port( D, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFRPB1
      port( D, CK, RB : in std_logic;  Q, QB : out std_logic);
   end component;
   
   component DFFRPQL
      port( D, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFSPQ1
      port( D, CK, SB : in std_logic;  Q : out std_logic);
   end component;
   
   signal req_port, data_out_15_port, data_out_14_port, data_out_13_port, 
      data_out_12_port, data_out_11_port, data_out_10_port, data_out_9_port, 
      data_out_8_port, data_out_7_port, data_out_6_port, data_out_5_port, 
      data_out_4_port, data_out_3_port, data_out_2_port, data_out_1_port, 
      data_out_0_port, num2_15_port, num2_14_port, num2_13_port, num2_12_port, 
      num2_11_port, num2_10_port, num2_9_port, num2_8_port, num2_7_port, 
      num2_6_port, num2_5_port, num2_4_port, num2_2_port, num2_0_port, odd, 
      sub_res_15, sub_res_14, sub_res_13, sub_res_12, sub_res_11, sub_res_10, 
      sub_res_9, sub_res_8, sub_res_7, sub_res_6, sub_res_5, sub_res_4, 
      sub_res_3, sub_res_2, sub_res_1, sub_res_0, N82, N83, N84, N85, N86, N87,
      N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, n1, n56, n57, n58, n59,
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n820, n830, n840, n850, n860, n870, 
      n880, n890, N810, N800, N790, N780, N770, N760, N750, N740, N730, N720, 
      N710, N700, N690, N680, N670, N660, n900, n910, n920, n930, n940, n950, 
      n960, n970, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n170, n171, n172, n173, n174, n175, n176, n_1003, sub_63_n224
      , sub_63_n223, sub_63_n222, sub_63_n221, sub_63_n220, sub_63_n219, 
      sub_63_n218, sub_63_n217, sub_63_n216, sub_63_n215, sub_63_n214, 
      sub_63_n213, sub_63_n212, sub_63_n211, sub_63_n210, sub_63_n209, 
      sub_63_n208, sub_63_n207, sub_63_n206, sub_63_n205, sub_63_n204, 
      sub_63_n203, sub_63_n202, sub_63_n146, sub_63_n145, sub_63_n144, 
      sub_63_n143, sub_63_n142, sub_63_n141, sub_63_n140, sub_63_n139, 
      sub_63_n138, sub_63_n137, sub_63_n136, sub_63_n135, sub_63_n134, 
      sub_63_n133, sub_63_n132, sub_63_n131, sub_63_n125, sub_63_n122, 
      sub_63_n121, sub_63_n120, sub_63_n119, sub_63_n118, sub_63_n115, 
      sub_63_n114, sub_63_n113, sub_63_n112, sub_63_n111, sub_63_n110, 
      sub_63_n109, sub_63_n108, sub_63_n107, sub_63_n106, sub_63_n105, 
      sub_63_n104, sub_63_n103, sub_63_n102, sub_63_n101, sub_63_n100, 
      sub_63_n99, sub_63_n98, sub_63_n97, sub_63_n96, sub_63_n90, sub_63_n89, 
      sub_63_n88, sub_63_n87, sub_63_n84, sub_63_n83, sub_63_n82, sub_63_n81, 
      sub_63_n80, sub_63_n79, sub_63_n78, sub_63_n77, sub_63_n76, sub_63_n75, 
      sub_63_n73, sub_63_n72, sub_63_n70, sub_63_n69, sub_63_n68, sub_63_n67, 
      sub_63_n62, sub_63_n61, sub_63_n60, sub_63_n59, sub_63_n56, sub_63_n55, 
      sub_63_n54, sub_63_n53, sub_63_n52, sub_63_n51, sub_63_n50, sub_63_n49, 
      sub_63_n48, sub_63_n47, sub_63_n45, sub_63_n42, sub_63_n41, sub_63_n40, 
      sub_63_n39, sub_63_n38, sub_63_n37, sub_63_n36, sub_63_n35, sub_63_n34, 
      sub_63_n33, sub_63_n32, sub_63_n31, sub_63_n30, sub_63_n29, sub_63_n25, 
      sub_63_n24, sub_63_n23, sub_63_n22, sub_63_n21, sub_63_n20, sub_63_n18, 
      sub_63_n17, sub_63_n16, sub_63_n15, sub_63_n14, sub_63_n12, sub_63_n11, 
      sub_63_n6, sub_63_n4, sub_63_n3, sub_63_n2, sub_63_n1, 
      add_0_root_add_80_ni_n89, add_0_root_add_80_ni_n88, 
      add_0_root_add_80_ni_n51, add_0_root_add_80_ni_n50, 
      add_0_root_add_80_ni_n47, add_0_root_add_80_ni_n46, 
      add_0_root_add_80_ni_n45, add_0_root_add_80_ni_n44, 
      add_0_root_add_80_ni_n43, add_0_root_add_80_ni_n42, 
      add_0_root_add_80_ni_n41, add_0_root_add_80_ni_n40, 
      add_0_root_add_80_ni_n39, add_0_root_add_80_ni_n38, 
      add_0_root_add_80_ni_n37, add_0_root_add_80_ni_n35, 
      add_0_root_add_80_ni_n34, add_0_root_add_80_ni_n33, 
      add_0_root_add_80_ni_n32, add_0_root_add_80_ni_n29, 
      add_0_root_add_80_ni_n28, add_0_root_add_80_ni_n27, 
      add_0_root_add_80_ni_n26, add_0_root_add_80_ni_n23, 
      add_0_root_add_80_ni_n19, add_0_root_add_80_ni_n18, 
      add_0_root_add_80_ni_n17, add_0_root_add_80_ni_n14, 
      add_0_root_add_80_ni_n13, add_0_root_add_80_ni_n10, 
      add_0_root_add_80_ni_n9, add_0_root_add_80_ni_n8, add_0_root_add_80_ni_n7
      , add_0_root_add_80_ni_n6, add_0_root_add_80_ni_n3, 
      add_0_root_add_80_ni_n1 : std_logic;

begin
   req <= req_port;
   data_out <= ( data_out_15_port, data_out_14_port, data_out_13_port, 
      data_out_12_port, data_out_11_port, data_out_10_port, data_out_9_port, 
      data_out_8_port, data_out_7_port, data_out_6_port, data_out_5_port, 
      data_out_4_port, data_out_3_port, data_out_2_port, data_out_1_port, 
      data_out_0_port );
   
   req_i_reg : DFFSPQ1 port map( D => n890, CK => clk, SB => n175, Q => 
                           req_port);
   odd_reg : DFFRPQ1 port map( D => n880, CK => clk, RB => n175, Q => odd);
   num2_reg_15 : DFFRPQ1 port map( D => n56, CK => clk, RB => n175, Q => 
                           num2_15_port);
   num1_reg_14 : DFFRPQ1 port map( D => n73, CK => clk, RB => n175, Q => 
                           data_out_14_port);
   num2_reg_14 : DFFRPQ1 port map( D => n57, CK => clk, RB => n175, Q => 
                           num2_14_port);
   num1_reg_12 : DFFRPQ1 port map( D => n75, CK => clk, RB => n175, Q => 
                           data_out_12_port);
   num2_reg_12 : DFFRPQ1 port map( D => n59, CK => clk, RB => n175, Q => 
                           num2_12_port);
   num1_reg_13 : DFFRPQ1 port map( D => n74, CK => clk, RB => n175, Q => 
                           data_out_13_port);
   num2_reg_13 : DFFRPQ1 port map( D => n58, CK => clk, RB => n175, Q => 
                           num2_13_port);
   num1_reg_4 : DFFRPQ1 port map( D => n830, CK => clk, RB => n175, Q => 
                           data_out_4_port);
   num2_reg_4 : DFFRPQ1 port map( D => n67, CK => clk, RB => n175, Q => 
                           num2_4_port);
   num1_reg_10 : DFFRPQ1 port map( D => n77, CK => clk, RB => n175, Q => 
                           data_out_10_port);
   num1_reg_8 : DFFRPQ1 port map( D => n79, CK => clk, RB => n175, Q => 
                           data_out_8_port);
   num1_reg_6 : DFFRPQ1 port map( D => n81, CK => clk, RB => n175, Q => 
                           data_out_6_port);
   num2_reg_8 : DFFRPQ1 port map( D => n63, CK => clk, RB => n175, Q => 
                           num2_8_port);
   num1_reg_2 : DFFRPQ1 port map( D => n850, CK => clk, RB => n175, Q => 
                           data_out_2_port);
   num2_reg_6 : DFFRPQ1 port map( D => n65, CK => clk, RB => n175, Q => 
                           num2_6_port);
   num1_reg_9 : DFFRPQ1 port map( D => n78, CK => clk, RB => n175, Q => 
                           data_out_9_port);
   num2_reg_10 : DFFRPQ1 port map( D => n61, CK => clk, RB => n175, Q => 
                           num2_10_port);
   num1_reg_11 : DFFRPQ1 port map( D => n76, CK => clk, RB => n175, Q => 
                           data_out_11_port);
   num2_reg_2 : DFFRPQ1 port map( D => n69, CK => clk, RB => n175, Q => 
                           num2_2_port);
   num1_reg_3 : DFFRPQ1 port map( D => n840, CK => clk, RB => n175, Q => 
                           data_out_3_port);
   num1_reg_7 : DFFRPQ1 port map( D => n80, CK => clk, RB => n175, Q => 
                           data_out_7_port);
   num1_reg_5 : DFFRPQ1 port map( D => n820, CK => clk, RB => n175, Q => 
                           data_out_5_port);
   num1_reg_0 : DFFRPQ1 port map( D => n870, CK => clk, RB => n175, Q => 
                           data_out_0_port);
   num2_reg_9 : DFFRPQ1 port map( D => n62, CK => clk, RB => n175, Q => 
                           num2_9_port);
   num2_reg_5 : DFFRPQ1 port map( D => n66, CK => clk, RB => n175, Q => 
                           num2_5_port);
   num2_reg_11 : DFFRPQ1 port map( D => n60, CK => clk, RB => n175, Q => 
                           num2_11_port);
   num2_reg_0 : DFFRPQ1 port map( D => n71, CK => clk, RB => n175, Q => 
                           num2_0_port);
   num2_reg_7 : DFFRPQ1 port map( D => n64, CK => clk, RB => n175, Q => 
                           num2_7_port);
   ready_reg : DFFRPQ1 port map( D => n176, CK => clk, RB => n175, Q => ready);
   num1_reg_15 : DFFRPQL port map( D => n72, CK => clk, RB => n175, Q => 
                           data_out_15_port);
   num2_reg_1 : DFFRPB1 port map( D => n70, CK => clk, RB => n175, Q => n98, QB
                           => n970);
   num2_reg_3 : DFFRPQ1 port map( D => n68, CK => clk, RB => n175, Q => n104);
   num1_reg_1 : DFFRPQ1 port map( D => n860, CK => clk, RB => n175, Q => 
                           data_out_1_port);
   U87 : NAN4M2D1 port map( A1 => sub_res_9, A2 => sub_res_8, A3 => N700, A4 =>
                           N710, Z => n115);
   U88 : INVD2 port map( A => sub_res_15, Z => N660);
   U89 : INVD1 port map( A => n173, Z => n119);
   U90 : INVD1 port map( A => sub_res_6, Z => N750);
   U91 : OAI21D1 port map( A1 => sub_res_15, A2 => n138, B => n110, Z => n169);
   U92 : OAI22M20DL port map( B1 => n140, B2 => n137, A1 => n910, A2 => 
                           data_out_15_port, Z => n72);
   U93 : OAI21DL port map( A1 => n148, A2 => n137, B => n124, Z => n76);
   U94 : OAI21DL port map( A1 => n160, A2 => n137, B => n129, Z => n820);
   U95 : OAI21DL port map( A1 => n150, A2 => n110, B => n125, Z => n77);
   U96 : OAI21DL port map( A1 => n146, A2 => n111, B => n123, Z => n75);
   U97 : OAI21DL port map( A1 => n142, A2 => n137, B => n121, Z => n73);
   U98 : OAI21DL port map( A1 => n144, A2 => n110, B => n122, Z => n74);
   U99 : OAI21DL port map( A1 => n152, A2 => n111, B => n126, Z => n78);
   U100 : OAI21DL port map( A1 => n154, A2 => n137, B => n127, Z => n79);
   U101 : OAI21DL port map( A1 => n162, A2 => n110, B => n130, Z => n830);
   U102 : OAI21DL port map( A1 => n166, A2 => n137, B => n132, Z => n850);
   U103 : INVD1 port map( A => sub_res_11, Z => N700);
   U104 : INVD1 port map( A => sub_res_10, Z => N710);
   U105 : INVD1 port map( A => sub_res_12, Z => N690);
   U106 : INVD1 port map( A => sub_res_13, Z => N680);
   U107 : INVD1 port map( A => n110, Z => n920);
   U108 : NAN2D1 port map( A1 => n120, A2 => n172, Z => n900);
   U109 : NAN2D1 port map( A1 => n120, A2 => n172, Z => n910);
   U110 : NAN2D1 port map( A1 => n120, A2 => n172, Z => n134);
   U111 : NAN2D1 port map( A1 => data_out_7_port, A2 => n134, Z => n101);
   U112 : AO21D1 port map( A1 => data_in(7), A2 => n920, B => n930, Z => n80);
   U113 : NAN2D1 port map( A1 => n100, A2 => n101, Z => n930);
   U114 : OR2D1 port map( A1 => n172, A2 => n148, Z => n940);
   U115 : NAN2D1 port map( A1 => n940, A2 => n147, Z => n60);
   U116 : AOI22D1 port map( A1 => num2_11_port, A2 => n169, B1 => N93, B2 => 
                           n107, Z => n147);
   U117 : INVDL port map( A => sub_res_8, Z => N730);
   U118 : OAI21M20D1 port map( A1 => n138, A2 => data_in(14), B => n141, Z => 
                           n57);
   U119 : NAN2D1 port map( A1 => N96, A2 => n107, Z => n950);
   U120 : INVD1 port map( A => num2_15_port, Z => n103);
   U121 : NAN2DL port map( A1 => num2_14_port, A2 => n169, Z => n960);
   U122 : AND2D1 port map( A1 => n950, A2 => n960, Z => n141);
   U123 : INVD1 port map( A => n970, Z => n99);
   U124 : NAN4DL port map( A1 => N760, A2 => N770, A3 => N740, A4 => N750, Z =>
                           n114);
   U125 : NAN2D1 port map( A1 => odd, A2 => req_port, Z => n172);
   U126 : NAN2DL port map( A1 => n106, A2 => sub_res_7, Z => n100);
   U127 : OR2D1 port map( A1 => n172, A2 => n140, Z => n102);
   U128 : NAN2D1 port map( A1 => n102, A2 => n139, Z => n56);
   U129 : AOI22M10D1 port map( B1 => N97, B2 => n107, A1 => n103, A2 => n169, Z
                           => n139);
   U130 : AOI22DL port map( A1 => num2_10_port, A2 => n169, B1 => N92, B2 => 
                           n107, Z => n149);
   U131 : INVD1 port map( A => num2_12_port, Z => n105);
   U132 : AOI22M10DL port map( B1 => N94, B2 => n107, A1 => n105, A2 => n169, Z
                           => n145);
   U133 : AOI22M10DL port map( B1 => data_out_6_port, B2 => n900, A1 => N750, 
                           A2 => n106, Z => n128);
   U134 : AOI22M10DL port map( B1 => data_out_1_port, B2 => n910, A1 => N800, 
                           A2 => n106, Z => n133);
   U135 : AOI22DL port map( A1 => n106, A2 => sub_res_2, B1 => data_out_2_port,
                           B2 => n910, Z => n132);
   U136 : AOI22DL port map( A1 => n106, A2 => sub_res_5, B1 => data_out_5_port,
                           B2 => n910, Z => n129);
   U137 : AOI22DL port map( A1 => n106, A2 => sub_res_8, B1 => data_out_8_port,
                           B2 => n900, Z => n127);
   U138 : AOI22DL port map( A1 => n106, A2 => sub_res_11, B1 => 
                           data_out_11_port, B2 => n900, Z => n124);
   U139 : AOI22DL port map( A1 => n106, A2 => sub_res_14, B1 => 
                           data_out_14_port, B2 => n900, Z => n121);
   U140 : AOI22DL port map( A1 => n106, A2 => sub_res_3, B1 => data_out_3_port,
                           B2 => n134, Z => n131);
   U141 : AOI22DL port map( A1 => n106, A2 => n109, B1 => data_out_9_port, B2 
                           => n910, Z => n126);
   U142 : AOI22DL port map( A1 => n106, A2 => sub_res_12, B1 => 
                           data_out_12_port, B2 => n910, Z => n123);
   U143 : AOI22DL port map( A1 => n106, A2 => sub_res_4, B1 => data_out_4_port,
                           B2 => n900, Z => n130);
   U144 : AOI22DL port map( A1 => n106, A2 => sub_res_10, B1 => 
                           data_out_10_port, B2 => n900, Z => n125);
   U145 : AOI22DL port map( A1 => n106, A2 => sub_res_13, B1 => 
                           data_out_13_port, B2 => n910, Z => n122);
   U146 : NAN4DL port map( A1 => N800, A2 => N810, A3 => N780, A4 => N790, Z =>
                           n113);
   U147 : AOI22DL port map( A1 => n106, A2 => sub_res_0, B1 => data_out_0_port,
                           B2 => n900, Z => n135);
   U148 : AOI22DL port map( A1 => n99, A2 => n169, B1 => N83, B2 => n107, Z => 
                           n167);
   U149 : NAN2D1 port map( A1 => n117, A2 => n118, Z => n173);
   U150 : NOR2D1 port map( A1 => n114, A2 => n113, Z => n118);
   U151 : NOR2D1 port map( A1 => n116, A2 => n115, Z => n117);
   U152 : NAN4D1 port map( A1 => N680, A2 => N690, A3 => N660, A4 => N670, Z =>
                           n116);
   U153 : INVD1 port map( A => sub_res_7, Z => N740);
   U154 : INVD1 port map( A => sub_res_5, Z => N760);
   U155 : INVD1 port map( A => sub_res_2, Z => N790);
   U156 : INVD1 port map( A => sub_res_4, Z => N770);
   U157 : INVD1 port map( A => sub_res_3, Z => N780);
   U158 : AND2D1 port map( A1 => n136, A2 => N660, Z => n106);
   U159 : INVD1 port map( A => n174, Z => n136);
   U160 : INVD1 port map( A => sub_res_14, Z => N670);
   U161 : AND2DL port map( A1 => n136, A2 => sub_res_15, Z => n107);
   U162 : INVD1 port map( A => sub_res_0, Z => N810);
   U163 : INVD1 port map( A => n172, Z => n138);
   U164 : AOI22DL port map( A1 => n169, A2 => num2_0_port, B1 => N82, B2 => 
                           n107, Z => n170);
   U165 : INVD1 port map( A => odd, Z => n112);
   U166 : INVD1 port map( A => data_in(15), Z => n140);
   U167 : INVD1 port map( A => data_in(3), Z => n164);
   U168 : INVD1 port map( A => data_in(1), Z => n168);
   U169 : INVD1 port map( A => data_in(2), Z => n166);
   U170 : INVD1 port map( A => data_in(4), Z => n162);
   U171 : INVD1 port map( A => data_in(5), Z => n160);
   U172 : INVD1 port map( A => data_in(6), Z => n158);
   U173 : INVD1 port map( A => data_in(7), Z => n156);
   U174 : INVD1 port map( A => data_in(8), Z => n154);
   U175 : INVD1 port map( A => data_in(9), Z => n152);
   U176 : INVD1 port map( A => data_in(10), Z => n150);
   U177 : INVD1 port map( A => data_in(11), Z => n148);
   U178 : INVD1 port map( A => data_in(12), Z => n146);
   U179 : INVD1 port map( A => data_in(13), Z => n144);
   U180 : INVD1 port map( A => data_in(14), Z => n142);
   U181 : INVD1 port map( A => reset, Z => n175);
   U182 : TIELO port map( Z => n1);
   U183 : INVDL port map( A => sub_res_9, Z => N720);
   U184 : INVDL port map( A => n119, Z => n108);
   U185 : INVD1 port map( A => sub_res_1, Z => N800);
   U186 : AOI22DL port map( A1 => num2_2_port, A2 => n169, B1 => N84, B2 => 
                           n107, Z => n165);
   U187 : AOI22DL port map( A1 => num2_4_port, A2 => n169, B1 => N86, B2 => 
                           n107, Z => n161);
   U188 : AOI22DL port map( A1 => num2_6_port, A2 => n169, B1 => N88, B2 => 
                           n107, Z => n157);
   U189 : AOI22DL port map( A1 => num2_7_port, A2 => n169, B1 => N89, B2 => 
                           n107, Z => n155);
   U190 : AOI22DL port map( A1 => num2_8_port, A2 => n169, B1 => N90, B2 => 
                           n107, Z => n153);
   U191 : OAI21M20DL port map( A1 => data_in(0), A2 => n920, B => n135, Z => 
                           n870);
   U192 : INVD1 port map( A => data_in(0), Z => n171);
   U193 : AOI22DL port map( A1 => n104, A2 => n169, B1 => N85, B2 => n107, Z =>
                           n163);
   U194 : AOI22DL port map( A1 => num2_5_port, A2 => n169, B1 => N87, B2 => 
                           n107, Z => n159);
   U195 : INVDL port map( A => N720, Z => n109);
   U196 : NAN2D1 port map( A1 => req_port, A2 => n112, Z => n110);
   U197 : NAN2D1 port map( A1 => req_port, A2 => n112, Z => n111);
   U198 : NAN2D1 port map( A1 => req_port, A2 => n112, Z => n137);
   U199 : OAI21D1 port map( A1 => n138, A2 => n112, B => n110, Z => n880);
   U200 : OAI21D1 port map( A1 => n138, A2 => n108, B => n111, Z => n890);
   U201 : OAI21D1 port map( A1 => n119, A2 => sub_res_15, B => n137, Z => n120)
                           ;
   U202 : NAN2D1 port map( A1 => n172, A2 => n111, Z => n174);
   U203 : OAI21D1 port map( A1 => n158, A2 => n111, B => n128, Z => n81);
   U204 : OAI21D1 port map( A1 => n164, A2 => n111, B => n131, Z => n840);
   U205 : OAI21D1 port map( A1 => n168, A2 => n110, B => n133, Z => n860);
   U206 : AOI22D1 port map( A1 => N95, A2 => n107, B1 => num2_13_port, B2 => 
                           n169, Z => n143);
   U207 : OAI21D1 port map( A1 => n172, A2 => n144, B => n143, Z => n58);
   U208 : OAI21D1 port map( A1 => n172, A2 => n146, B => n145, Z => n59);
   U209 : OAI21D1 port map( A1 => n172, A2 => n150, B => n149, Z => n61);
   U210 : AOI22D1 port map( A1 => num2_9_port, A2 => n169, B1 => N91, B2 => 
                           n107, Z => n151);
   U211 : OAI21D1 port map( A1 => n172, A2 => n152, B => n151, Z => n62);
   U212 : OAI21D1 port map( A1 => n172, A2 => n154, B => n153, Z => n63);
   U213 : OAI21D1 port map( A1 => n172, A2 => n156, B => n155, Z => n64);
   U214 : OAI21D1 port map( A1 => n172, A2 => n158, B => n157, Z => n65);
   U215 : OAI21D1 port map( A1 => n172, A2 => n160, B => n159, Z => n66);
   U216 : OAI21D1 port map( A1 => n172, A2 => n162, B => n161, Z => n67);
   U217 : OAI21D1 port map( A1 => n172, A2 => n164, B => n163, Z => n68);
   U218 : OAI21D1 port map( A1 => n172, A2 => n166, B => n165, Z => n69);
   U219 : OAI21D1 port map( A1 => n172, A2 => n168, B => n167, Z => n70);
   U220 : OAI21D1 port map( A1 => n172, A2 => n171, B => n170, Z => n71);
   U221 : NOR2D1 port map( A1 => n174, A2 => n108, Z => n176);
   sub_63_U292 : AOI21DL port map( A1 => sub_63_n1, A2 => sub_63_n31, B => 
                           sub_63_n32, Z => sub_63_n30);
   sub_63_U291 : AOI21DL port map( A1 => sub_63_n1, A2 => sub_63_n40, B => 
                           sub_63_n41, Z => sub_63_n39);
   sub_63_U290 : EXNOR2DL port map( A1 => sub_63_n211, A2 => sub_63_n11, Z => 
                           sub_res_8);
   sub_63_U289 : EXOR2D2 port map( A1 => sub_63_n21, A2 => sub_63_n4, Z => 
                           sub_res_15);
   sub_63_U288 : NAN2D1 port map( A1 => sub_63_n145, A2 => data_out_1_port, Z 
                           => sub_63_n114);
   sub_63_U287 : NAN2DL port map( A1 => sub_63_n215, A2 => sub_63_n114, Z => 
                           sub_63_n18);
   sub_63_U286 : AOI21DL port map( A1 => sub_63_n1, A2 => sub_63_n70, B => 
                           sub_63_n224, Z => sub_63_n69);
   sub_63_U285 : EXOR2DL port map( A1 => sub_63_n18, A2 => sub_63_n222, Z => 
                           sub_res_1);
   sub_63_U284 : EXNOR2DL port map( A1 => sub_63_n216, A2 => data_out_0_port, Z
                           => sub_res_0);
   sub_63_U283 : OAI21DL port map( A1 => sub_63_n2, A2 => sub_63_n33, B => 
                           sub_63_n34, Z => sub_63_n32);
   sub_63_U282 : OAI21DL port map( A1 => sub_63_n2, A2 => sub_63_n42, B => 
                           sub_63_n45, Z => sub_63_n41);
   sub_63_U281 : INVDL port map( A => sub_63_n2, Z => sub_63_n48);
   sub_63_U280 : NOR2D1 port map( A1 => sub_63_n106, A2 => sub_63_n109, Z => 
                           sub_63_n104);
   sub_63_U279 : AND2D1 port map( A1 => sub_63_n209, A2 => sub_63_n29, Z => 
                           sub_63_n223);
   sub_63_U278 : EXNOR2D1 port map( A1 => sub_63_n223, A2 => sub_63_n30, Z => 
                           sub_res_14);
   sub_63_U277 : NOR2DL port map( A1 => sub_63_n216, A2 => data_out_0_port, Z 
                           => sub_63_n222);
   sub_63_U276 : AND2D1 port map( A1 => sub_63_n122, A2 => sub_63_n68, Z => 
                           sub_63_n221);
   sub_63_U275 : EXNOR2D1 port map( A1 => sub_63_n221, A2 => sub_63_n69, Z => 
                           sub_res_9);
   sub_63_U274 : OAI21DL port map( A1 => sub_63_n111, A2 => sub_63_n217, B => 
                           sub_63_n110, Z => sub_63_n108);
   sub_63_U273 : INVDL port map( A => sub_63_n112, Z => sub_63_n111);
   sub_63_U272 : NAN2D1 port map( A1 => sub_63_n142, A2 => data_out_4_port, Z 
                           => sub_63_n101);
   sub_63_U271 : NAN2DL port map( A1 => sub_63_n142, A2 => data_out_4_port, Z 
                           => sub_63_n220);
   sub_63_U270 : NOR2D1 port map( A1 => sub_63_n141, A2 => data_out_5_port, Z 
                           => sub_63_n218);
   sub_63_U269 : NOR2D1 port map( A1 => sub_63_n144, A2 => data_out_2_port, Z 
                           => sub_63_n109);
   sub_63_U268 : NOR2DL port map( A1 => sub_63_n144, A2 => data_out_2_port, Z 
                           => sub_63_n217);
   sub_63_U267 : BUFDL port map( A => sub_63_n146, Z => sub_63_n216);
   sub_63_U266 : OR2DL port map( A1 => sub_63_n145, A2 => data_out_1_port, Z =>
                           sub_63_n215);
   sub_63_U265 : OAI21DL port map( A1 => sub_63_n67, A2 => sub_63_n73, B => 
                           sub_63_n68, Z => sub_63_n214);
   sub_63_U264 : INVD1 port map( A => sub_63_n103, Z => sub_63_n102);
   sub_63_U263 : NOR2D1 port map( A1 => sub_63_n141, A2 => data_out_5_port, Z 
                           => sub_63_n219);
   sub_63_U262 : OAI21DL port map( A1 => sub_63_n219, A2 => sub_63_n101, B => 
                           sub_63_n96, Z => sub_63_n213);
   sub_63_U261 : INVD1 port map( A => sub_63_n84, Z => sub_63_n125);
   sub_63_U260 : OAI21D1 port map( A1 => sub_63_n206, A2 => sub_63_n75, B => 
                           sub_63_n76, Z => sub_63_n212);
   sub_63_U259 : BUFDL port map( A => sub_63_n212, Z => sub_63_n211);
   sub_63_U258 : NOR2D1 port map( A1 => sub_63_n56, A2 => sub_63_n51, Z => 
                           sub_63_n49);
   sub_63_U257 : OR2D1 port map( A1 => sub_63_n131, A2 => data_out_15_port, Z 
                           => sub_63_n210);
   sub_63_U256 : INVD1 port map( A => num2_15_port, Z => sub_63_n131);
   sub_63_U255 : NAN2D1 port map( A1 => sub_63_n132, A2 => data_out_14_port, Z 
                           => sub_63_n29);
   sub_63_U254 : OR2D1 port map( A1 => sub_63_n132, A2 => data_out_14_port, Z 
                           => sub_63_n209);
   sub_63_U253 : INVD1 port map( A => num2_14_port, Z => sub_63_n132);
   sub_63_U252 : NAN2D1 port map( A1 => sub_63_n137, A2 => data_out_9_port, Z 
                           => sub_63_n68);
   sub_63_U251 : NOR2D1 port map( A1 => sub_63_n138, A2 => data_out_8_port, Z 
                           => sub_63_n72);
   sub_63_U250 : NAN2D1 port map( A1 => sub_63_n140, A2 => data_out_6_port, Z 
                           => sub_63_n87);
   sub_63_U249 : NOR2D1 port map( A1 => sub_63_n134, A2 => data_out_12_port, Z 
                           => sub_63_n42);
   sub_63_U248 : NAN2D1 port map( A1 => sub_63_n141, A2 => data_out_5_port, Z 
                           => sub_63_n96);
   sub_63_U247 : NOR2D1 port map( A1 => sub_63_n133, A2 => data_out_13_port, Z 
                           => sub_63_n37);
   sub_63_U246 : NOR2D1 port map( A1 => sub_63_n142, A2 => data_out_4_port, Z 
                           => sub_63_n100);
   sub_63_U245 : NAN2D1 port map( A1 => sub_63_n138, A2 => data_out_8_port, Z 
                           => sub_63_n73);
   sub_63_U244 : INVD1 port map( A => num2_6_port, Z => sub_63_n140);
   sub_63_U243 : NAN2D1 port map( A1 => sub_63_n144, A2 => data_out_2_port, Z 
                           => sub_63_n110);
   sub_63_U242 : NOR2D1 port map( A1 => sub_63_n143, A2 => data_out_3_port, Z 
                           => sub_63_n106);
   sub_63_U241 : INVDL port map( A => num2_11_port, Z => sub_63_n135);
   sub_63_U240 : NAN2D1 port map( A1 => sub_63_n131, A2 => data_out_15_port, Z 
                           => sub_63_n20);
   sub_63_U239 : NAN2D1 port map( A1 => sub_63_n210, A2 => sub_63_n20, Z => 
                           sub_63_n4);
   sub_63_U238 : NOR2D1 port map( A1 => sub_63_n146, A2 => data_out_0_port, Z 
                           => sub_63_n115);
   sub_63_U237 : NOR2D1 port map( A1 => sub_63_n202, A2 => data_out_1_port, Z 
                           => sub_63_n113);
   sub_63_U236 : INVD1 port map( A => num2_7_port, Z => sub_63_n139);
   sub_63_U235 : INVD1 port map( A => sub_63_n220, Z => sub_63_n99);
   sub_63_U234 : NAN2D1 port map( A1 => sub_63_n98, A2 => sub_63_n220, Z => 
                           sub_63_n15);
   sub_63_U233 : NAN2D1 port map( A1 => sub_63_n35, A2 => sub_63_n209, Z => 
                           sub_63_n24);
   sub_63_U232 : NOR2D1 port map( A1 => sub_63_n42, A2 => sub_63_n37, Z => 
                           sub_63_n35);
   sub_63_U231 : NAN2D1 port map( A1 => sub_63_n89, A2 => sub_63_n77, Z => 
                           sub_63_n75);
   sub_63_U230 : NOR2D1 port map( A1 => sub_63_n72, A2 => sub_63_n67, Z => 
                           sub_63_n61);
   sub_63_U229 : AND2D1 port map( A1 => sub_63_n119, A2 => sub_63_n45, Z => 
                           sub_63_n208);
   sub_63_U228 : AOI21DL port map( A1 => sub_63_n212, A2 => sub_63_n47, B => 
                           sub_63_n48, Z => sub_63_n207);
   sub_63_U227 : EXNOR2D1 port map( A1 => sub_63_n207, A2 => sub_63_n208, Z => 
                           sub_res_12);
   sub_63_U226 : NAN2D1 port map( A1 => sub_63_n118, A2 => sub_63_n38, Z => 
                           sub_63_n6);
   sub_63_U225 : OA21M20D1 port map( A1 => sub_63_n36, A2 => sub_63_n209, B => 
                           sub_63_n29, Z => sub_63_n25);
   sub_63_U224 : NOR2D1 port map( A1 => sub_63_n84, A2 => sub_63_n79, Z => 
                           sub_63_n77);
   sub_63_U223 : NOR2D1 port map( A1 => sub_63_n3, A2 => sub_63_n24, Z => 
                           sub_63_n22);
   sub_63_U222 : NAN2D1 port map( A1 => sub_63_n61, A2 => sub_63_n49, Z => 
                           sub_63_n3);
   sub_63_U221 : NAN2DL port map( A1 => sub_63_n133, A2 => data_out_13_port, Z 
                           => sub_63_n38);
   sub_63_U220 : NAN2DL port map( A1 => sub_63_n135, A2 => data_out_11_port, Z 
                           => sub_63_n52);
   sub_63_U219 : NAN2DL port map( A1 => sub_63_n139, A2 => data_out_7_port, Z 
                           => sub_63_n80);
   sub_63_U218 : NAN2DL port map( A1 => sub_63_n136, A2 => data_out_10_port, Z 
                           => sub_63_n59);
   sub_63_U217 : INVDL port map( A => num2_13_port, Z => sub_63_n133);
   sub_63_U216 : INVDL port map( A => num2_12_port, Z => sub_63_n134);
   sub_63_U215 : NAN2DL port map( A1 => sub_63_n143, A2 => data_out_3_port, Z 
                           => sub_63_n107);
   sub_63_U214 : INVDL port map( A => sub_63_n37, Z => sub_63_n118);
   sub_63_U213 : INVDL port map( A => sub_63_n51, Z => sub_63_n120);
   sub_63_U212 : INVDL port map( A => sub_63_n42, Z => sub_63_n119);
   sub_63_U211 : INVDL port map( A => sub_63_n73, Z => sub_63_n224);
   sub_63_U210 : INVDL port map( A => sub_63_n72, Z => sub_63_n70);
   sub_63_U209 : INVDL port map( A => sub_63_n100, Z => sub_63_n98);
   sub_63_U208 : NAN2M1DL port map( A1 => sub_63_n106, A2 => sub_63_n107, Z => 
                           sub_63_n16);
   sub_63_U207 : NAN2M1DL port map( A1 => sub_63_n217, A2 => sub_63_n110, Z => 
                           sub_63_n17);
   sub_63_U206 : NOR2M1DL port map( A1 => sub_63_n89, A2 => sub_63_n84, Z => 
                           sub_63_n82);
   sub_63_U205 : OAI21M10DL port map( A1 => sub_63_n213, A2 => sub_63_n84, B =>
                           sub_63_n87, Z => sub_63_n83);
   sub_63_U204 : EXNOR2D1 port map( A1 => sub_63_n60, A2 => sub_63_n205, Z => 
                           sub_res_10);
   sub_63_U203 : NOR2DL port map( A1 => sub_63_n3, A2 => sub_63_n42, Z => 
                           sub_63_n40);
   sub_63_U202 : NAN2DL port map( A1 => sub_63_n70, A2 => sub_63_n73, Z => 
                           sub_63_n11);
   sub_63_U201 : AND2D1 port map( A1 => sub_63_n120, A2 => sub_63_n52, Z => 
                           sub_63_n204);
   sub_63_U200 : EXNOR2D1 port map( A1 => sub_63_n53, A2 => sub_63_n204, Z => 
                           sub_res_11);
   sub_63_U199 : INVDL port map( A => sub_63_n67, Z => sub_63_n122);
   sub_63_U198 : AND2DL port map( A1 => sub_63_n125, A2 => sub_63_n87, Z => 
                           sub_63_n203);
   sub_63_U197 : NAN2M1DL port map( A1 => sub_63_n218, A2 => sub_63_n96, Z => 
                           sub_63_n14);
   sub_63_U196 : NAN2M1DL port map( A1 => sub_63_n79, A2 => sub_63_n80, Z => 
                           sub_63_n12);
   sub_63_U195 : INVDL port map( A => sub_63_n35, Z => sub_63_n33);
   sub_63_U194 : INVDL port map( A => sub_63_n36, Z => sub_63_n34);
   sub_63_U193 : INVDL port map( A => sub_63_n3, Z => sub_63_n47);
   sub_63_U192 : NOR2DL port map( A1 => sub_63_n3, A2 => sub_63_n33, Z => 
                           sub_63_n31);
   sub_63_U191 : NOR2D1 port map( A1 => sub_63_n136, A2 => data_out_10_port, Z 
                           => sub_63_n56);
   sub_63_U190 : INVD1 port map( A => num2_8_port, Z => sub_63_n138);
   sub_63_U189 : NAN2D1 port map( A1 => sub_63_n134, A2 => data_out_12_port, Z 
                           => sub_63_n45);
   sub_63_U188 : INVD1 port map( A => num2_9_port, Z => sub_63_n137);
   sub_63_U187 : INVD1 port map( A => num2_10_port, Z => sub_63_n136);
   sub_63_U186 : AND2DL port map( A1 => sub_63_n121, A2 => sub_63_n59, Z => 
                           sub_63_n205);
   sub_63_U185 : INVD1 port map( A => num2_4_port, Z => sub_63_n142);
   sub_63_U184 : INVDL port map( A => num2_2_port, Z => sub_63_n144);
   sub_63_U183 : INVDL port map( A => n104, Z => sub_63_n143);
   sub_63_U182 : INVDL port map( A => num2_0_port, Z => sub_63_n146);
   sub_63_U181 : INVDL port map( A => n98, Z => sub_63_n145);
   sub_63_U180 : AOI21DL port map( A1 => sub_63_n104, A2 => sub_63_n112, B => 
                           sub_63_n105, Z => sub_63_n206);
   sub_63_U179 : OAI21D1 port map( A1 => sub_63_n75, A2 => sub_63_n103, B => 
                           sub_63_n76, Z => sub_63_n1);
   sub_63_U178 : INVDL port map( A => n98, Z => sub_63_n202);
   sub_63_U177 : AOI21DL port map( A1 => sub_63_n102, A2 => sub_63_n89, B => 
                           sub_63_n213, Z => sub_63_n88);
   sub_63_U176 : EXNOR2DL port map( A1 => sub_63_n102, A2 => sub_63_n15, Z => 
                           sub_res_4);
   sub_63_U175 : NOR2M1DL port map( A1 => sub_63_n61, A2 => sub_63_n56, Z => 
                           sub_63_n54);
   sub_63_U174 : OAI21M10DL port map( A1 => sub_63_n214, A2 => sub_63_n56, B =>
                           sub_63_n59, Z => sub_63_n55);
   sub_63_U173 : INVDL port map( A => sub_63_n56, Z => sub_63_n121);
   sub_63_U172 : OAI21D1 port map( A1 => sub_63_n2, A2 => sub_63_n24, B => 
                           sub_63_n25, Z => sub_63_n23);
   sub_63_U171 : NOR2D1 port map( A1 => sub_63_n135, A2 => data_out_11_port, Z 
                           => sub_63_n51);
   sub_63_U170 : NOR2D1 port map( A1 => sub_63_n139, A2 => data_out_7_port, Z 
                           => sub_63_n79);
   sub_63_U169 : NOR2D1 port map( A1 => sub_63_n137, A2 => data_out_9_port, Z 
                           => sub_63_n67);
   sub_63_U168 : INVD1 port map( A => num2_5_port, Z => sub_63_n141);
   sub_63_U167 : NOR2D1 port map( A1 => sub_63_n100, A2 => sub_63_n218, Z => 
                           sub_63_n89);
   sub_63_U166 : EXNOR2DL port map( A1 => sub_63_n88, A2 => sub_63_n203, Z => 
                           sub_res_6);
   sub_63_U140 : OAI21D1 port map( A1 => sub_63_n115, A2 => sub_63_n113, B => 
                           sub_63_n114, Z => sub_63_n112);
   sub_63_U132 : EXOR2D1 port map( A1 => sub_63_n111, A2 => sub_63_n17, Z => 
                           sub_res_2);
   sub_63_U127 : OAI21D1 port map( A1 => sub_63_n106, A2 => sub_63_n110, B => 
                           sub_63_n107, Z => sub_63_n105);
   sub_63_U125 : AOI21D1 port map( A1 => sub_63_n104, A2 => sub_63_n112, B => 
                           sub_63_n105, Z => sub_63_n103);
   sub_63_U123 : EXNOR2D1 port map( A1 => sub_63_n108, A2 => sub_63_n16, Z => 
                           sub_res_3);
   sub_63_U116 : AOI21D1 port map( A1 => sub_63_n102, A2 => sub_63_n98, B => 
                           sub_63_n99, Z => sub_63_n97);
   sub_63_U110 : OAI21D1 port map( A1 => sub_63_n219, A2 => sub_63_n101, B => 
                           sub_63_n96, Z => sub_63_n90);
   sub_63_U103 : EXOR2D1 port map( A1 => sub_63_n97, A2 => sub_63_n14, Z => 
                           sub_res_5);
   sub_63_U101 : NOR2D2 port map( A1 => sub_63_n140, A2 => data_out_6_port, Z 
                           => sub_63_n84);
   sub_63_U94 : AOI21D1 port map( A1 => sub_63_n102, A2 => sub_63_n82, B => 
                           sub_63_n83, Z => sub_63_n81);
   sub_63_U88 : OAI21D1 port map( A1 => sub_63_n79, A2 => sub_63_n87, B => 
                           sub_63_n80, Z => sub_63_n78);
   sub_63_U86 : AOI21D1 port map( A1 => sub_63_n77, A2 => sub_63_n90, B => 
                           sub_63_n78, Z => sub_63_n76);
   sub_63_U83 : EXOR2D1 port map( A1 => sub_63_n81, A2 => sub_63_n12, Z => 
                           sub_res_7);
   sub_63_U70 : OAI21D1 port map( A1 => sub_63_n67, A2 => sub_63_n73, B => 
                           sub_63_n68, Z => sub_63_n62);
   sub_63_U64 : AOI21D1 port map( A1 => sub_63_n212, A2 => sub_63_n61, B => 
                           sub_63_n214, Z => sub_63_n60);
   sub_63_U54 : AOI21D1 port map( A1 => sub_63_n212, A2 => sub_63_n54, B => 
                           sub_63_n55, Z => sub_63_n53);
   sub_63_U48 : OAI21D1 port map( A1 => sub_63_n51, A2 => sub_63_n59, B => 
                           sub_63_n52, Z => sub_63_n50);
   sub_63_U46 : AOI21D1 port map( A1 => sub_63_n49, A2 => sub_63_n62, B => 
                           sub_63_n50, Z => sub_63_n2);
   sub_63_U26 : OAI21D1 port map( A1 => sub_63_n37, A2 => sub_63_n45, B => 
                           sub_63_n38, Z => sub_63_n36);
   sub_63_U19 : EXOR2D1 port map( A1 => sub_63_n6, A2 => sub_63_n39, Z => 
                           sub_res_13);
   sub_63_U8 : AOI21D1 port map( A1 => sub_63_n1, A2 => sub_63_n22, B => 
                           sub_63_n23, Z => sub_63_n21);
   add_0_root_add_80_ni_U114 : NAN2DL port map( A1 => N700, A2 => N690, Z => 
                           add_0_root_add_80_ni_n10);
   add_0_root_add_80_ni_U113 : NAN2DL port map( A1 => add_0_root_add_80_ni_n19,
                           A2 => N700, Z => add_0_root_add_80_ni_n14);
   add_0_root_add_80_ni_U112 : INVDL port map( A => N720, Z => 
                           add_0_root_add_80_ni_n26);
   add_0_root_add_80_ni_U111 : NAN2D1 port map( A1 => N720, A2 => N710, Z => 
                           add_0_root_add_80_ni_n18);
   add_0_root_add_80_ni_U110 : INVDL port map( A => N670, Z => 
                           add_0_root_add_80_ni_n6);
   add_0_root_add_80_ni_U109 : NOR2D1 port map( A1 => add_0_root_add_80_ni_n27,
                           A2 => add_0_root_add_80_ni_n26, Z => 
                           add_0_root_add_80_ni_n23);
   add_0_root_add_80_ni_U108 : EXOR2D1 port map( A1 => add_0_root_add_80_ni_n3,
                           A2 => N660, Z => N97);
   add_0_root_add_80_ni_U107 : INVD1 port map( A => N810, Z => N82);
   add_0_root_add_80_ni_U106 : INVD1 port map( A => N680, Z => 
                           add_0_root_add_80_ni_n8);
   add_0_root_add_80_ni_U105 : NOR2D1 port map( A1 => add_0_root_add_80_ni_n51,
                           A2 => N82, Z => add_0_root_add_80_ni_n50);
   add_0_root_add_80_ni_U104 : INVD1 port map( A => N750, Z => 
                           add_0_root_add_80_ni_n37);
   add_0_root_add_80_ni_U103 : NOR2D1 port map( A1 => add_0_root_add_80_ni_n18,
                           A2 => add_0_root_add_80_ni_n10, Z => 
                           add_0_root_add_80_ni_n9);
   add_0_root_add_80_ni_U102 : NAN2D1 port map( A1 => add_0_root_add_80_ni_n9, 
                           A2 => add_0_root_add_80_ni_n28, Z => 
                           add_0_root_add_80_ni_n1);
   add_0_root_add_80_ni_U101 : NOR2D1 port map( A1 => add_0_root_add_80_ni_n14,
                           A2 => add_0_root_add_80_ni_n27, Z => 
                           add_0_root_add_80_ni_n13);
   add_0_root_add_80_ni_U100 : NAN2D1 port map( A1 => N730, A2 => 
                           add_0_root_add_80_ni_n33, Z => 
                           add_0_root_add_80_ni_n29);
   add_0_root_add_80_ni_U99 : INVD1 port map( A => N780, Z => 
                           add_0_root_add_80_ni_n46);
   add_0_root_add_80_ni_U98 : INVD1 port map( A => N770, Z => 
                           add_0_root_add_80_ni_n43);
   add_0_root_add_80_ni_U97 : NAN2D1 port map( A1 => N790, A2 => 
                           add_0_root_add_80_ni_n50, Z => 
                           add_0_root_add_80_ni_n47);
   add_0_root_add_80_ni_U96 : NOR2D1 port map( A1 => add_0_root_add_80_ni_n18, 
                           A2 => add_0_root_add_80_ni_n27, Z => 
                           add_0_root_add_80_ni_n17);
   add_0_root_add_80_ni_U95 : NOR2D1 port map( A1 => add_0_root_add_80_ni_n1, 
                           A2 => add_0_root_add_80_ni_n88, Z => 
                           add_0_root_add_80_ni_n3);
   add_0_root_add_80_ni_U94 : NOR2D1 port map( A1 => add_0_root_add_80_ni_n46, 
                           A2 => add_0_root_add_80_ni_n47, Z => 
                           add_0_root_add_80_ni_n45);
   add_0_root_add_80_ni_U93 : EXOR2DL port map( A1 => add_0_root_add_80_ni_n51,
                           A2 => N82, Z => N83);
   add_0_root_add_80_ni_U92 : EXNOR2DL port map( A1 => add_0_root_add_80_ni_n32
                           , A2 => N730, Z => N90);
   add_0_root_add_80_ni_U91 : EXOR2DL port map( A1 => add_0_root_add_80_ni_n35,
                           A2 => add_0_root_add_80_ni_n34, Z => N89);
   add_0_root_add_80_ni_U90 : NAN2DL port map( A1 => add_0_root_add_80_ni_n38, 
                           A2 => N750, Z => add_0_root_add_80_ni_n35);
   add_0_root_add_80_ni_U89 : EXNOR2DL port map( A1 => add_0_root_add_80_ni_n41
                           , A2 => add_0_root_add_80_ni_n42, Z => N87);
   add_0_root_add_80_ni_U88 : NOR2DL port map( A1 => add_0_root_add_80_ni_n43, 
                           A2 => add_0_root_add_80_ni_n44, Z => 
                           add_0_root_add_80_ni_n42);
   add_0_root_add_80_ni_U87 : EXOR2DL port map( A1 => N790, A2 => 
                           add_0_root_add_80_ni_n50, Z => N84);
   add_0_root_add_80_ni_U86 : INVDL port map( A => N800, Z => 
                           add_0_root_add_80_ni_n51);
   add_0_root_add_80_ni_U85 : INVDL port map( A => add_0_root_add_80_ni_n18, Z 
                           => add_0_root_add_80_ni_n19);
   add_0_root_add_80_ni_U84 : INVDL port map( A => N760, Z => 
                           add_0_root_add_80_ni_n41);
   add_0_root_add_80_ni_U83 : INVDL port map( A => N740, Z => 
                           add_0_root_add_80_ni_n34);
   add_0_root_add_80_ni_U82 : NAN2DL port map( A1 => add_0_root_add_80_ni_n38, 
                           A2 => add_0_root_add_80_ni_n33, Z => 
                           add_0_root_add_80_ni_n32);
   add_0_root_add_80_ni_U81 : INVDL port map( A => add_0_root_add_80_ni_n45, Z 
                           => add_0_root_add_80_ni_n44);
   add_0_root_add_80_ni_U80 : INVDL port map( A => add_0_root_add_80_ni_n39, Z 
                           => add_0_root_add_80_ni_n38);
   add_0_root_add_80_ni_U79 : EXOR2DL port map( A1 => add_0_root_add_80_ni_n13,
                           A2 => N690, Z => N94);
   add_0_root_add_80_ni_U78 : EXOR2DL port map( A1 => add_0_root_add_80_ni_n23,
                           A2 => N710, Z => N92);
   add_0_root_add_80_ni_U77 : INVD2 port map( A => add_0_root_add_80_ni_n28, Z 
                           => add_0_root_add_80_ni_n27);
   add_0_root_add_80_ni_U76 : BUFDL port map( A => add_0_root_add_80_ni_n27, Z 
                           => add_0_root_add_80_ni_n89);
   add_0_root_add_80_ni_U75 : NOR2D1 port map( A1 => add_0_root_add_80_ni_n1, 
                           A2 => add_0_root_add_80_ni_n8, Z => 
                           add_0_root_add_80_ni_n7);
   add_0_root_add_80_ni_U74 : EXOR2D1 port map( A1 => add_0_root_add_80_ni_n17,
                           A2 => N700, Z => N93);
   add_0_root_add_80_ni_U73 : AND2D1 port map( A1 => N750, A2 => N740, Z => 
                           add_0_root_add_80_ni_n33);
   add_0_root_add_80_ni_U72 : NOR2D2 port map( A1 => add_0_root_add_80_ni_n41, 
                           A2 => add_0_root_add_80_ni_n43, Z => 
                           add_0_root_add_80_ni_n40);
   add_0_root_add_80_ni_U71 : NAN2D2 port map( A1 => add_0_root_add_80_ni_n40, 
                           A2 => add_0_root_add_80_ni_n45, Z => 
                           add_0_root_add_80_ni_n39);
   add_0_root_add_80_ni_U70 : OR2D1 port map( A1 => add_0_root_add_80_ni_n8, A2
                           => add_0_root_add_80_ni_n6, Z => 
                           add_0_root_add_80_ni_n88);
   add_0_root_add_80_ni_U56 : EXOR2D1 port map( A1 => add_0_root_add_80_ni_n46,
                           A2 => add_0_root_add_80_ni_n47, Z => N85);
   add_0_root_add_80_ni_U53 : EXOR2D1 port map( A1 => add_0_root_add_80_ni_n43,
                           A2 => add_0_root_add_80_ni_n44, Z => N86);
   add_0_root_add_80_ni_U44 : EXNOR2D1 port map( A1 => add_0_root_add_80_ni_n38
                           , A2 => add_0_root_add_80_ni_n37, Z => N88);
   add_0_root_add_80_ni_U36 : NOR2D2 port map( A1 => add_0_root_add_80_ni_n29, 
                           A2 => add_0_root_add_80_ni_n39, Z => 
                           add_0_root_add_80_ni_n28);
   add_0_root_add_80_ni_U29 : EXOR2D1 port map( A1 => add_0_root_add_80_ni_n89,
                           A2 => add_0_root_add_80_ni_n26, Z => N91);
   add_0_root_add_80_ni_U8 : EXOR2D1 port map( A1 => add_0_root_add_80_ni_n8, 
                           A2 => add_0_root_add_80_ni_n1, Z => N95);
   add_0_root_add_80_ni_U3 : EXNOR2D1 port map( A1 => add_0_root_add_80_ni_n7, 
                           A2 => add_0_root_add_80_ni_n6, Z => N96);

end flat_gcd_16_1p5;
