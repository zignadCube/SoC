
library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

package CONV_PACK_siso_gen is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_siso_gen;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_siso_gen.all;

architecture flat_sec_par_16_5 of siso_gen is

   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component ADHALFD1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AO21D2
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22D2
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVBD32
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22DL
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVDL
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component ADFULD2
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI22M10D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR3D4
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFDL
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AO21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR3D2
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFD2
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component NAN2M1DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21M10D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFD2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN3D2
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M10D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN3M1D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D4
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component ADFULDL
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component EXOR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR3DL
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFD4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AO21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21M10DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OA22DL
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21M20DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22D4
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22M10D1
      port( B1, B2, A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVBD2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21M20DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M20DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AO21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M10DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD16
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD20
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M20D2
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AO21M10DL
      port( A2, A1, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN3M1DL
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D4
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFD20
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AO21M20DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OA22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component TIELO
      port( Z : out std_logic);
   end component;
   
   component TIEHI
      port( Z : out std_logic);
   end component;
   
   component BUFD8
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INVBD4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFERPQ1
      port( D, CEB, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component DFERPQ4
      port( D, CEB, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component DFERPQL
      port( D, CEB, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component DFERPQ2
      port( D, CEB, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFRPQ1
      port( D, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   signal ready_port, coeff_memory_79_port, coeff_memory_78_port, 
      coeff_memory_77_port, coeff_memory_76_port, coeff_memory_75_port, 
      coeff_memory_74_port, coeff_memory_73_port, coeff_memory_72_port, 
      coeff_memory_71_port, coeff_memory_70_port, coeff_memory_69_port, 
      coeff_memory_68_port, coeff_memory_67_port, coeff_memory_66_port, 
      coeff_memory_65_port, coeff_memory_64_port, coeff_memory_63_port, 
      coeff_memory_62_port, coeff_memory_61_port, coeff_memory_60_port, 
      coeff_memory_59_port, coeff_memory_58_port, coeff_memory_57_port, 
      coeff_memory_56_port, coeff_memory_55_port, coeff_memory_54_port, 
      coeff_memory_53_port, coeff_memory_52_port, coeff_memory_51_port, 
      coeff_memory_50_port, coeff_memory_49_port, coeff_memory_48_port, 
      coeff_memory_47_port, coeff_memory_46_port, coeff_memory_45_port, 
      coeff_memory_44_port, coeff_memory_43_port, coeff_memory_42_port, 
      coeff_memory_41_port, coeff_memory_40_port, coeff_memory_39_port, 
      coeff_memory_38_port, coeff_memory_37_port, coeff_memory_36_port, 
      coeff_memory_35_port, coeff_memory_34_port, coeff_memory_33_port, 
      coeff_memory_32_port, coeff_memory_31_port, coeff_memory_30_port, 
      coeff_memory_29_port, coeff_memory_28_port, coeff_memory_27_port, 
      coeff_memory_26_port, coeff_memory_25_port, coeff_memory_24_port, 
      coeff_memory_23_port, coeff_memory_22_port, coeff_memory_21_port, 
      coeff_memory_20_port, coeff_memory_19_port, coeff_memory_18_port, 
      coeff_memory_17_port, coeff_memory_16_port, coeff_memory_15_port, 
      coeff_memory_14_port, coeff_memory_13_port, coeff_memory_12_port, 
      coeff_memory_11_port, coeff_memory_10_port, coeff_memory_9_port, 
      coeff_memory_8_port, coeff_memory_7_port, coeff_memory_6_port, 
      coeff_memory_5_port, coeff_memory_4_port, coeff_memory_3_port, 
      coeff_memory_2_port, coeff_memory_1_port, coeff_memory_0_port, 
      coeff_counter_2_port, coeff_counter_1_port, coeff_counter_0_port, 
      z1_15_port, z1_14_port, z1_13_port, z1_12_port, z1_11_port, z1_10_port, 
      z1_9_port, z1_8_port, z1_7_port, z1_6_port, z1_5_port, z1_4_port, 
      z1_3_port, z1_2_port, z1_1_port, z1_0_port, z2_15_port, z2_14_port, 
      z2_13_port, z2_12_port, z2_11_port, z2_10_port, z2_9_port, z2_8_port, 
      z2_7_port, z2_6_port, z2_5_port, z2_4_port, z2_3_port, z2_2_port, 
      z2_1_port, z2_0_port, z1_next_15_port, z1_next_14_port, z1_next_13_port, 
      z1_next_12_port, z1_next_11_port, z1_next_10_port, z1_next_9_port, 
      z1_next_8_port, z1_next_7_port, z1_next_6_port, z1_next_5_port, 
      z1_next_4_port, z1_next_3_port, z1_next_2_port, z1_next_1_port, 
      z1_next_0_port, z2_next_15_port, z2_next_14_port, z2_next_13_port, 
      z2_next_12_port, z2_next_11_port, z2_next_10_port, z2_next_9_port, 
      z2_next_8_port, z2_next_7_port, z2_next_6_port, z2_next_5_port, 
      z2_next_4_port, z2_next_3_port, z2_next_2_port, z2_next_1_port, 
      z2_next_0_port, y_15_port, y_14_port, y_13_port, y_12_port, y_11_port, 
      y_10_port, y_9_port, y_8_port, y_7_port, y_6_port, y_5_port, y_4_port, 
      y_3_port, y_2_port, y_1_port, y_0_port, n22, n23, n25, n26, n27, n28, n29
      , n30, n31, n32, z2_temp_9, z2_temp_8, z2_temp_7, z2_temp_6, z2_temp_5, 
      z2_temp_4, z2_temp_3, z2_temp_2, z2_temp_1, z2_temp_15, z2_temp_14, 
      z2_temp_13, z2_temp_12, z2_temp_11, z2_temp_10, z2_temp_0, m3_9, m3_8, 
      m3_7, m3_6, m3_5, m3_4, m3_3, m3_2, m3_1, m3_15, m3_14, m3_13, m3_12, 
      m3_11, m3_10, m3_0, m2_9, m2_8, m2_7, m2_6, m2_5, m2_4, m2_3, m2_2, m2_1,
      m2_15, m2_14, m2_13, m2_12, m2_11, m2_10, m2_0, m5_9, m5_8, m5_7, m5_6, 
      m5_5, m5_4, m5_3, m5_2, m5_1, m5_15, m5_14, m5_13, m5_12, m5_11, m5_10, 
      m5_0, m4_9, m4_8, m4_7, m4_6, m4_5, m4_4, m4_3, m4_2, m4_1, m4_15, m4_14,
      m4_13, m4_12, m4_11, m4_10, m4_0, m1_9, m1_8, m1_7, m1_6, m1_5, m1_4, 
      m1_3, m1_2, m1_1, m1_15, m1_14, m1_13, m1_12, m1_11, m1_10, m1_0, n33, 
      n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48
      , n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n_1091
      , n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100,
      n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, 
      n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, 
      n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, 
      n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, 
      n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, 
      n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, 
      n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, 
      n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, 
      n_1173, n_1174, mult_28_C94_n940, mult_28_C94_n939, mult_28_C94_n938, 
      mult_28_C94_n937, mult_28_C94_n936, mult_28_C94_n935, mult_28_C94_n934, 
      mult_28_C94_n933, mult_28_C94_n932, mult_28_C94_n931, mult_28_C94_n930, 
      mult_28_C94_n929, mult_28_C94_n928, mult_28_C94_n927, mult_28_C94_n926, 
      mult_28_C94_n925, mult_28_C94_n924, mult_28_C94_n923, mult_28_C94_n922, 
      mult_28_C94_n921, mult_28_C94_n920, mult_28_C94_n919, mult_28_C94_n918, 
      mult_28_C94_n917, mult_28_C94_n916, mult_28_C94_n915, mult_28_C94_n914, 
      mult_28_C94_n913, mult_28_C94_n912, mult_28_C94_n911, mult_28_C94_n910, 
      mult_28_C94_n842, mult_28_C94_n840, mult_28_C94_n839, mult_28_C94_n838, 
      mult_28_C94_n837, mult_28_C94_n834, mult_28_C94_n833, mult_28_C94_n832, 
      mult_28_C94_n831, mult_28_C94_n830, mult_28_C94_n829, mult_28_C94_n828, 
      mult_28_C94_n827, mult_28_C94_n826, mult_28_C94_n825, mult_28_C94_n824, 
      mult_28_C94_n823, mult_28_C94_n822, mult_28_C94_n821, mult_28_C94_n820, 
      mult_28_C94_n819, mult_28_C94_n818, mult_28_C94_n817, mult_28_C94_n816, 
      mult_28_C94_n815, mult_28_C94_n814, mult_28_C94_n813, mult_28_C94_n812, 
      mult_28_C94_n811, mult_28_C94_n809, mult_28_C94_n808, mult_28_C94_n807, 
      mult_28_C94_n806, mult_28_C94_n805, mult_28_C94_n803, mult_28_C94_n802, 
      mult_28_C94_n801, mult_28_C94_n800, mult_28_C94_n799, mult_28_C94_n798, 
      mult_28_C94_n797, mult_28_C94_n796, mult_28_C94_n795, mult_28_C94_n794, 
      mult_28_C94_n793, mult_28_C94_n792, mult_28_C94_n791, mult_28_C94_n790, 
      mult_28_C94_n789, mult_28_C94_n788, mult_28_C94_n787, mult_28_C94_n786, 
      mult_28_C94_n785, mult_28_C94_n784, mult_28_C94_n783, mult_28_C94_n782, 
      mult_28_C94_n781, mult_28_C94_n780, mult_28_C94_n779, mult_28_C94_n778, 
      mult_28_C94_n777, mult_28_C94_n776, mult_28_C94_n775, mult_28_C94_n774, 
      mult_28_C94_n773, mult_28_C94_n772, mult_28_C94_n771, mult_28_C94_n770, 
      mult_28_C94_n769, mult_28_C94_n768, mult_28_C94_n767, mult_28_C94_n766, 
      mult_28_C94_n765, mult_28_C94_n764, mult_28_C94_n763, mult_28_C94_n762, 
      mult_28_C94_n761, mult_28_C94_n760, mult_28_C94_n759, mult_28_C94_n758, 
      mult_28_C94_n757, mult_28_C94_n756, mult_28_C94_n755, mult_28_C94_n754, 
      mult_28_C94_n753, mult_28_C94_n752, mult_28_C94_n751, mult_28_C94_n750, 
      mult_28_C94_n749, mult_28_C94_n748, mult_28_C94_n747, mult_28_C94_n746, 
      mult_28_C94_n745, mult_28_C94_n744, mult_28_C94_n743, mult_28_C94_n742, 
      mult_28_C94_n741, mult_28_C94_n740, mult_28_C94_n739, mult_28_C94_n738, 
      mult_28_C94_n737, mult_28_C94_n736, mult_28_C94_n735, mult_28_C94_n734, 
      mult_28_C94_n733, mult_28_C94_n732, mult_28_C94_n731, mult_28_C94_n730, 
      mult_28_C94_n729, mult_28_C94_n728, mult_28_C94_n727, mult_28_C94_n726, 
      mult_28_C94_n725, mult_28_C94_n724, mult_28_C94_n723, mult_28_C94_n722, 
      mult_28_C94_n721, mult_28_C94_n720, mult_28_C94_n719, mult_28_C94_n718, 
      mult_28_C94_n717, mult_28_C94_n716, mult_28_C94_n715, mult_28_C94_n714, 
      mult_28_C94_n713, mult_28_C94_n712, mult_28_C94_n711, mult_28_C94_n710, 
      mult_28_C94_n709, mult_28_C94_n708, mult_28_C94_n707, mult_28_C94_n706, 
      mult_28_C94_n705, mult_28_C94_n704, mult_28_C94_n703, mult_28_C94_n702, 
      mult_28_C94_n701, mult_28_C94_n700, mult_28_C94_n699, mult_28_C94_n698, 
      mult_28_C94_n697, mult_28_C94_n696, mult_28_C94_n695, mult_28_C94_n694, 
      mult_28_C94_n693, mult_28_C94_n692, mult_28_C94_n691, mult_28_C94_n690, 
      mult_28_C94_n689, mult_28_C94_n688, mult_28_C94_n687, mult_28_C94_n686, 
      mult_28_C94_n685, mult_28_C94_n684, mult_28_C94_n683, mult_28_C94_n682, 
      mult_28_C94_n681, mult_28_C94_n680, mult_28_C94_n679, mult_28_C94_n678, 
      mult_28_C94_n677, mult_28_C94_n676, mult_28_C94_n675, mult_28_C94_n674, 
      mult_28_C94_n673, mult_28_C94_n672, mult_28_C94_n671, mult_28_C94_n670, 
      mult_28_C94_n669, mult_28_C94_n668, mult_28_C94_n667, mult_28_C94_n666, 
      mult_28_C94_n665, mult_28_C94_n664, mult_28_C94_n663, mult_28_C94_n662, 
      mult_28_C94_n661, mult_28_C94_n660, mult_28_C94_n659, mult_28_C94_n658, 
      mult_28_C94_n657, mult_28_C94_n656, mult_28_C94_n655, mult_28_C94_n654, 
      mult_28_C94_n653, mult_28_C94_n652, mult_28_C94_n651, mult_28_C94_n650, 
      mult_28_C94_n649, mult_28_C94_n648, mult_28_C94_n647, mult_28_C94_n646, 
      mult_28_C94_n645, mult_28_C94_n644, mult_28_C94_n643, mult_28_C94_n642, 
      mult_28_C94_n641, mult_28_C94_n640, mult_28_C94_n639, mult_28_C94_n638, 
      mult_28_C94_n637, mult_28_C94_n636, mult_28_C94_n635, mult_28_C94_n634, 
      mult_28_C94_n633, mult_28_C94_n632, mult_28_C94_n631, mult_28_C94_n630, 
      mult_28_C94_n629, mult_28_C94_n628, mult_28_C94_n627, mult_28_C94_n626, 
      mult_28_C94_n625, mult_28_C94_n624, mult_28_C94_n623, mult_28_C94_n622, 
      mult_28_C94_n621, mult_28_C94_n620, mult_28_C94_n619, mult_28_C94_n618, 
      mult_28_C94_n617, mult_28_C94_n616, mult_28_C94_n615, mult_28_C94_n614, 
      mult_28_C94_n613, mult_28_C94_n612, mult_28_C94_n611, mult_28_C94_n610, 
      mult_28_C94_n609, mult_28_C94_n608, mult_28_C94_n607, mult_28_C94_n606, 
      mult_28_C94_n605, mult_28_C94_n604, mult_28_C94_n603, mult_28_C94_n602, 
      mult_28_C94_n601, mult_28_C94_n600, mult_28_C94_n599, mult_28_C94_n598, 
      mult_28_C94_n597, mult_28_C94_n596, mult_28_C94_n595, mult_28_C94_n594, 
      mult_28_C94_n593, mult_28_C94_n592, mult_28_C94_n591, mult_28_C94_n590, 
      mult_28_C94_n589, mult_28_C94_n588, mult_28_C94_n587, mult_28_C94_n586, 
      mult_28_C94_n585, mult_28_C94_n584, mult_28_C94_n583, mult_28_C94_n582, 
      mult_28_C94_n581, mult_28_C94_n580, mult_28_C94_n579, mult_28_C94_n578, 
      mult_28_C94_n577, mult_28_C94_n576, mult_28_C94_n575, mult_28_C94_n574, 
      mult_28_C94_n573, mult_28_C94_n572, mult_28_C94_n571, mult_28_C94_n570, 
      mult_28_C94_n569, mult_28_C94_n568, mult_28_C94_n567, mult_28_C94_n566, 
      mult_28_C94_n565, mult_28_C94_n564, mult_28_C94_n563, mult_28_C94_n562, 
      mult_28_C94_n561, mult_28_C94_n560, mult_28_C94_n559, mult_28_C94_n558, 
      mult_28_C94_n557, mult_28_C94_n556, mult_28_C94_n555, mult_28_C94_n554, 
      mult_28_C94_n553, mult_28_C94_n552, mult_28_C94_n551, mult_28_C94_n550, 
      mult_28_C94_n549, mult_28_C94_n548, mult_28_C94_n547, mult_28_C94_n546, 
      mult_28_C94_n545, mult_28_C94_n544, mult_28_C94_n543, mult_28_C94_n542, 
      mult_28_C94_n541, mult_28_C94_n540, mult_28_C94_n539, mult_28_C94_n538, 
      mult_28_C94_n537, mult_28_C94_n536, mult_28_C94_n535, mult_28_C94_n534, 
      mult_28_C94_n533, mult_28_C94_n532, mult_28_C94_n530, mult_28_C94_n529, 
      mult_28_C94_n528, mult_28_C94_n527, mult_28_C94_n526, mult_28_C94_n525, 
      mult_28_C94_n524, mult_28_C94_n523, mult_28_C94_n522, mult_28_C94_n521, 
      mult_28_C94_n520, mult_28_C94_n519, mult_28_C94_n518, mult_28_C94_n517, 
      mult_28_C94_n516, mult_28_C94_n515, mult_28_C94_n514, mult_28_C94_n513, 
      mult_28_C94_n512, mult_28_C94_n511, mult_28_C94_n510, mult_28_C94_n509, 
      mult_28_C94_n508, mult_28_C94_n507, mult_28_C94_n506, mult_28_C94_n505, 
      mult_28_C94_n504, mult_28_C94_n503, mult_28_C94_n502, mult_28_C94_n501, 
      mult_28_C94_n500, mult_28_C94_n499, mult_28_C94_n498, mult_28_C94_n497, 
      mult_28_C94_n496, mult_28_C94_n495, mult_28_C94_n494, mult_28_C94_n493, 
      mult_28_C94_n492, mult_28_C94_n491, mult_28_C94_n490, mult_28_C94_n489, 
      mult_28_C94_n488, mult_28_C94_n487, mult_28_C94_n486, mult_28_C94_n485, 
      mult_28_C94_n484, mult_28_C94_n483, mult_28_C94_n482, mult_28_C94_n481, 
      mult_28_C94_n480, mult_28_C94_n479, mult_28_C94_n478, mult_28_C94_n477, 
      mult_28_C94_n476, mult_28_C94_n475, mult_28_C94_n474, mult_28_C94_n473, 
      mult_28_C94_n472, mult_28_C94_n471, mult_28_C94_n470, mult_28_C94_n469, 
      mult_28_C94_n468, mult_28_C94_n467, mult_28_C94_n466, mult_28_C94_n465, 
      mult_28_C94_n464, mult_28_C94_n463, mult_28_C94_n462, mult_28_C94_n461, 
      mult_28_C94_n460, mult_28_C94_n459, mult_28_C94_n458, mult_28_C94_n457, 
      mult_28_C94_n456, mult_28_C94_n455, mult_28_C94_n454, mult_28_C94_n453, 
      mult_28_C94_n452, mult_28_C94_n451, mult_28_C94_n450, mult_28_C94_n449, 
      mult_28_C94_n448, mult_28_C94_n447, mult_28_C94_n446, mult_28_C94_n445, 
      mult_28_C94_n444, mult_28_C94_n443, mult_28_C94_n442, mult_28_C94_n441, 
      mult_28_C94_n440, mult_28_C94_n439, mult_28_C94_n438, mult_28_C94_n437, 
      mult_28_C94_n436, mult_28_C94_n435, mult_28_C94_n434, mult_28_C94_n433, 
      mult_28_C94_n432, mult_28_C94_n431, mult_28_C94_n430, mult_28_C94_n429, 
      mult_28_C94_n428, mult_28_C94_n427, mult_28_C94_n426, mult_28_C94_n425, 
      mult_28_C94_n424, mult_28_C94_n423, mult_28_C94_n422, mult_28_C94_n421, 
      mult_28_C94_n420, mult_28_C94_n419, mult_28_C94_n418, mult_28_C94_n417, 
      mult_28_C94_n416, mult_28_C94_n415, mult_28_C94_n414, mult_28_C94_n413, 
      mult_28_C94_n412, mult_28_C94_n411, mult_28_C94_n410, mult_28_C94_n409, 
      mult_28_C94_n408, mult_28_C94_n407, mult_28_C94_n406, mult_28_C94_n405, 
      mult_28_C94_n404, mult_28_C94_n403, mult_28_C94_n402, mult_28_C94_n401, 
      mult_28_C94_n400, mult_28_C94_n399, mult_28_C94_n398, mult_28_C94_n397, 
      mult_28_C94_n396, mult_28_C94_n395, mult_28_C94_n394, mult_28_C94_n393, 
      mult_28_C94_n392, mult_28_C94_n391, mult_28_C94_n390, mult_28_C94_n389, 
      mult_28_C94_n388, mult_28_C94_n387, mult_28_C94_n386, mult_28_C94_n385, 
      mult_28_C94_n384, mult_28_C94_n383, mult_28_C94_n382, mult_28_C94_n381, 
      mult_28_C94_n380, mult_28_C94_n379, mult_28_C94_n378, mult_28_C94_n377, 
      mult_28_C94_n376, mult_28_C94_n375, mult_28_C94_n374, mult_28_C94_n373, 
      mult_28_C94_n372, mult_28_C94_n371, mult_28_C94_n370, mult_28_C94_n369, 
      mult_28_C94_n368, mult_28_C94_n367, mult_28_C94_n366, mult_28_C94_n365, 
      mult_28_C94_n364, mult_28_C94_n363, mult_28_C94_n362, mult_28_C94_n361, 
      mult_28_C94_n360, mult_28_C94_n359, mult_28_C94_n358, mult_28_C94_n357, 
      mult_28_C94_n356, mult_28_C94_n355, mult_28_C94_n354, mult_28_C94_n353, 
      mult_28_C94_n352, mult_28_C94_n351, mult_28_C94_n350, mult_28_C94_n349, 
      mult_28_C94_n348, mult_28_C94_n347, mult_28_C94_n346, mult_28_C94_n345, 
      mult_28_C94_n344, mult_28_C94_n343, mult_28_C94_n342, mult_28_C94_n341, 
      mult_28_C94_n340, mult_28_C94_n339, mult_28_C94_n338, mult_28_C94_n337, 
      mult_28_C94_n336, mult_28_C94_n335, mult_28_C94_n334, mult_28_C94_n333, 
      mult_28_C94_n332, mult_28_C94_n331, mult_28_C94_n330, mult_28_C94_n329, 
      mult_28_C94_n328, mult_28_C94_n327, mult_28_C94_n326, mult_28_C94_n325, 
      mult_28_C94_n324, mult_28_C94_n323, mult_28_C94_n322, mult_28_C94_n321, 
      mult_28_C94_n320, mult_28_C94_n319, mult_28_C94_n318, mult_28_C94_n317, 
      mult_28_C94_n316, mult_28_C94_n315, mult_28_C94_n294, mult_28_C94_n277, 
      mult_28_C94_n276, mult_28_C94_n275, mult_28_C94_n274, mult_28_C94_n269, 
      mult_28_C94_n268, mult_28_C94_n267, mult_28_C94_n266, mult_28_C94_n261, 
      mult_28_C94_n250, mult_28_C94_n249, mult_28_C94_n248, mult_28_C94_n243, 
      mult_28_C94_n232, mult_28_C94_n231, mult_28_C94_n230, mult_28_C94_n229, 
      mult_28_C94_n217, mult_28_C94_n216, mult_28_C94_n215, mult_28_C94_n214, 
      mult_28_C94_n213, mult_28_C94_n210, mult_28_C94_n209, mult_28_C94_n208, 
      mult_28_C94_n207, mult_28_C94_n206, mult_28_C94_n205, mult_28_C94_n204, 
      mult_28_C94_n203, mult_28_C94_n202, mult_28_C94_n201, mult_28_C94_n200, 
      mult_28_C94_n199, mult_28_C94_n198, mult_28_C94_n197, mult_28_C94_n195, 
      mult_28_C94_n194, mult_28_C94_n193, mult_28_C94_n192, mult_28_C94_n191, 
      mult_28_C94_n190, mult_28_C94_n189, mult_28_C94_n188, mult_28_C94_n187, 
      mult_28_C94_n186, mult_28_C94_n185, mult_28_C94_n184, mult_28_C94_n183, 
      mult_28_C94_n182, mult_28_C94_n181, mult_28_C94_n180, mult_28_C94_n179, 
      mult_28_C94_n178, mult_28_C94_n177, mult_28_C94_n176, mult_28_C94_n175, 
      mult_28_C94_n174, mult_28_C94_n173, mult_28_C94_n172, mult_28_C94_n171, 
      mult_28_C94_n170, mult_28_C94_n168, mult_28_C94_n167, mult_28_C94_n166, 
      mult_28_C94_n165, mult_28_C94_n164, mult_28_C94_n163, mult_28_C94_n162, 
      mult_28_C94_n161, mult_28_C94_n160, mult_28_C94_n159, mult_28_C94_n158, 
      mult_28_C94_n157, mult_28_C94_n156, mult_28_C94_n155, mult_28_C94_n154, 
      mult_28_C94_n152, mult_28_C94_n151, mult_28_C94_n150, mult_28_C94_n149, 
      mult_28_C94_n148, mult_28_C94_n147, mult_28_C94_n146, mult_28_C94_n145, 
      mult_28_C94_n144, mult_28_C94_n143, mult_28_C94_n142, mult_28_C94_n141, 
      mult_28_C94_n139, mult_28_C94_n136, mult_28_C94_n135, mult_28_C94_n134, 
      mult_28_C94_n133, mult_28_C94_n132, mult_28_C94_n129, mult_28_C94_n128, 
      mult_28_C94_n127, mult_28_C94_n126, mult_28_C94_n125, mult_28_C94_n124, 
      mult_28_C94_n123, mult_28_C94_n121, mult_28_C94_n116, mult_28_C94_n115, 
      mult_28_C94_n114, mult_28_C94_n113, mult_28_C94_n112, mult_28_C94_n110, 
      mult_28_C94_n109, mult_28_C94_n108, mult_28_C94_n107, mult_28_C94_n106, 
      mult_28_C94_n105, mult_28_C94_n104, mult_28_C94_n103, mult_28_C94_n102, 
      mult_28_C94_n101, mult_28_C94_n100, mult_28_C94_n99, mult_28_C94_n96, 
      mult_28_C94_n95, mult_28_C94_n94, mult_28_C94_n93, mult_28_C94_n92, 
      mult_28_C94_n87, mult_28_C94_n86, mult_28_C94_n85, mult_28_C94_n84, 
      mult_28_C94_n69, mult_28_C94_n68, mult_28_C94_n67, mult_28_C94_n66, 
      mult_28_C94_n65, mult_28_C94_n64, mult_28_C94_n62, mult_28_C94_n61, 
      mult_28_C94_n60, mult_28_C94_n59, mult_28_C94_n58, mult_28_C94_n57, 
      mult_28_C94_n56, mult_28_C94_n55, mult_28_C94_n54, mult_28_C94_n51, 
      mult_28_C94_n48, mult_28_C94_n47, mult_28_C94_n46, mult_28_C94_n45, 
      mult_28_C94_n43, mult_28_C94_n42, mult_28_C94_n41, mult_28_C94_n40, 
      mult_28_C94_n39, mult_28_C94_n37, mult_28_C94_n36, mult_28_C94_n35, 
      mult_28_C94_n34, mult_28_C94_n33, mult_28_C94_n31, mult_28_C94_n30, 
      mult_28_C94_n29, mult_28_C94_n28, mult_28_C94_n27, mult_28_C94_n25, 
      mult_28_C94_n24, mult_28_C94_n23, mult_28_C94_n22, mult_28_C94_n21, 
      mult_28_C94_n19, mult_28_C94_n18, mult_28_C94_n17, mult_28_C94_n16, 
      mult_28_C94_n15, mult_28_C94_n13, mult_28_C94_n12, mult_28_C94_n11, 
      mult_28_C94_n10, mult_28_C94_n9, mult_28_C94_n7, mult_28_C94_n6, 
      mult_28_C94_n5, mult_28_C94_n4, mult_28_C94_n3, mult_28_C94_n1, 
      mult_28_C93_n938, mult_28_C93_n937, mult_28_C93_n936, mult_28_C93_n935, 
      mult_28_C93_n934, mult_28_C93_n933, mult_28_C93_n932, mult_28_C93_n931, 
      mult_28_C93_n930, mult_28_C93_n929, mult_28_C93_n928, mult_28_C93_n927, 
      mult_28_C93_n926, mult_28_C93_n925, mult_28_C93_n924, mult_28_C93_n923, 
      mult_28_C93_n922, mult_28_C93_n921, mult_28_C93_n920, mult_28_C93_n919, 
      mult_28_C93_n918, mult_28_C93_n917, mult_28_C93_n916, mult_28_C93_n915, 
      mult_28_C93_n914, mult_28_C93_n913, mult_28_C93_n912, mult_28_C93_n911, 
      mult_28_C93_n910, mult_28_C93_n842, mult_28_C93_n840, mult_28_C93_n839, 
      mult_28_C93_n838, mult_28_C93_n837, mult_28_C93_n834, mult_28_C93_n833, 
      mult_28_C93_n832, mult_28_C93_n831, mult_28_C93_n830, mult_28_C93_n829, 
      mult_28_C93_n828, mult_28_C93_n827, mult_28_C93_n826, mult_28_C93_n825, 
      mult_28_C93_n824, mult_28_C93_n823, mult_28_C93_n822, mult_28_C93_n821, 
      mult_28_C93_n820, mult_28_C93_n819, mult_28_C93_n818, mult_28_C93_n817, 
      mult_28_C93_n816, mult_28_C93_n815, mult_28_C93_n814, mult_28_C93_n813, 
      mult_28_C93_n812, mult_28_C93_n811, mult_28_C93_n809, mult_28_C93_n808, 
      mult_28_C93_n807, mult_28_C93_n806, mult_28_C93_n805, mult_28_C93_n803, 
      mult_28_C93_n802, mult_28_C93_n801, mult_28_C93_n800, mult_28_C93_n799, 
      mult_28_C93_n798, mult_28_C93_n797, mult_28_C93_n796, mult_28_C93_n795, 
      mult_28_C93_n794, mult_28_C93_n793, mult_28_C93_n792, mult_28_C93_n791, 
      mult_28_C93_n790, mult_28_C93_n789, mult_28_C93_n788, mult_28_C93_n787, 
      mult_28_C93_n786, mult_28_C93_n785, mult_28_C93_n784, mult_28_C93_n783, 
      mult_28_C93_n782, mult_28_C93_n781, mult_28_C93_n780, mult_28_C93_n779, 
      mult_28_C93_n778, mult_28_C93_n777, mult_28_C93_n776, mult_28_C93_n775, 
      mult_28_C93_n774, mult_28_C93_n773, mult_28_C93_n772, mult_28_C93_n771, 
      mult_28_C93_n770, mult_28_C93_n769, mult_28_C93_n768, mult_28_C93_n767, 
      mult_28_C93_n766, mult_28_C93_n765, mult_28_C93_n764, mult_28_C93_n763, 
      mult_28_C93_n762, mult_28_C93_n761, mult_28_C93_n760, mult_28_C93_n759, 
      mult_28_C93_n758, mult_28_C93_n757, mult_28_C93_n756, mult_28_C93_n755, 
      mult_28_C93_n754, mult_28_C93_n753, mult_28_C93_n752, mult_28_C93_n751, 
      mult_28_C93_n750, mult_28_C93_n749, mult_28_C93_n748, mult_28_C93_n747, 
      mult_28_C93_n746, mult_28_C93_n745, mult_28_C93_n744, mult_28_C93_n743, 
      mult_28_C93_n742, mult_28_C93_n741, mult_28_C93_n740, mult_28_C93_n739, 
      mult_28_C93_n738, mult_28_C93_n737, mult_28_C93_n736, mult_28_C93_n735, 
      mult_28_C93_n734, mult_28_C93_n733, mult_28_C93_n732, mult_28_C93_n731, 
      mult_28_C93_n730, mult_28_C93_n729, mult_28_C93_n728, mult_28_C93_n727, 
      mult_28_C93_n726, mult_28_C93_n725, mult_28_C93_n724, mult_28_C93_n723, 
      mult_28_C93_n722, mult_28_C93_n721, mult_28_C93_n720, mult_28_C93_n719, 
      mult_28_C93_n718, mult_28_C93_n717, mult_28_C93_n716, mult_28_C93_n715, 
      mult_28_C93_n714, mult_28_C93_n713, mult_28_C93_n712, mult_28_C93_n711, 
      mult_28_C93_n710, mult_28_C93_n709, mult_28_C93_n708, mult_28_C93_n707, 
      mult_28_C93_n706, mult_28_C93_n705, mult_28_C93_n704, mult_28_C93_n703, 
      mult_28_C93_n702, mult_28_C93_n701, mult_28_C93_n700, mult_28_C93_n699, 
      mult_28_C93_n698, mult_28_C93_n697, mult_28_C93_n696, mult_28_C93_n695, 
      mult_28_C93_n694, mult_28_C93_n693, mult_28_C93_n692, mult_28_C93_n691, 
      mult_28_C93_n690, mult_28_C93_n689, mult_28_C93_n688, mult_28_C93_n687, 
      mult_28_C93_n686, mult_28_C93_n685, mult_28_C93_n684, mult_28_C93_n683, 
      mult_28_C93_n682, mult_28_C93_n681, mult_28_C93_n680, mult_28_C93_n679, 
      mult_28_C93_n678, mult_28_C93_n677, mult_28_C93_n676, mult_28_C93_n675, 
      mult_28_C93_n674, mult_28_C93_n673, mult_28_C93_n672, mult_28_C93_n671, 
      mult_28_C93_n670, mult_28_C93_n669, mult_28_C93_n668, mult_28_C93_n667, 
      mult_28_C93_n666, mult_28_C93_n665, mult_28_C93_n664, mult_28_C93_n663, 
      mult_28_C93_n662, mult_28_C93_n661, mult_28_C93_n660, mult_28_C93_n659, 
      mult_28_C93_n658, mult_28_C93_n657, mult_28_C93_n656, mult_28_C93_n655, 
      mult_28_C93_n654, mult_28_C93_n653, mult_28_C93_n652, mult_28_C93_n651, 
      mult_28_C93_n650, mult_28_C93_n649, mult_28_C93_n648, mult_28_C93_n647, 
      mult_28_C93_n646, mult_28_C93_n645, mult_28_C93_n644, mult_28_C93_n643, 
      mult_28_C93_n642, mult_28_C93_n641, mult_28_C93_n640, mult_28_C93_n639, 
      mult_28_C93_n638, mult_28_C93_n637, mult_28_C93_n636, mult_28_C93_n635, 
      mult_28_C93_n634, mult_28_C93_n633, mult_28_C93_n632, mult_28_C93_n631, 
      mult_28_C93_n630, mult_28_C93_n629, mult_28_C93_n628, mult_28_C93_n627, 
      mult_28_C93_n626, mult_28_C93_n625, mult_28_C93_n624, mult_28_C93_n623, 
      mult_28_C93_n622, mult_28_C93_n621, mult_28_C93_n620, mult_28_C93_n619, 
      mult_28_C93_n618, mult_28_C93_n617, mult_28_C93_n616, mult_28_C93_n615, 
      mult_28_C93_n614, mult_28_C93_n613, mult_28_C93_n612, mult_28_C93_n611, 
      mult_28_C93_n610, mult_28_C93_n609, mult_28_C93_n608, mult_28_C93_n607, 
      mult_28_C93_n606, mult_28_C93_n605, mult_28_C93_n604, mult_28_C93_n603, 
      mult_28_C93_n602, mult_28_C93_n601, mult_28_C93_n600, mult_28_C93_n599, 
      mult_28_C93_n598, mult_28_C93_n597, mult_28_C93_n596, mult_28_C93_n595, 
      mult_28_C93_n594, mult_28_C93_n593, mult_28_C93_n592, mult_28_C93_n591, 
      mult_28_C93_n590, mult_28_C93_n589, mult_28_C93_n588, mult_28_C93_n587, 
      mult_28_C93_n586, mult_28_C93_n585, mult_28_C93_n584, mult_28_C93_n583, 
      mult_28_C93_n582, mult_28_C93_n581, mult_28_C93_n580, mult_28_C93_n579, 
      mult_28_C93_n578, mult_28_C93_n577, mult_28_C93_n576, mult_28_C93_n575, 
      mult_28_C93_n574, mult_28_C93_n573, mult_28_C93_n572, mult_28_C93_n571, 
      mult_28_C93_n570, mult_28_C93_n569, mult_28_C93_n568, mult_28_C93_n567, 
      mult_28_C93_n566, mult_28_C93_n565, mult_28_C93_n564, mult_28_C93_n563, 
      mult_28_C93_n562, mult_28_C93_n561, mult_28_C93_n560, mult_28_C93_n559, 
      mult_28_C93_n558, mult_28_C93_n557, mult_28_C93_n556, mult_28_C93_n555, 
      mult_28_C93_n554, mult_28_C93_n553, mult_28_C93_n552, mult_28_C93_n551, 
      mult_28_C93_n550, mult_28_C93_n549, mult_28_C93_n548, mult_28_C93_n547, 
      mult_28_C93_n546, mult_28_C93_n545, mult_28_C93_n544, mult_28_C93_n543, 
      mult_28_C93_n542, mult_28_C93_n541, mult_28_C93_n540, mult_28_C93_n539, 
      mult_28_C93_n538, mult_28_C93_n537, mult_28_C93_n536, mult_28_C93_n535, 
      mult_28_C93_n534, mult_28_C93_n533, mult_28_C93_n532, mult_28_C93_n530, 
      mult_28_C93_n529, mult_28_C93_n528, mult_28_C93_n527, mult_28_C93_n526, 
      mult_28_C93_n525, mult_28_C93_n524, mult_28_C93_n523, mult_28_C93_n522, 
      mult_28_C93_n521, mult_28_C93_n520, mult_28_C93_n519, mult_28_C93_n518, 
      mult_28_C93_n517, mult_28_C93_n516, mult_28_C93_n515, mult_28_C93_n514, 
      mult_28_C93_n513, mult_28_C93_n512, mult_28_C93_n511, mult_28_C93_n510, 
      mult_28_C93_n509, mult_28_C93_n508, mult_28_C93_n507, mult_28_C93_n506, 
      mult_28_C93_n505, mult_28_C93_n504, mult_28_C93_n503, mult_28_C93_n502, 
      mult_28_C93_n501, mult_28_C93_n500, mult_28_C93_n499, mult_28_C93_n498, 
      mult_28_C93_n497, mult_28_C93_n496, mult_28_C93_n495, mult_28_C93_n494, 
      mult_28_C93_n493, mult_28_C93_n492, mult_28_C93_n491, mult_28_C93_n490, 
      mult_28_C93_n489, mult_28_C93_n488, mult_28_C93_n487, mult_28_C93_n486, 
      mult_28_C93_n485, mult_28_C93_n484, mult_28_C93_n483, mult_28_C93_n482, 
      mult_28_C93_n481, mult_28_C93_n480, mult_28_C93_n479, mult_28_C93_n478, 
      mult_28_C93_n477, mult_28_C93_n476, mult_28_C93_n475, mult_28_C93_n474, 
      mult_28_C93_n473, mult_28_C93_n472, mult_28_C93_n471, mult_28_C93_n470, 
      mult_28_C93_n469, mult_28_C93_n468, mult_28_C93_n467, mult_28_C93_n466, 
      mult_28_C93_n465, mult_28_C93_n464, mult_28_C93_n463, mult_28_C93_n462, 
      mult_28_C93_n461, mult_28_C93_n460, mult_28_C93_n459, mult_28_C93_n458, 
      mult_28_C93_n457, mult_28_C93_n456, mult_28_C93_n455, mult_28_C93_n454, 
      mult_28_C93_n453, mult_28_C93_n452, mult_28_C93_n451, mult_28_C93_n450, 
      mult_28_C93_n449, mult_28_C93_n448, mult_28_C93_n447, mult_28_C93_n446, 
      mult_28_C93_n445, mult_28_C93_n444, mult_28_C93_n443, mult_28_C93_n442, 
      mult_28_C93_n441, mult_28_C93_n440, mult_28_C93_n439, mult_28_C93_n438, 
      mult_28_C93_n437, mult_28_C93_n436, mult_28_C93_n435, mult_28_C93_n434, 
      mult_28_C93_n433, mult_28_C93_n432, mult_28_C93_n431, mult_28_C93_n430, 
      mult_28_C93_n429, mult_28_C93_n428, mult_28_C93_n427, mult_28_C93_n426, 
      mult_28_C93_n425, mult_28_C93_n424, mult_28_C93_n423, mult_28_C93_n422, 
      mult_28_C93_n421, mult_28_C93_n420, mult_28_C93_n419, mult_28_C93_n418, 
      mult_28_C93_n417, mult_28_C93_n416, mult_28_C93_n415, mult_28_C93_n414, 
      mult_28_C93_n413, mult_28_C93_n412, mult_28_C93_n411, mult_28_C93_n410, 
      mult_28_C93_n409, mult_28_C93_n408, mult_28_C93_n407, mult_28_C93_n406, 
      mult_28_C93_n405, mult_28_C93_n404, mult_28_C93_n403, mult_28_C93_n402, 
      mult_28_C93_n401, mult_28_C93_n400, mult_28_C93_n399, mult_28_C93_n398, 
      mult_28_C93_n397, mult_28_C93_n396, mult_28_C93_n395, mult_28_C93_n394, 
      mult_28_C93_n393, mult_28_C93_n392, mult_28_C93_n391, mult_28_C93_n390, 
      mult_28_C93_n389, mult_28_C93_n388, mult_28_C93_n387, mult_28_C93_n386, 
      mult_28_C93_n385, mult_28_C93_n384, mult_28_C93_n383, mult_28_C93_n382, 
      mult_28_C93_n381, mult_28_C93_n380, mult_28_C93_n379, mult_28_C93_n378, 
      mult_28_C93_n377, mult_28_C93_n376, mult_28_C93_n375, mult_28_C93_n374, 
      mult_28_C93_n373, mult_28_C93_n372, mult_28_C93_n371, mult_28_C93_n370, 
      mult_28_C93_n369, mult_28_C93_n368, mult_28_C93_n367, mult_28_C93_n366, 
      mult_28_C93_n365, mult_28_C93_n364, mult_28_C93_n363, mult_28_C93_n362, 
      mult_28_C93_n361, mult_28_C93_n360, mult_28_C93_n359, mult_28_C93_n358, 
      mult_28_C93_n357, mult_28_C93_n356, mult_28_C93_n355, mult_28_C93_n354, 
      mult_28_C93_n353, mult_28_C93_n352, mult_28_C93_n351, mult_28_C93_n350, 
      mult_28_C93_n349, mult_28_C93_n348, mult_28_C93_n347, mult_28_C93_n346, 
      mult_28_C93_n345, mult_28_C93_n344, mult_28_C93_n343, mult_28_C93_n342, 
      mult_28_C93_n341, mult_28_C93_n340, mult_28_C93_n339, mult_28_C93_n338, 
      mult_28_C93_n337, mult_28_C93_n336, mult_28_C93_n335, mult_28_C93_n334, 
      mult_28_C93_n333, mult_28_C93_n332, mult_28_C93_n331, mult_28_C93_n330, 
      mult_28_C93_n329, mult_28_C93_n328, mult_28_C93_n327, mult_28_C93_n326, 
      mult_28_C93_n325, mult_28_C93_n324, mult_28_C93_n323, mult_28_C93_n322, 
      mult_28_C93_n321, mult_28_C93_n320, mult_28_C93_n319, mult_28_C93_n318, 
      mult_28_C93_n317, mult_28_C93_n316, mult_28_C93_n315, mult_28_C93_n298, 
      mult_28_C93_n297, mult_28_C93_n296, mult_28_C93_n294, mult_28_C93_n293, 
      mult_28_C93_n292, mult_28_C93_n277, mult_28_C93_n276, mult_28_C93_n275, 
      mult_28_C93_n274, mult_28_C93_n269, mult_28_C93_n268, mult_28_C93_n267, 
      mult_28_C93_n266, mult_28_C93_n261, mult_28_C93_n250, mult_28_C93_n249, 
      mult_28_C93_n248, mult_28_C93_n243, mult_28_C93_n232, mult_28_C93_n231, 
      mult_28_C93_n230, mult_28_C93_n229, mult_28_C93_n217, mult_28_C93_n216, 
      mult_28_C93_n215, mult_28_C93_n214, mult_28_C93_n213, mult_28_C93_n210, 
      mult_28_C93_n209, mult_28_C93_n208, mult_28_C93_n207, mult_28_C93_n206, 
      mult_28_C93_n205, mult_28_C93_n204, mult_28_C93_n203, mult_28_C93_n202, 
      mult_28_C93_n201, mult_28_C93_n200, mult_28_C93_n199, mult_28_C93_n198, 
      mult_28_C93_n197, mult_28_C93_n195, mult_28_C93_n194, mult_28_C93_n193, 
      mult_28_C93_n192, mult_28_C93_n191, mult_28_C93_n190, mult_28_C93_n189, 
      mult_28_C93_n188, mult_28_C93_n187, mult_28_C93_n186, mult_28_C93_n185, 
      mult_28_C93_n184, mult_28_C93_n183, mult_28_C93_n182, mult_28_C93_n181, 
      mult_28_C93_n180, mult_28_C93_n179, mult_28_C93_n178, mult_28_C93_n177, 
      mult_28_C93_n176, mult_28_C93_n175, mult_28_C93_n174, mult_28_C93_n173, 
      mult_28_C93_n172, mult_28_C93_n171, mult_28_C93_n170, mult_28_C93_n169, 
      mult_28_C93_n168, mult_28_C93_n167, mult_28_C93_n166, mult_28_C93_n165, 
      mult_28_C93_n164, mult_28_C93_n163, mult_28_C93_n161, mult_28_C93_n160, 
      mult_28_C93_n159, mult_28_C93_n158, mult_28_C93_n157, mult_28_C93_n156, 
      mult_28_C93_n155, mult_28_C93_n152, mult_28_C93_n151, mult_28_C93_n150, 
      mult_28_C93_n149, mult_28_C93_n148, mult_28_C93_n147, mult_28_C93_n146, 
      mult_28_C93_n145, mult_28_C93_n144, mult_28_C93_n143, mult_28_C93_n142, 
      mult_28_C93_n141, mult_28_C93_n140, mult_28_C93_n139, mult_28_C93_n138, 
      mult_28_C93_n136, mult_28_C93_n135, mult_28_C93_n134, mult_28_C93_n133, 
      mult_28_C93_n132, mult_28_C93_n131, mult_28_C93_n130, mult_28_C93_n129, 
      mult_28_C93_n128, mult_28_C93_n127, mult_28_C93_n126, mult_28_C93_n125, 
      mult_28_C93_n124, mult_28_C93_n123, mult_28_C93_n117, mult_28_C93_n116, 
      mult_28_C93_n115, mult_28_C93_n114, mult_28_C93_n113, mult_28_C93_n112, 
      mult_28_C93_n110, mult_28_C93_n109, mult_28_C93_n108, mult_28_C93_n107, 
      mult_28_C93_n106, mult_28_C93_n105, mult_28_C93_n104, mult_28_C93_n103, 
      mult_28_C93_n102, mult_28_C93_n101, mult_28_C93_n100, mult_28_C93_n99, 
      mult_28_C93_n98, mult_28_C93_n97, mult_28_C93_n96, mult_28_C93_n95, 
      mult_28_C93_n94, mult_28_C93_n93, mult_28_C93_n92, mult_28_C93_n87, 
      mult_28_C93_n86, mult_28_C93_n85, mult_28_C93_n84, mult_28_C93_n69, 
      mult_28_C93_n68, mult_28_C93_n67, mult_28_C93_n66, mult_28_C93_n65, 
      mult_28_C93_n64, mult_28_C93_n63, mult_28_C93_n62, mult_28_C93_n60, 
      mult_28_C93_n59, mult_28_C93_n58, mult_28_C93_n57, mult_28_C93_n56, 
      mult_28_C93_n55, mult_28_C93_n54, mult_28_C93_n52, mult_28_C93_n51, 
      mult_28_C93_n48, mult_28_C93_n47, mult_28_C93_n46, mult_28_C93_n45, 
      mult_28_C93_n43, mult_28_C93_n42, mult_28_C93_n41, mult_28_C93_n40, 
      mult_28_C93_n39, mult_28_C93_n37, mult_28_C93_n36, mult_28_C93_n35, 
      mult_28_C93_n34, mult_28_C93_n33, mult_28_C93_n31, mult_28_C93_n30, 
      mult_28_C93_n29, mult_28_C93_n28, mult_28_C93_n27, mult_28_C93_n25, 
      mult_28_C93_n24, mult_28_C93_n23, mult_28_C93_n22, mult_28_C93_n21, 
      mult_28_C93_n19, mult_28_C93_n18, mult_28_C93_n17, mult_28_C93_n16, 
      mult_28_C93_n15, mult_28_C93_n13, mult_28_C93_n12, mult_28_C93_n11, 
      mult_28_C93_n10, mult_28_C93_n9, mult_28_C93_n7, mult_28_C93_n6, 
      mult_28_C93_n5, mult_28_C93_n4, mult_28_C93_n3, mult_28_C93_n1, 
      add_1_root_add_0_root_add_101_n193, add_1_root_add_0_root_add_101_n191, 
      add_1_root_add_0_root_add_101_n190, add_1_root_add_0_root_add_101_n189, 
      add_1_root_add_0_root_add_101_n130, add_1_root_add_0_root_add_101_n128, 
      add_1_root_add_0_root_add_101_n126, add_1_root_add_0_root_add_101_n124, 
      add_1_root_add_0_root_add_101_n122, add_1_root_add_0_root_add_101_n117, 
      add_1_root_add_0_root_add_101_n115, add_1_root_add_0_root_add_101_n114, 
      add_1_root_add_0_root_add_101_n113, add_1_root_add_0_root_add_101_n112, 
      add_1_root_add_0_root_add_101_n111, add_1_root_add_0_root_add_101_n110, 
      add_1_root_add_0_root_add_101_n109, add_1_root_add_0_root_add_101_n108, 
      add_1_root_add_0_root_add_101_n107, add_1_root_add_0_root_add_101_n104, 
      add_1_root_add_0_root_add_101_n103, add_1_root_add_0_root_add_101_n102, 
      add_1_root_add_0_root_add_101_n101, add_1_root_add_0_root_add_101_n100, 
      add_1_root_add_0_root_add_101_n99, add_1_root_add_0_root_add_101_n98, 
      add_1_root_add_0_root_add_101_n97, add_1_root_add_0_root_add_101_n96, 
      add_1_root_add_0_root_add_101_n95, add_1_root_add_0_root_add_101_n94, 
      add_1_root_add_0_root_add_101_n93, add_1_root_add_0_root_add_101_n92, 
      add_1_root_add_0_root_add_101_n89, add_1_root_add_0_root_add_101_n88, 
      add_1_root_add_0_root_add_101_n87, add_1_root_add_0_root_add_101_n86, 
      add_1_root_add_0_root_add_101_n85, add_1_root_add_0_root_add_101_n84, 
      add_1_root_add_0_root_add_101_n83, add_1_root_add_0_root_add_101_n82, 
      add_1_root_add_0_root_add_101_n81, add_1_root_add_0_root_add_101_n80, 
      add_1_root_add_0_root_add_101_n79, add_1_root_add_0_root_add_101_n78, 
      add_1_root_add_0_root_add_101_n77, add_1_root_add_0_root_add_101_n76, 
      add_1_root_add_0_root_add_101_n75, add_1_root_add_0_root_add_101_n74, 
      add_1_root_add_0_root_add_101_n73, add_1_root_add_0_root_add_101_n72, 
      add_1_root_add_0_root_add_101_n71, add_1_root_add_0_root_add_101_n70, 
      add_1_root_add_0_root_add_101_n69, add_1_root_add_0_root_add_101_n68, 
      add_1_root_add_0_root_add_101_n67, add_1_root_add_0_root_add_101_n66, 
      add_1_root_add_0_root_add_101_n65, add_1_root_add_0_root_add_101_n64, 
      add_1_root_add_0_root_add_101_n63, add_1_root_add_0_root_add_101_n62, 
      add_1_root_add_0_root_add_101_n61, add_1_root_add_0_root_add_101_n60, 
      add_1_root_add_0_root_add_101_n59, add_1_root_add_0_root_add_101_n58, 
      add_1_root_add_0_root_add_101_n57, add_1_root_add_0_root_add_101_n56, 
      add_1_root_add_0_root_add_101_n55, add_1_root_add_0_root_add_101_n54, 
      add_1_root_add_0_root_add_101_n53, add_1_root_add_0_root_add_101_n52, 
      add_1_root_add_0_root_add_101_n51, add_1_root_add_0_root_add_101_n50, 
      add_1_root_add_0_root_add_101_n49, add_1_root_add_0_root_add_101_n48, 
      add_1_root_add_0_root_add_101_n47, add_1_root_add_0_root_add_101_n46, 
      add_1_root_add_0_root_add_101_n45, add_1_root_add_0_root_add_101_n44, 
      add_1_root_add_0_root_add_101_n43, add_1_root_add_0_root_add_101_n42, 
      add_1_root_add_0_root_add_101_n41, add_1_root_add_0_root_add_101_n40, 
      add_1_root_add_0_root_add_101_n39, add_1_root_add_0_root_add_101_n38, 
      add_1_root_add_0_root_add_101_n37, add_1_root_add_0_root_add_101_n36, 
      add_1_root_add_0_root_add_101_n35, add_1_root_add_0_root_add_101_n34, 
      add_1_root_add_0_root_add_101_n33, add_1_root_add_0_root_add_101_n32, 
      add_1_root_add_0_root_add_101_n31, add_1_root_add_0_root_add_101_n30, 
      add_1_root_add_0_root_add_101_n29, add_1_root_add_0_root_add_101_n27, 
      add_1_root_add_0_root_add_101_n26, add_1_root_add_0_root_add_101_n25, 
      add_1_root_add_0_root_add_101_n24, add_1_root_add_0_root_add_101_n23, 
      add_1_root_add_0_root_add_101_n22, add_1_root_add_0_root_add_101_n21, 
      add_1_root_add_0_root_add_101_n18, add_1_root_add_0_root_add_101_n17, 
      add_1_root_add_0_root_add_101_n16, add_1_root_add_0_root_add_101_n15, 
      add_1_root_add_0_root_add_101_n14, add_1_root_add_0_root_add_101_n13, 
      add_1_root_add_0_root_add_101_n12, add_1_root_add_0_root_add_101_n11, 
      add_1_root_add_0_root_add_101_n10, add_1_root_add_0_root_add_101_n9, 
      add_1_root_add_0_root_add_101_n8, add_1_root_add_0_root_add_101_n7, 
      add_1_root_add_0_root_add_101_n6, add_1_root_add_0_root_add_101_n5, 
      add_1_root_add_0_root_add_101_n4, add_1_root_add_0_root_add_101_n3, 
      add_1_root_add_0_root_add_101_n2, add_1_root_add_0_root_add_101_n1, 
      mult_28_C92_n1157, mult_28_C92_n1156, mult_28_C92_n1155, 
      mult_28_C92_n1154, mult_28_C92_n1153, mult_28_C92_n1152, 
      mult_28_C92_n1151, mult_28_C92_n1150, mult_28_C92_n1149, 
      mult_28_C92_n1148, mult_28_C92_n1147, mult_28_C92_n1146, 
      mult_28_C92_n1145, mult_28_C92_n1144, mult_28_C92_n1143, 
      mult_28_C92_n1142, mult_28_C92_n1141, mult_28_C92_n1140, 
      mult_28_C92_n1139, mult_28_C92_n1138, mult_28_C92_n1137, 
      mult_28_C92_n1136, mult_28_C92_n1135, mult_28_C92_n1134, 
      mult_28_C92_n1133, mult_28_C92_n1132, mult_28_C92_n1131, 
      mult_28_C92_n1130, mult_28_C92_n1129, mult_28_C92_n1128, 
      mult_28_C92_n1127, mult_28_C92_n1126, mult_28_C92_n1125, 
      mult_28_C92_n1124, mult_28_C92_n1123, mult_28_C92_n1122, 
      mult_28_C92_n1121, mult_28_C92_n1120, mult_28_C92_n1119, 
      mult_28_C92_n1118, mult_28_C92_n1117, mult_28_C92_n1116, 
      mult_28_C92_n1115, mult_28_C92_n1114, mult_28_C92_n1113, 
      mult_28_C92_n1112, mult_28_C92_n1111, mult_28_C92_n1110, 
      mult_28_C92_n1109, mult_28_C92_n1108, mult_28_C92_n1107, 
      mult_28_C92_n1106, mult_28_C92_n1105, mult_28_C92_n1104, 
      mult_28_C92_n1103, mult_28_C92_n1102, mult_28_C92_n1101, 
      mult_28_C92_n1100, mult_28_C92_n1099, mult_28_C92_n1098, 
      mult_28_C92_n1097, mult_28_C92_n1096, mult_28_C92_n1095, 
      mult_28_C92_n1094, mult_28_C92_n1093, mult_28_C92_n1092, 
      mult_28_C92_n1091, mult_28_C92_n1090, mult_28_C92_n1089, 
      mult_28_C92_n1088, mult_28_C92_n1087, mult_28_C92_n1086, 
      mult_28_C92_n1085, mult_28_C92_n1084, mult_28_C92_n1083, 
      mult_28_C92_n1082, mult_28_C92_n1081, mult_28_C92_n1080, 
      mult_28_C92_n1079, mult_28_C92_n1078, mult_28_C92_n1077, 
      mult_28_C92_n1076, mult_28_C92_n1075, mult_28_C92_n1074, 
      mult_28_C92_n1073, mult_28_C92_n1072, mult_28_C92_n1071, 
      mult_28_C92_n1070, mult_28_C92_n1069, mult_28_C92_n1068, 
      mult_28_C92_n1067, mult_28_C92_n1066, mult_28_C92_n1065, 
      mult_28_C92_n1064, mult_28_C92_n1063, mult_28_C92_n1062, 
      mult_28_C92_n1061, mult_28_C92_n1060, mult_28_C92_n1059, 
      mult_28_C92_n1058, mult_28_C92_n1057, mult_28_C92_n1056, 
      mult_28_C92_n1055, mult_28_C92_n1054, mult_28_C92_n1053, 
      mult_28_C92_n1052, mult_28_C92_n1051, mult_28_C92_n1050, 
      mult_28_C92_n1049, mult_28_C92_n1048, mult_28_C92_n1047, 
      mult_28_C92_n1046, mult_28_C92_n1045, mult_28_C92_n1044, 
      mult_28_C92_n1043, mult_28_C92_n1042, mult_28_C92_n1041, 
      mult_28_C92_n1040, mult_28_C92_n1039, mult_28_C92_n1038, 
      mult_28_C92_n1037, mult_28_C92_n1036, mult_28_C92_n1035, 
      mult_28_C92_n1034, mult_28_C92_n1033, mult_28_C92_n1032, 
      mult_28_C92_n1031, mult_28_C92_n1030, mult_28_C92_n1029, 
      mult_28_C92_n1028, mult_28_C92_n1027, mult_28_C92_n1026, 
      mult_28_C92_n1025, mult_28_C92_n1024, mult_28_C92_n1023, 
      mult_28_C92_n1022, mult_28_C92_n1021, mult_28_C92_n1020, 
      mult_28_C92_n1019, mult_28_C92_n1018, mult_28_C92_n1017, 
      mult_28_C92_n1016, mult_28_C92_n1015, mult_28_C92_n1014, 
      mult_28_C92_n1013, mult_28_C92_n1012, mult_28_C92_n1011, 
      mult_28_C92_n1010, mult_28_C92_n1009, mult_28_C92_n1008, 
      mult_28_C92_n1007, mult_28_C92_n1006, mult_28_C92_n1005, 
      mult_28_C92_n1004, mult_28_C92_n1003, mult_28_C92_n1002, 
      mult_28_C92_n1001, mult_28_C92_n1000, mult_28_C92_n999, mult_28_C92_n998,
      mult_28_C92_n997, mult_28_C92_n996, mult_28_C92_n995, mult_28_C92_n994, 
      mult_28_C92_n993, mult_28_C92_n992, mult_28_C92_n991, mult_28_C92_n990, 
      mult_28_C92_n989, mult_28_C92_n988, mult_28_C92_n987, mult_28_C92_n986, 
      mult_28_C92_n985, mult_28_C92_n984, mult_28_C92_n983, mult_28_C92_n982, 
      mult_28_C92_n981, mult_28_C92_n980, mult_28_C92_n979, mult_28_C92_n978, 
      mult_28_C92_n977, mult_28_C92_n976, mult_28_C92_n975, mult_28_C92_n974, 
      mult_28_C92_n973, mult_28_C92_n972, mult_28_C92_n971, mult_28_C92_n970, 
      mult_28_C92_n969, mult_28_C92_n968, mult_28_C92_n967, mult_28_C92_n966, 
      mult_28_C92_n965, mult_28_C92_n964, mult_28_C92_n963, mult_28_C92_n962, 
      mult_28_C92_n961, mult_28_C92_n960, mult_28_C92_n959, mult_28_C92_n958, 
      mult_28_C92_n957, mult_28_C92_n956, mult_28_C92_n955, mult_28_C92_n954, 
      mult_28_C92_n953, mult_28_C92_n952, mult_28_C92_n951, mult_28_C92_n950, 
      mult_28_C92_n949, mult_28_C92_n948, mult_28_C92_n947, mult_28_C92_n946, 
      mult_28_C92_n945, mult_28_C92_n944, mult_28_C92_n943, mult_28_C92_n942, 
      mult_28_C92_n941, mult_28_C92_n940, mult_28_C92_n939, mult_28_C92_n938, 
      mult_28_C92_n937, mult_28_C92_n936, mult_28_C92_n935, mult_28_C92_n934, 
      mult_28_C92_n933, mult_28_C92_n932, mult_28_C92_n931, mult_28_C92_n930, 
      mult_28_C92_n929, mult_28_C92_n928, mult_28_C92_n927, mult_28_C92_n926, 
      mult_28_C92_n925, mult_28_C92_n924, mult_28_C92_n923, mult_28_C92_n922, 
      mult_28_C92_n921, mult_28_C92_n920, mult_28_C92_n919, mult_28_C92_n918, 
      mult_28_C92_n917, mult_28_C92_n916, mult_28_C92_n915, mult_28_C92_n914, 
      mult_28_C92_n913, mult_28_C92_n912, mult_28_C92_n911, mult_28_C92_n910, 
      mult_28_C92_n464, mult_28_C92_n473, mult_28_C92_net11020, 
      mult_28_C92_net11797, mult_28_C92_net11803, mult_28_C92_n466, 
      mult_28_C92_n470, mult_28_C92_n472, mult_28_C92_n477, mult_28_C92_n478, 
      mult_28_C92_n481, mult_28_C92_n482, mult_28_C92_n525, mult_28_C92_n591, 
      mult_28_C92_n605, mult_28_C92_n633, mult_28_C92_n709, 
      mult_28_C92_net11337, mult_28_C92_n230, mult_28_C92_n231, 
      mult_28_C92_n233, mult_28_C92_n235, mult_28_C92_n243, mult_28_C92_n248, 
      mult_28_C92_n250, mult_28_C92_n261, mult_28_C92_n266, mult_28_C92_n268, 
      mult_28_C92_n269, mult_28_C92_n483, mult_28_C92_n484, 
      mult_28_C92_net12275, mult_28_C92_n576, mult_28_C92_n604, 
      mult_28_C92_n632, mult_28_C92_n767, mult_28_C92_net11996, 
      mult_28_C92_n174, mult_28_C92_n175, mult_28_C92_n176, mult_28_C92_n178, 
      mult_28_C92_n179, mult_28_C92_n180, mult_28_C92_n183, mult_28_C92_n184, 
      mult_28_C92_n185, mult_28_C92_n199, mult_28_C92_n294, mult_28_C92_n295, 
      mult_28_C92_n63, mult_28_C92_net12274, mult_28_C92_n468, mult_28_C92_n475
      , mult_28_C92_net11941, mult_28_C92_net12148, mult_28_C92_n217, 
      mult_28_C92_n218, mult_28_C92_n219, mult_28_C92_n221, mult_28_C92_n451, 
      mult_28_C92_n452, mult_28_C92_n455, mult_28_C92_n456, mult_28_C92_n465, 
      mult_28_C92_n469, mult_28_C92_net11961, mult_28_C92_net11981, 
      mult_28_C92_net11982, mult_28_C92_net9967, mult_28_C92_net9968, 
      mult_28_C92_net9969, mult_28_C92_net9971, mult_28_C92_net9972, 
      mult_28_C92_net9974, mult_28_C92_net9975, mult_28_C92_net9976, 
      mult_28_C92_n211, mult_28_C92_n212, mult_28_C92_n213, mult_28_C92_n214, 
      mult_28_C92_n300, mult_28_C92_n186, mult_28_C92_n187, mult_28_C92_n191, 
      mult_28_C92_n194, mult_28_C92_n196, mult_28_C92_n197, mult_28_C92_n206, 
      mult_28_C92_n737, mult_28_C92_net11920, mult_28_C92_net12350, 
      mult_28_C92_net12321, mult_28_C92_net12315, mult_28_C92_net12273, 
      mult_28_C92_net12262, mult_28_C92_net12187, mult_28_C92_net12184, 
      mult_28_C92_net12160, mult_28_C92_net12114, mult_28_C92_net12088, 
      mult_28_C92_net12005, mult_28_C92_net11946, mult_28_C92_net11942, 
      mult_28_C92_net11943, mult_28_C92_net11944, mult_28_C92_net11792, 
      mult_28_C92_net11686, mult_28_C92_net11523, mult_28_C92_net11524, 
      mult_28_C92_net11339, mult_28_C92_net11247, mult_28_C92_net11021, 
      mult_28_C92_net10923, mult_28_C92_net10919, mult_28_C92_net9959, 
      mult_28_C92_net9957, mult_28_C92_n842, mult_28_C92_n835, mult_28_C92_n834
      , mult_28_C92_n814, mult_28_C92_n812, mult_28_C92_n811, mult_28_C92_n794,
      mult_28_C92_n793, mult_28_C92_n792, mult_28_C92_n791, mult_28_C92_n790, 
      mult_28_C92_n789, mult_28_C92_n788, mult_28_C92_n787, mult_28_C92_n786, 
      mult_28_C92_n785, mult_28_C92_n784, mult_28_C92_n783, mult_28_C92_n782, 
      mult_28_C92_n781, mult_28_C92_n780, mult_28_C92_n779, mult_28_C92_n778, 
      mult_28_C92_n777, mult_28_C92_n776, mult_28_C92_n775, mult_28_C92_n774, 
      mult_28_C92_n773, mult_28_C92_n772, mult_28_C92_n771, mult_28_C92_n770, 
      mult_28_C92_n769, mult_28_C92_n768, mult_28_C92_n766, mult_28_C92_n765, 
      mult_28_C92_n764, mult_28_C92_n763, mult_28_C92_n762, mult_28_C92_n761, 
      mult_28_C92_n760, mult_28_C92_n759, mult_28_C92_n758, mult_28_C92_n757, 
      mult_28_C92_n756, mult_28_C92_n755, mult_28_C92_n754, mult_28_C92_n753, 
      mult_28_C92_n752, mult_28_C92_n751, mult_28_C92_n750, mult_28_C92_n749, 
      mult_28_C92_n748, mult_28_C92_n747, mult_28_C92_n746, mult_28_C92_n745, 
      mult_28_C92_n744, mult_28_C92_n743, mult_28_C92_n742, mult_28_C92_n741, 
      mult_28_C92_n740, mult_28_C92_n739, mult_28_C92_n738, mult_28_C92_n736, 
      mult_28_C92_n735, mult_28_C92_n734, mult_28_C92_n733, mult_28_C92_n732, 
      mult_28_C92_n731, mult_28_C92_n730, mult_28_C92_n729, mult_28_C92_n728, 
      mult_28_C92_n727, mult_28_C92_n726, mult_28_C92_n725, mult_28_C92_n724, 
      mult_28_C92_n723, mult_28_C92_n722, mult_28_C92_n721, mult_28_C92_n720, 
      mult_28_C92_n719, mult_28_C92_n718, mult_28_C92_n717, mult_28_C92_n716, 
      mult_28_C92_n715, mult_28_C92_n714, mult_28_C92_n713, mult_28_C92_n712, 
      mult_28_C92_n711, mult_28_C92_n710, mult_28_C92_n708, mult_28_C92_n707, 
      mult_28_C92_n706, mult_28_C92_n705, mult_28_C92_n704, mult_28_C92_n703, 
      mult_28_C92_n702, mult_28_C92_n701, mult_28_C92_n700, mult_28_C92_n699, 
      mult_28_C92_n698, mult_28_C92_n697, mult_28_C92_n696, mult_28_C92_n695, 
      mult_28_C92_n694, mult_28_C92_n693, mult_28_C92_n692, mult_28_C92_n691, 
      mult_28_C92_n690, mult_28_C92_n689, mult_28_C92_n688, mult_28_C92_n687, 
      mult_28_C92_n686, mult_28_C92_n685, mult_28_C92_n684, mult_28_C92_n683, 
      mult_28_C92_n682, mult_28_C92_n681, mult_28_C92_n680, mult_28_C92_n679, 
      mult_28_C92_n678, mult_28_C92_n677, mult_28_C92_n676, mult_28_C92_n675, 
      mult_28_C92_n674, mult_28_C92_n673, mult_28_C92_n672, mult_28_C92_n671, 
      mult_28_C92_n670, mult_28_C92_n669, mult_28_C92_n668, mult_28_C92_n667, 
      mult_28_C92_n666, mult_28_C92_n665, mult_28_C92_n664, mult_28_C92_n663, 
      mult_28_C92_n662, mult_28_C92_n661, mult_28_C92_n660, mult_28_C92_n659, 
      mult_28_C92_n658, mult_28_C92_n657, mult_28_C92_n656, mult_28_C92_n655, 
      mult_28_C92_n654, mult_28_C92_n653, mult_28_C92_n652, mult_28_C92_n651, 
      mult_28_C92_n650, mult_28_C92_n649, mult_28_C92_n648, mult_28_C92_n647, 
      mult_28_C92_n646, mult_28_C92_n645, mult_28_C92_n644, mult_28_C92_n643, 
      mult_28_C92_n642, mult_28_C92_n641, mult_28_C92_n640, mult_28_C92_n639, 
      mult_28_C92_n638, mult_28_C92_n637, mult_28_C92_n636, mult_28_C92_n635, 
      mult_28_C92_n634, mult_28_C92_n631, mult_28_C92_n630, mult_28_C92_n629, 
      mult_28_C92_n628, mult_28_C92_n627, mult_28_C92_n626, mult_28_C92_n625, 
      mult_28_C92_n624, mult_28_C92_n623, mult_28_C92_n622, mult_28_C92_n621, 
      mult_28_C92_n620, mult_28_C92_n619, mult_28_C92_n618, mult_28_C92_n617, 
      mult_28_C92_n616, mult_28_C92_n615, mult_28_C92_n614, mult_28_C92_n613, 
      mult_28_C92_n612, mult_28_C92_n611, mult_28_C92_n610, mult_28_C92_n609, 
      mult_28_C92_n608, mult_28_C92_n607, mult_28_C92_n606, mult_28_C92_n603, 
      mult_28_C92_n602, mult_28_C92_n601, mult_28_C92_n600, mult_28_C92_n599, 
      mult_28_C92_n598, mult_28_C92_n597, mult_28_C92_n596, mult_28_C92_n595, 
      mult_28_C92_n594, mult_28_C92_n593, mult_28_C92_n592, mult_28_C92_n590, 
      mult_28_C92_n589, mult_28_C92_n588, mult_28_C92_n587, mult_28_C92_n586, 
      mult_28_C92_n585, mult_28_C92_n584, mult_28_C92_n583, mult_28_C92_n582, 
      mult_28_C92_n581, mult_28_C92_n580, mult_28_C92_n579, mult_28_C92_n578, 
      mult_28_C92_n577, mult_28_C92_n574, mult_28_C92_n573, mult_28_C92_n572, 
      mult_28_C92_n571, mult_28_C92_n570, mult_28_C92_n569, mult_28_C92_n568, 
      mult_28_C92_n567, mult_28_C92_n566, mult_28_C92_n565, mult_28_C92_n564, 
      mult_28_C92_n563, mult_28_C92_n562, mult_28_C92_n561, mult_28_C92_n560, 
      mult_28_C92_n559, mult_28_C92_n558, mult_28_C92_n557, mult_28_C92_n556, 
      mult_28_C92_n555, mult_28_C92_n554, mult_28_C92_n553, mult_28_C92_n552, 
      mult_28_C92_n551, mult_28_C92_n550, mult_28_C92_n549, mult_28_C92_n548, 
      mult_28_C92_n547, mult_28_C92_n546, mult_28_C92_n545, mult_28_C92_n544, 
      mult_28_C92_n543, mult_28_C92_n542, mult_28_C92_n541, mult_28_C92_n540, 
      mult_28_C92_n539, mult_28_C92_n538, mult_28_C92_n537, mult_28_C92_n536, 
      mult_28_C92_n535, mult_28_C92_n534, mult_28_C92_n533, mult_28_C92_n532, 
      mult_28_C92_n530, mult_28_C92_n529, mult_28_C92_n528, mult_28_C92_n527, 
      mult_28_C92_n526, mult_28_C92_n524, mult_28_C92_n523, mult_28_C92_n522, 
      mult_28_C92_n521, mult_28_C92_n520, mult_28_C92_n519, mult_28_C92_n518, 
      mult_28_C92_n517, mult_28_C92_n516, mult_28_C92_n515, mult_28_C92_n514, 
      mult_28_C92_n513, mult_28_C92_n512, mult_28_C92_n511, mult_28_C92_n510, 
      mult_28_C92_n509, mult_28_C92_n508, mult_28_C92_n507, mult_28_C92_n506, 
      mult_28_C92_n505, mult_28_C92_n504, mult_28_C92_n503, mult_28_C92_n502, 
      mult_28_C92_n501, mult_28_C92_n500, mult_28_C92_n499, mult_28_C92_n498, 
      mult_28_C92_n497, mult_28_C92_n496, mult_28_C92_n495, mult_28_C92_n494, 
      mult_28_C92_n493, mult_28_C92_n492, mult_28_C92_n491, mult_28_C92_n490, 
      mult_28_C92_n489, mult_28_C92_n488, mult_28_C92_n487, mult_28_C92_n486, 
      mult_28_C92_n485, mult_28_C92_n480, mult_28_C92_n479, mult_28_C92_n476, 
      mult_28_C92_n474, mult_28_C92_n471, mult_28_C92_n467, mult_28_C92_n463, 
      mult_28_C92_n462, mult_28_C92_n460, mult_28_C92_n459, mult_28_C92_n458, 
      mult_28_C92_n457, mult_28_C92_n454, mult_28_C92_n453, mult_28_C92_n450, 
      mult_28_C92_n449, mult_28_C92_n448, mult_28_C92_n447, mult_28_C92_n446, 
      mult_28_C92_n445, mult_28_C92_n444, mult_28_C92_n443, mult_28_C92_n442, 
      mult_28_C92_n441, mult_28_C92_n440, mult_28_C92_n439, mult_28_C92_n438, 
      mult_28_C92_n437, mult_28_C92_n436, mult_28_C92_n435, mult_28_C92_n434, 
      mult_28_C92_n433, mult_28_C92_n432, mult_28_C92_n431, mult_28_C92_n430, 
      mult_28_C92_n429, mult_28_C92_n428, mult_28_C92_n427, mult_28_C92_n426, 
      mult_28_C92_n425, mult_28_C92_n424, mult_28_C92_n423, mult_28_C92_n422, 
      mult_28_C92_n421, mult_28_C92_n420, mult_28_C92_n419, mult_28_C92_n418, 
      mult_28_C92_n417, mult_28_C92_n416, mult_28_C92_n415, mult_28_C92_n414, 
      mult_28_C92_n413, mult_28_C92_n412, mult_28_C92_n411, mult_28_C92_n410, 
      mult_28_C92_n409, mult_28_C92_n408, mult_28_C92_n407, mult_28_C92_n406, 
      mult_28_C92_n405, mult_28_C92_n404, mult_28_C92_n403, mult_28_C92_n402, 
      mult_28_C92_n401, mult_28_C92_n400, mult_28_C92_n399, mult_28_C92_n398, 
      mult_28_C92_n397, mult_28_C92_n396, mult_28_C92_n395, mult_28_C92_n394, 
      mult_28_C92_n393, mult_28_C92_n392, mult_28_C92_n391, mult_28_C92_n390, 
      mult_28_C92_n389, mult_28_C92_n388, mult_28_C92_n387, mult_28_C92_n386, 
      mult_28_C92_n385, mult_28_C92_n384, mult_28_C92_n383, mult_28_C92_n382, 
      mult_28_C92_n381, mult_28_C92_n380, mult_28_C92_n379, mult_28_C92_n378, 
      mult_28_C92_n377, mult_28_C92_n376, mult_28_C92_n375, mult_28_C92_n374, 
      mult_28_C92_n373, mult_28_C92_n372, mult_28_C92_n371, mult_28_C92_n370, 
      mult_28_C92_n369, mult_28_C92_n368, mult_28_C92_n367, mult_28_C92_n366, 
      mult_28_C92_n365, mult_28_C92_n364, mult_28_C92_n363, mult_28_C92_n362, 
      mult_28_C92_n361, mult_28_C92_n360, mult_28_C92_n359, mult_28_C92_n358, 
      mult_28_C92_n357, mult_28_C92_n356, mult_28_C92_n355, mult_28_C92_n354, 
      mult_28_C92_n353, mult_28_C92_n352, mult_28_C92_n351, mult_28_C92_n350, 
      mult_28_C92_n349, mult_28_C92_n348, mult_28_C92_n347, mult_28_C92_n346, 
      mult_28_C92_n345, mult_28_C92_n344, mult_28_C92_n343, mult_28_C92_n342, 
      mult_28_C92_n341, mult_28_C92_n340, mult_28_C92_n339, mult_28_C92_n338, 
      mult_28_C92_n337, mult_28_C92_n336, mult_28_C92_n335, mult_28_C92_n334, 
      mult_28_C92_n333, mult_28_C92_n332, mult_28_C92_n331, mult_28_C92_n330, 
      mult_28_C92_n329, mult_28_C92_n328, mult_28_C92_n327, mult_28_C92_n326, 
      mult_28_C92_n325, mult_28_C92_n324, mult_28_C92_n323, mult_28_C92_n322, 
      mult_28_C92_n321, mult_28_C92_n320, mult_28_C92_n319, mult_28_C92_n318, 
      mult_28_C92_n317, mult_28_C92_n316, mult_28_C92_n315, mult_28_C92_n299, 
      mult_28_C92_n298, mult_28_C92_n297, mult_28_C92_n296, mult_28_C92_n293, 
      mult_28_C92_n290, mult_28_C92_n289, mult_28_C92_n288, mult_28_C92_n287, 
      mult_28_C92_n277, mult_28_C92_n276, mult_28_C92_n275, mult_28_C92_n274, 
      mult_28_C92_n267, mult_28_C92_n220, mult_28_C92_n216, mult_28_C92_n215, 
      mult_28_C92_n208, mult_28_C92_n207, mult_28_C92_n204, mult_28_C92_n203, 
      mult_28_C92_n202, mult_28_C92_n195, mult_28_C92_n190, mult_28_C92_n189, 
      mult_28_C92_n188, mult_28_C92_n171, mult_28_C92_n170, mult_28_C92_n169, 
      mult_28_C92_n168, mult_28_C92_n167, mult_28_C92_n164, mult_28_C92_n162, 
      mult_28_C92_n161, mult_28_C92_n160, mult_28_C92_n159, mult_28_C92_n158, 
      mult_28_C92_n157, mult_28_C92_n155, mult_28_C92_n151, mult_28_C92_n150, 
      mult_28_C92_n149, mult_28_C92_n148, mult_28_C92_n147, mult_28_C92_n146, 
      mult_28_C92_n142, mult_28_C92_n141, mult_28_C92_n140, mult_28_C92_n139, 
      mult_28_C92_n136, mult_28_C92_n135, mult_28_C92_n134, mult_28_C92_n133, 
      mult_28_C92_n130, mult_28_C92_n129, mult_28_C92_n128, mult_28_C92_n127, 
      mult_28_C92_n126, mult_28_C92_n125, mult_28_C92_n120, mult_28_C92_n119, 
      mult_28_C92_n118, mult_28_C92_n117, mult_28_C92_n116, mult_28_C92_n115, 
      mult_28_C92_n114, mult_28_C92_n113, mult_28_C92_n112, mult_28_C92_n109, 
      mult_28_C92_n108, mult_28_C92_n107, mult_28_C92_n106, mult_28_C92_n105, 
      mult_28_C92_n104, mult_28_C92_n103, mult_28_C92_n102, mult_28_C92_n101, 
      mult_28_C92_n100, mult_28_C92_n97, mult_28_C92_n96, mult_28_C92_n95, 
      mult_28_C92_n94, mult_28_C92_n93, mult_28_C92_n92, mult_28_C92_n87, 
      mult_28_C92_n86, mult_28_C92_n85, mult_28_C92_n84, mult_28_C92_n69, 
      mult_28_C92_n64, mult_28_C92_n62, mult_28_C92_n61, mult_28_C92_n60, 
      mult_28_C92_n57, mult_28_C92_n55, mult_28_C92_n54, mult_28_C92_n53, 
      mult_28_C92_n52, mult_28_C92_n48, mult_28_C92_n46, mult_28_C92_n42, 
      mult_28_C92_n40, mult_28_C92_n36, mult_28_C92_n34, mult_28_C92_n30, 
      mult_28_C92_n28, mult_28_C92_n24, mult_28_C92_n22, mult_28_C92_n18, 
      mult_28_C92_n16, mult_28_C92_n12, mult_28_C92_n9, mult_28_C92_n6, 
      add_102_n202, add_102_n201, add_102_n200, add_102_n199, add_102_n198, 
      add_102_n197, add_102_n196, add_102_n195, add_102_n194, add_102_n193, 
      add_102_n192, add_102_n191, add_102_n190, add_102_n189, add_102_n188, 
      add_102_n187, add_102_n123, add_102_n65, add_102_n67, add_102_n72, 
      add_102_n83, add_102_n122, add_102_n61, add_102_n62, add_102_n63, 
      add_102_n64, add_102_n66, add_102_n70, add_102_n73, add_102_n75, 
      add_102_n79, add_102_n8, add_102_n84, add_102_n86, add_102_n87, 
      add_102_n88, add_102_net11440, add_102_net11486, add_102_net12276, 
      add_102_n60, add_102_n78, add_102_net12241, add_102_net12242, 
      add_102_net11859, add_102_net11615, add_102_net11439, add_102_net11441, 
      add_102_net11329, add_102_n129, add_102_n120, add_102_n119, add_102_n118,
      add_102_n117, add_102_n115, add_102_n113, add_102_n112, add_102_n108, 
      add_102_n107, add_102_n106, add_102_n105, add_102_n104, add_102_n102, 
      add_102_n101, add_102_n100, add_102_n98, add_102_n97, add_102_n96, 
      add_102_n95, add_102_n94, add_102_n93, add_102_n92, add_102_n91, 
      add_102_n90, add_102_n89, add_102_n82, add_102_n81, add_102_n80, 
      add_102_n71, add_102_n59, add_102_n58, add_102_n56, add_102_n55, 
      add_102_n53, add_102_n52, add_102_n51, add_102_n50, add_102_n47, 
      add_102_n45, add_102_n44, add_102_n43, add_102_n42, add_102_n39, 
      add_102_n38, add_102_n37, add_102_n36, add_102_n35, add_102_n34, 
      add_102_n33, add_102_n32, add_102_n31, add_102_n30, add_102_n28, 
      add_102_n27, add_102_n26, add_102_n23, add_102_n22, add_102_n21, 
      add_102_n20, add_102_n19, add_102_n17, add_102_n16, add_102_n15, 
      add_102_n14, add_102_n13, add_102_n12, add_102_n10, add_102_n9, 
      add_102_n7, add_102_n6, add_102_n5, add_102_n4, add_102_n3, add_102_n2, 
      add_102_n1, add_0_root_add_0_root_add_101_n201, 
      add_0_root_add_0_root_add_101_n199, add_0_root_add_0_root_add_101_n198, 
      add_0_root_add_0_root_add_101_n197, add_0_root_add_0_root_add_101_n196, 
      add_0_root_add_0_root_add_101_n195, add_0_root_add_0_root_add_101_n194, 
      add_0_root_add_0_root_add_101_n193, add_0_root_add_0_root_add_101_n192, 
      add_0_root_add_0_root_add_101_n191, add_0_root_add_0_root_add_101_n190, 
      add_0_root_add_0_root_add_101_n189, add_0_root_add_0_root_add_101_n188, 
      add_0_root_add_0_root_add_101_n187, add_0_root_add_0_root_add_101_n186, 
      add_0_root_add_0_root_add_101_n185, add_0_root_add_0_root_add_101_n184, 
      add_0_root_add_0_root_add_101_n183, add_0_root_add_0_root_add_101_n182, 
      add_0_root_add_0_root_add_101_n181, add_0_root_add_0_root_add_101_n180, 
      add_0_root_add_0_root_add_101_n179, add_0_root_add_0_root_add_101_n1, 
      add_0_root_add_0_root_add_101_n109, add_0_root_add_0_root_add_101_n19, 
      add_0_root_add_0_root_add_101_n20, add_0_root_add_0_root_add_101_n21, 
      add_0_root_add_0_root_add_101_n22, add_0_root_add_0_root_add_101_n23, 
      add_0_root_add_0_root_add_101_n26, add_0_root_add_0_root_add_101_n30, 
      add_0_root_add_0_root_add_101_n31, add_0_root_add_0_root_add_101_n32, 
      add_0_root_add_0_root_add_101_n33, add_0_root_add_0_root_add_101_n38, 
      add_0_root_add_0_root_add_101_n58, add_0_root_add_0_root_add_101_n59, 
      add_0_root_add_0_root_add_101_net11559, 
      add_0_root_add_0_root_add_101_net11588, add_0_root_add_0_root_add_101_n60
      , add_0_root_add_0_root_add_101_n61, add_0_root_add_0_root_add_101_n62, 
      add_0_root_add_0_root_add_101_n63, add_0_root_add_0_root_add_101_n67, 
      add_0_root_add_0_root_add_101_n72, add_0_root_add_0_root_add_101_n37, 
      add_0_root_add_0_root_add_101_n116, add_0_root_add_0_root_add_101_n73, 
      add_0_root_add_0_root_add_101_n87, add_0_root_add_0_root_add_101_n88, 
      add_0_root_add_0_root_add_101_net12354, 
      add_0_root_add_0_root_add_101_net12355, 
      add_0_root_add_0_root_add_101_net12169, 
      add_0_root_add_0_root_add_101_net12025, 
      add_0_root_add_0_root_add_101_net11959, 
      add_0_root_add_0_root_add_101_net9993, add_0_root_add_0_root_add_101_n107
      , add_0_root_add_0_root_add_101_n105, add_0_root_add_0_root_add_101_n104,
      add_0_root_add_0_root_add_101_n103, add_0_root_add_0_root_add_101_n102, 
      add_0_root_add_0_root_add_101_n100, add_0_root_add_0_root_add_101_n98, 
      add_0_root_add_0_root_add_101_n97, add_0_root_add_0_root_add_101_n96, 
      add_0_root_add_0_root_add_101_n95, add_0_root_add_0_root_add_101_n94, 
      add_0_root_add_0_root_add_101_n93, add_0_root_add_0_root_add_101_n92, 
      add_0_root_add_0_root_add_101_n91, add_0_root_add_0_root_add_101_n90, 
      add_0_root_add_0_root_add_101_n89, add_0_root_add_0_root_add_101_n85, 
      add_0_root_add_0_root_add_101_n84, add_0_root_add_0_root_add_101_n83, 
      add_0_root_add_0_root_add_101_n82, add_0_root_add_0_root_add_101_n81, 
      add_0_root_add_0_root_add_101_n80, add_0_root_add_0_root_add_101_n79, 
      add_0_root_add_0_root_add_101_n78, add_0_root_add_0_root_add_101_n75, 
      add_0_root_add_0_root_add_101_n71, add_0_root_add_0_root_add_101_n70, 
      add_0_root_add_0_root_add_101_n66, add_0_root_add_0_root_add_101_n65, 
      add_0_root_add_0_root_add_101_n56, add_0_root_add_0_root_add_101_n55, 
      add_0_root_add_0_root_add_101_n54, add_0_root_add_0_root_add_101_n53, 
      add_0_root_add_0_root_add_101_n52, add_0_root_add_0_root_add_101_n51, 
      add_0_root_add_0_root_add_101_n50, add_0_root_add_0_root_add_101_n45, 
      add_0_root_add_0_root_add_101_n44, add_0_root_add_0_root_add_101_n43, 
      add_0_root_add_0_root_add_101_n42, add_0_root_add_0_root_add_101_n39, 
      add_0_root_add_0_root_add_101_n36, add_0_root_add_0_root_add_101_n35, 
      add_0_root_add_0_root_add_101_n34, add_0_root_add_0_root_add_101_n29, 
      add_0_root_add_0_root_add_101_n28, add_0_root_add_0_root_add_101_n27, 
      add_0_root_add_0_root_add_101_n16, add_0_root_add_0_root_add_101_n15, 
      add_0_root_add_0_root_add_101_n14, add_0_root_add_0_root_add_101_n13, 
      add_0_root_add_0_root_add_101_n12, add_0_root_add_0_root_add_101_n9, 
      add_0_root_add_0_root_add_101_n8, add_0_root_add_0_root_add_101_n7, 
      add_0_root_add_0_root_add_101_n6, add_0_root_add_0_root_add_101_n5, 
      add_0_root_add_0_root_add_101_n4, add_99_n209, add_99_n208, add_99_n207, 
      add_99_n206, add_99_n205, add_99_n203, add_99_n202, add_99_n201, 
      add_99_n200, add_99_n199, add_99_n198, add_99_n197, add_99_n196, 
      add_99_n195, add_99_n194, add_99_n193, add_99_n192, add_99_n191, 
      add_99_n190, add_99_n189, add_99_n188, add_99_n187, add_99_n186, 
      add_99_n185, add_99_n184, add_99_n183, add_99_n182, add_99_n181, 
      add_99_n180, add_99_n179, add_99_n116, add_99_n112, add_99_n110, 
      add_99_n109, add_99_n107, add_99_n105, add_99_n104, add_99_n103, 
      add_99_n102, add_99_n98, add_99_n97, add_99_n96, add_99_n95, add_99_n94, 
      add_99_n93, add_99_n92, add_99_n91, add_99_n90, add_99_n89, add_99_n88, 
      add_99_n87, add_99_n86, add_99_n85, add_99_n84, add_99_n83, add_99_n82, 
      add_99_n81, add_99_n80, add_99_n79, add_99_n78, add_99_n75, add_99_n73, 
      add_99_n72, add_99_n71, add_99_n70, add_99_n67, add_99_n66, add_99_n65, 
      add_99_n64, add_99_n63, add_99_n62, add_99_n61, add_99_n60, add_99_n59, 
      add_99_n58, add_99_n56, add_99_n55, add_99_n53, add_99_n52, add_99_n51, 
      add_99_n50, add_99_n47, add_99_n45, add_99_n44, add_99_n43, add_99_n42, 
      add_99_n39, add_99_n38, add_99_n37, add_99_n36, add_99_n35, add_99_n34, 
      add_99_n33, add_99_n32, add_99_n31, add_99_n30, add_99_n29, add_99_n28, 
      add_99_n27, add_99_n26, add_99_n23, add_99_n22, add_99_n21, add_99_n20, 
      add_99_n19, add_99_n16, add_99_n15, add_99_n14, add_99_n13, add_99_n12, 
      add_99_n11, add_99_n10, add_99_n9, add_99_n8, add_99_n5, add_99_n1, 
      mult_28_C95_n_1033, mult_28_C95_n1013, mult_28_C95_n1012, 
      mult_28_C95_n1011, mult_28_C95_n1010, mult_28_C95_n1009, 
      mult_28_C95_n1008, mult_28_C95_n1007, mult_28_C95_n1006, 
      mult_28_C95_n1005, mult_28_C95_n1004, mult_28_C95_n1003, 
      mult_28_C95_n1002, mult_28_C95_n1001, mult_28_C95_n1000, mult_28_C95_n999
      , mult_28_C95_n998, mult_28_C95_n997, mult_28_C95_n996, mult_28_C95_n995,
      mult_28_C95_n994, mult_28_C95_n993, mult_28_C95_n992, mult_28_C95_n991, 
      mult_28_C95_n990, mult_28_C95_n989, mult_28_C95_n988, mult_28_C95_n987, 
      mult_28_C95_n986, mult_28_C95_n985, mult_28_C95_n984, mult_28_C95_n983, 
      mult_28_C95_n982, mult_28_C95_n981, mult_28_C95_n980, mult_28_C95_n979, 
      mult_28_C95_n978, mult_28_C95_n977, mult_28_C95_n976, mult_28_C95_n975, 
      mult_28_C95_n974, mult_28_C95_n973, mult_28_C95_n972, mult_28_C95_n971, 
      mult_28_C95_n970, mult_28_C95_n969, mult_28_C95_n968, mult_28_C95_n967, 
      mult_28_C95_n966, mult_28_C95_n965, mult_28_C95_n964, mult_28_C95_n963, 
      mult_28_C95_n962, mult_28_C95_n961, mult_28_C95_n960, mult_28_C95_n959, 
      mult_28_C95_n958, mult_28_C95_n957, mult_28_C95_n956, mult_28_C95_n955, 
      mult_28_C95_n954, mult_28_C95_n953, mult_28_C95_n952, mult_28_C95_n951, 
      mult_28_C95_n950, mult_28_C95_n949, mult_28_C95_n948, mult_28_C95_n947, 
      mult_28_C95_n946, mult_28_C95_n945, mult_28_C95_n944, mult_28_C95_n943, 
      mult_28_C95_n942, mult_28_C95_n941, mult_28_C95_n940, mult_28_C95_n939, 
      mult_28_C95_n938, mult_28_C95_n937, mult_28_C95_n936, mult_28_C95_n935, 
      mult_28_C95_n934, mult_28_C95_n933, mult_28_C95_n932, mult_28_C95_n931, 
      mult_28_C95_n930, mult_28_C95_n929, mult_28_C95_n928, mult_28_C95_n927, 
      mult_28_C95_n926, mult_28_C95_n925, mult_28_C95_n924, mult_28_C95_n923, 
      mult_28_C95_n922, mult_28_C95_n921, mult_28_C95_n920, mult_28_C95_n919, 
      mult_28_C95_n918, mult_28_C95_n917, mult_28_C95_n916, mult_28_C95_n915, 
      mult_28_C95_n914, mult_28_C95_n913, mult_28_C95_n912, mult_28_C95_n911, 
      mult_28_C95_n910, mult_28_C95_n909, mult_28_C95_n908, mult_28_C95_n907, 
      mult_28_C95_n906, mult_28_C95_n905, mult_28_C95_n904, mult_28_C95_n903, 
      mult_28_C95_n902, mult_28_C95_n901, mult_28_C95_n900, mult_28_C95_n706, 
      mult_28_C95_n175, mult_28_C95_n176, mult_28_C95_n177, mult_28_C95_n178, 
      mult_28_C95_n189, mult_28_C95_n134, mult_28_C95_n143, mult_28_C95_n144, 
      mult_28_C95_n150, mult_28_C95_n151, mult_28_C95_n152, mult_28_C95_n153, 
      mult_28_C95_n154, mult_28_C95_n155, mult_28_C95_n162, mult_28_C95_n163, 
      mult_28_C95_n164, mult_28_C95_n282, mult_28_C95_net10037, 
      mult_28_C95_net11096, mult_28_C95_net11621, mult_28_C95_net11675, 
      mult_28_C95_n179, mult_28_C95_n184, mult_28_C95_n375, mult_28_C95_n376, 
      mult_28_C95_net12019, mult_28_C95_n389, mult_28_C95_n390, 
      mult_28_C95_n405, mult_28_C95_n406, mult_28_C95_n421, mult_28_C95_n423, 
      mult_28_C95_n424, mult_28_C95_n439, mult_28_C95_n440, mult_28_C95_n545, 
      mult_28_C95_n589, mult_28_C95_n633, mult_28_C95_n634, mult_28_C95_n391, 
      mult_28_C95_n392, mult_28_C95_n395, mult_28_C95_n396, mult_28_C95_n409, 
      mult_28_C95_n411, mult_28_C95_n412, mult_28_C95_n414, mult_28_C95_n543, 
      mult_28_C95_n557, mult_28_C95_n558, mult_28_C95_n572, mult_28_C95_n617, 
      mult_28_C95_n692, mult_28_C95_n693, mult_28_C95_n707, mult_28_C95_n803, 
      mult_28_C95_n677, mult_28_C95_n678, mult_28_C95_n802, mult_28_C95_n387, 
      mult_28_C95_net11585, mult_28_C95_net11586, mult_28_C95_net11587, 
      mult_28_C95_n132, mult_28_C95_n161, mult_28_C95_n51, mult_28_C95_n377, 
      mult_28_C95_n378, mult_28_C95_n380, mult_28_C95_n384, mult_28_C95_n180, 
      mult_28_C95_n187, mult_28_C95_n203, mult_28_C95_n204, mult_28_C95_n205, 
      mult_28_C95_net12065, mult_28_C95_n804, mult_28_C95_net12285, 
      mult_28_C95_net12257, mult_28_C95_net12249, mult_28_C95_net12250, 
      mult_28_C95_net12183, mult_28_C95_net12151, mult_28_C95_net12152, 
      mult_28_C95_net12153, mult_28_C95_net12125, mult_28_C95_net12126, 
      mult_28_C95_net12127, mult_28_C95_net12095, mult_28_C95_net12078, 
      mult_28_C95_net12079, mult_28_C95_net12054, mult_28_C95_net12055, 
      mult_28_C95_net12033, mult_28_C95_net11829, mult_28_C95_net11745, 
      mult_28_C95_net11746, mult_28_C95_net11693, mult_28_C95_net11666, 
      mult_28_C95_net11667, mult_28_C95_net11662, mult_28_C95_net11503, 
      mult_28_C95_net11507, mult_28_C95_net11509, mult_28_C95_net11172, 
      mult_28_C95_net11083, mult_28_C95_net11025, mult_28_C95_n832, 
      mult_28_C95_n831, mult_28_C95_n830, mult_28_C95_n829, mult_28_C95_n828, 
      mult_28_C95_n827, mult_28_C95_n826, mult_28_C95_n824, mult_28_C95_n808, 
      mult_28_C95_n807, mult_28_C95_n806, mult_28_C95_n805, mult_28_C95_n801, 
      mult_28_C95_n784, mult_28_C95_n783, mult_28_C95_n782, mult_28_C95_n781, 
      mult_28_C95_n780, mult_28_C95_n779, mult_28_C95_n778, mult_28_C95_n777, 
      mult_28_C95_n776, mult_28_C95_n775, mult_28_C95_n774, mult_28_C95_n773, 
      mult_28_C95_n772, mult_28_C95_n771, mult_28_C95_n770, mult_28_C95_n769, 
      mult_28_C95_n768, mult_28_C95_n767, mult_28_C95_n766, mult_28_C95_n765, 
      mult_28_C95_n764, mult_28_C95_n763, mult_28_C95_n762, mult_28_C95_n761, 
      mult_28_C95_n760, mult_28_C95_n759, mult_28_C95_n758, mult_28_C95_n757, 
      mult_28_C95_n756, mult_28_C95_n755, mult_28_C95_n754, mult_28_C95_n753, 
      mult_28_C95_n752, mult_28_C95_n751, mult_28_C95_n750, mult_28_C95_n749, 
      mult_28_C95_n748, mult_28_C95_n747, mult_28_C95_n746, mult_28_C95_n745, 
      mult_28_C95_n744, mult_28_C95_n743, mult_28_C95_n742, mult_28_C95_n741, 
      mult_28_C95_n740, mult_28_C95_n739, mult_28_C95_n738, mult_28_C95_n737, 
      mult_28_C95_n736, mult_28_C95_n735, mult_28_C95_n734, mult_28_C95_n733, 
      mult_28_C95_n732, mult_28_C95_n731, mult_28_C95_n730, mult_28_C95_n729, 
      mult_28_C95_n728, mult_28_C95_n727, mult_28_C95_n726, mult_28_C95_n725, 
      mult_28_C95_n724, mult_28_C95_n723, mult_28_C95_n722, mult_28_C95_n721, 
      mult_28_C95_n720, mult_28_C95_n719, mult_28_C95_n718, mult_28_C95_n717, 
      mult_28_C95_n716, mult_28_C95_n715, mult_28_C95_n714, mult_28_C95_n713, 
      mult_28_C95_n712, mult_28_C95_n711, mult_28_C95_n710, mult_28_C95_n709, 
      mult_28_C95_n708, mult_28_C95_n705, mult_28_C95_n704, mult_28_C95_n703, 
      mult_28_C95_n702, mult_28_C95_n701, mult_28_C95_n700, mult_28_C95_n699, 
      mult_28_C95_n698, mult_28_C95_n697, mult_28_C95_n696, mult_28_C95_n695, 
      mult_28_C95_n694, mult_28_C95_n691, mult_28_C95_n690, mult_28_C95_n689, 
      mult_28_C95_n688, mult_28_C95_n687, mult_28_C95_n686, mult_28_C95_n685, 
      mult_28_C95_n684, mult_28_C95_n683, mult_28_C95_n682, mult_28_C95_n681, 
      mult_28_C95_n680, mult_28_C95_n679, mult_28_C95_n676, mult_28_C95_n675, 
      mult_28_C95_n674, mult_28_C95_n673, mult_28_C95_n672, mult_28_C95_n671, 
      mult_28_C95_n670, mult_28_C95_n669, mult_28_C95_n668, mult_28_C95_n667, 
      mult_28_C95_n666, mult_28_C95_n665, mult_28_C95_n664, mult_28_C95_n663, 
      mult_28_C95_n662, mult_28_C95_n661, mult_28_C95_n660, mult_28_C95_n659, 
      mult_28_C95_n658, mult_28_C95_n657, mult_28_C95_n656, mult_28_C95_n655, 
      mult_28_C95_n654, mult_28_C95_n653, mult_28_C95_n652, mult_28_C95_n651, 
      mult_28_C95_n650, mult_28_C95_n649, mult_28_C95_n648, mult_28_C95_n647, 
      mult_28_C95_n646, mult_28_C95_n645, mult_28_C95_n644, mult_28_C95_n643, 
      mult_28_C95_n642, mult_28_C95_n641, mult_28_C95_n640, mult_28_C95_n639, 
      mult_28_C95_n638, mult_28_C95_n637, mult_28_C95_n636, mult_28_C95_n635, 
      mult_28_C95_n632, mult_28_C95_n631, mult_28_C95_n630, mult_28_C95_n629, 
      mult_28_C95_n628, mult_28_C95_n627, mult_28_C95_n626, mult_28_C95_n625, 
      mult_28_C95_n624, mult_28_C95_n623, mult_28_C95_n622, mult_28_C95_n621, 
      mult_28_C95_n620, mult_28_C95_n619, mult_28_C95_n618, mult_28_C95_n616, 
      mult_28_C95_n615, mult_28_C95_n614, mult_28_C95_n613, mult_28_C95_n612, 
      mult_28_C95_n611, mult_28_C95_n610, mult_28_C95_n609, mult_28_C95_n608, 
      mult_28_C95_n607, mult_28_C95_n606, mult_28_C95_n605, mult_28_C95_n604, 
      mult_28_C95_n603, mult_28_C95_n602, mult_28_C95_n601, mult_28_C95_n600, 
      mult_28_C95_n599, mult_28_C95_n598, mult_28_C95_n597, mult_28_C95_n596, 
      mult_28_C95_n595, mult_28_C95_n594, mult_28_C95_n593, mult_28_C95_n592, 
      mult_28_C95_n591, mult_28_C95_n590, mult_28_C95_n588, mult_28_C95_n587, 
      mult_28_C95_n586, mult_28_C95_n585, mult_28_C95_n584, mult_28_C95_n583, 
      mult_28_C95_n582, mult_28_C95_n581, mult_28_C95_n580, mult_28_C95_n579, 
      mult_28_C95_n578, mult_28_C95_n577, mult_28_C95_n576, mult_28_C95_n575, 
      mult_28_C95_n574, mult_28_C95_n573, mult_28_C95_n571, mult_28_C95_n570, 
      mult_28_C95_n569, mult_28_C95_n568, mult_28_C95_n567, mult_28_C95_n566, 
      mult_28_C95_n565, mult_28_C95_n564, mult_28_C95_n563, mult_28_C95_n562, 
      mult_28_C95_n561, mult_28_C95_n560, mult_28_C95_n559, mult_28_C95_n556, 
      mult_28_C95_n555, mult_28_C95_n554, mult_28_C95_n553, mult_28_C95_n552, 
      mult_28_C95_n551, mult_28_C95_n550, mult_28_C95_n549, mult_28_C95_n548, 
      mult_28_C95_n547, mult_28_C95_n546, mult_28_C95_n544, mult_28_C95_n542, 
      mult_28_C95_n541, mult_28_C95_n540, mult_28_C95_n539, mult_28_C95_n538, 
      mult_28_C95_n537, mult_28_C95_n536, mult_28_C95_n535, mult_28_C95_n534, 
      mult_28_C95_n533, mult_28_C95_n532, mult_28_C95_n531, mult_28_C95_n530, 
      mult_28_C95_n529, mult_28_C95_n528, mult_28_C95_n527, mult_28_C95_n526, 
      mult_28_C95_n525, mult_28_C95_n524, mult_28_C95_n523, mult_28_C95_n522, 
      mult_28_C95_n520, mult_28_C95_n519, mult_28_C95_n518, mult_28_C95_n517, 
      mult_28_C95_n516, mult_28_C95_n515, mult_28_C95_n514, mult_28_C95_n513, 
      mult_28_C95_n512, mult_28_C95_n511, mult_28_C95_n510, mult_28_C95_n509, 
      mult_28_C95_n508, mult_28_C95_n507, mult_28_C95_n506, mult_28_C95_n505, 
      mult_28_C95_n504, mult_28_C95_n503, mult_28_C95_n502, mult_28_C95_n501, 
      mult_28_C95_n500, mult_28_C95_n499, mult_28_C95_n498, mult_28_C95_n497, 
      mult_28_C95_n496, mult_28_C95_n495, mult_28_C95_n494, mult_28_C95_n493, 
      mult_28_C95_n492, mult_28_C95_n491, mult_28_C95_n490, mult_28_C95_n489, 
      mult_28_C95_n488, mult_28_C95_n487, mult_28_C95_n486, mult_28_C95_n485, 
      mult_28_C95_n484, mult_28_C95_n483, mult_28_C95_n482, mult_28_C95_n481, 
      mult_28_C95_n480, mult_28_C95_n479, mult_28_C95_n478, mult_28_C95_n477, 
      mult_28_C95_n476, mult_28_C95_n475, mult_28_C95_n474, mult_28_C95_n473, 
      mult_28_C95_n472, mult_28_C95_n471, mult_28_C95_n470, mult_28_C95_n469, 
      mult_28_C95_n468, mult_28_C95_n467, mult_28_C95_n466, mult_28_C95_n465, 
      mult_28_C95_n464, mult_28_C95_n463, mult_28_C95_n462, mult_28_C95_n461, 
      mult_28_C95_n460, mult_28_C95_n459, mult_28_C95_n458, mult_28_C95_n457, 
      mult_28_C95_n456, mult_28_C95_n455, mult_28_C95_n454, mult_28_C95_n453, 
      mult_28_C95_n452, mult_28_C95_n451, mult_28_C95_n450, mult_28_C95_n449, 
      mult_28_C95_n448, mult_28_C95_n447, mult_28_C95_n446, mult_28_C95_n445, 
      mult_28_C95_n444, mult_28_C95_n443, mult_28_C95_n442, mult_28_C95_n441, 
      mult_28_C95_n438, mult_28_C95_n437, mult_28_C95_n436, mult_28_C95_n435, 
      mult_28_C95_n434, mult_28_C95_n433, mult_28_C95_n432, mult_28_C95_n431, 
      mult_28_C95_n430, mult_28_C95_n429, mult_28_C95_n428, mult_28_C95_n427, 
      mult_28_C95_n426, mult_28_C95_n425, mult_28_C95_n422, mult_28_C95_n420, 
      mult_28_C95_n419, mult_28_C95_n418, mult_28_C95_n417, mult_28_C95_n416, 
      mult_28_C95_n415, mult_28_C95_n413, mult_28_C95_n410, mult_28_C95_n408, 
      mult_28_C95_n407, mult_28_C95_n404, mult_28_C95_n403, mult_28_C95_n402, 
      mult_28_C95_n401, mult_28_C95_n400, mult_28_C95_n399, mult_28_C95_n398, 
      mult_28_C95_n397, mult_28_C95_n394, mult_28_C95_n393, mult_28_C95_n388, 
      mult_28_C95_n386, mult_28_C95_n385, mult_28_C95_n383, mult_28_C95_n382, 
      mult_28_C95_n381, mult_28_C95_n379, mult_28_C95_n374, mult_28_C95_n373, 
      mult_28_C95_n372, mult_28_C95_n371, mult_28_C95_n370, mult_28_C95_n369, 
      mult_28_C95_n368, mult_28_C95_n367, mult_28_C95_n366, mult_28_C95_n365, 
      mult_28_C95_n364, mult_28_C95_n363, mult_28_C95_n362, mult_28_C95_n361, 
      mult_28_C95_n360, mult_28_C95_n359, mult_28_C95_n358, mult_28_C95_n357, 
      mult_28_C95_n356, mult_28_C95_n355, mult_28_C95_n354, mult_28_C95_n353, 
      mult_28_C95_n352, mult_28_C95_n351, mult_28_C95_n350, mult_28_C95_n349, 
      mult_28_C95_n348, mult_28_C95_n347, mult_28_C95_n346, mult_28_C95_n345, 
      mult_28_C95_n344, mult_28_C95_n343, mult_28_C95_n342, mult_28_C95_n341, 
      mult_28_C95_n340, mult_28_C95_n339, mult_28_C95_n338, mult_28_C95_n337, 
      mult_28_C95_n336, mult_28_C95_n335, mult_28_C95_n334, mult_28_C95_n333, 
      mult_28_C95_n332, mult_28_C95_n331, mult_28_C95_n330, mult_28_C95_n329, 
      mult_28_C95_n328, mult_28_C95_n327, mult_28_C95_n326, mult_28_C95_n325, 
      mult_28_C95_n324, mult_28_C95_n323, mult_28_C95_n322, mult_28_C95_n321, 
      mult_28_C95_n320, mult_28_C95_n319, mult_28_C95_n318, mult_28_C95_n317, 
      mult_28_C95_n316, mult_28_C95_n315, mult_28_C95_n314, mult_28_C95_n313, 
      mult_28_C95_n312, mult_28_C95_n311, mult_28_C95_n310, mult_28_C95_n309, 
      mult_28_C95_n308, mult_28_C95_n307, mult_28_C95_n306, mult_28_C95_n305, 
      mult_28_C95_n288, mult_28_C95_n287, mult_28_C95_n285, mult_28_C95_n284, 
      mult_28_C95_n283, mult_28_C95_n279, mult_28_C95_n278, mult_28_C95_n267, 
      mult_28_C95_n266, mult_28_C95_n265, mult_28_C95_n264, mult_28_C95_n259, 
      mult_28_C95_n258, mult_28_C95_n257, mult_28_C95_n256, mult_28_C95_n251, 
      mult_28_C95_n250, mult_28_C95_n249, mult_28_C95_n248, mult_28_C95_n243, 
      mult_28_C95_n232, mult_28_C95_n231, mult_28_C95_n230, mult_28_C95_n225, 
      mult_28_C95_n214, mult_28_C95_n213, mult_28_C95_n212, mult_28_C95_n211, 
      mult_28_C95_n210, mult_28_C95_n209, mult_28_C95_n208, mult_28_C95_n207, 
      mult_28_C95_n206, mult_28_C95_n202, mult_28_C95_n201, mult_28_C95_n200, 
      mult_28_C95_n199, mult_28_C95_n197, mult_28_C95_n196, mult_28_C95_n195, 
      mult_28_C95_n192, mult_28_C95_n188, mult_28_C95_n183, mult_28_C95_n182, 
      mult_28_C95_n173, mult_28_C95_n172, mult_28_C95_n171, mult_28_C95_n169, 
      mult_28_C95_n168, mult_28_C95_n167, mult_28_C95_n160, mult_28_C95_n148, 
      mult_28_C95_n142, mult_28_C95_n141, mult_28_C95_n140, mult_28_C95_n139, 
      mult_28_C95_n135, mult_28_C95_n129, mult_28_C95_n128, mult_28_C95_n127, 
      mult_28_C95_n124, mult_28_C95_n118, mult_28_C95_n117, mult_28_C95_n116, 
      mult_28_C95_n115, mult_28_C95_n114, mult_28_C95_n113, mult_28_C95_n112, 
      mult_28_C95_n109, mult_28_C95_n108, mult_28_C95_n107, mult_28_C95_n106, 
      mult_28_C95_n105, mult_28_C95_n104, mult_28_C95_n103, mult_28_C95_n102, 
      mult_28_C95_n101, mult_28_C95_n100, mult_28_C95_n97, mult_28_C95_n96, 
      mult_28_C95_n95, mult_28_C95_n94, mult_28_C95_n93, mult_28_C95_n92, 
      mult_28_C95_n87, mult_28_C95_n86, mult_28_C95_n85, mult_28_C95_n84, 
      mult_28_C95_n69, mult_28_C95_n68, mult_28_C95_n67, mult_28_C95_n65, 
      mult_28_C95_n63, mult_28_C95_n56, mult_28_C95_n55, mult_28_C95_n54, 
      mult_28_C95_n53, mult_28_C95_n52, mult_28_C95_n48, mult_28_C95_n46, 
      mult_28_C95_n42, mult_28_C95_n40, mult_28_C95_n36, mult_28_C95_n34, 
      mult_28_C95_n30, mult_28_C95_n28, mult_28_C95_n24, mult_28_C95_n22, 
      mult_28_C95_n18, mult_28_C95_n16, mult_28_C95_n12, mult_28_C95_n9, 
      mult_28_C95_n6, mult_28_C96_n_1016, mult_28_C96_n1094, mult_28_C96_n1093,
      mult_28_C96_n1092, mult_28_C96_n1091, mult_28_C96_n1090, 
      mult_28_C96_n1089, mult_28_C96_n1088, mult_28_C96_n1087, 
      mult_28_C96_n1086, mult_28_C96_n1085, mult_28_C96_n1084, 
      mult_28_C96_n1083, mult_28_C96_n1082, mult_28_C96_n1081, 
      mult_28_C96_n1080, mult_28_C96_n1079, mult_28_C96_n1078, 
      mult_28_C96_n1077, mult_28_C96_n1076, mult_28_C96_n1075, 
      mult_28_C96_n1074, mult_28_C96_n1073, mult_28_C96_n1072, 
      mult_28_C96_n1071, mult_28_C96_n1070, mult_28_C96_n1069, 
      mult_28_C96_n1068, mult_28_C96_n1067, mult_28_C96_n1066, 
      mult_28_C96_n1065, mult_28_C96_n1064, mult_28_C96_n1063, 
      mult_28_C96_n1062, mult_28_C96_n1061, mult_28_C96_n1060, 
      mult_28_C96_n1059, mult_28_C96_n1058, mult_28_C96_n1057, 
      mult_28_C96_n1056, mult_28_C96_n1055, mult_28_C96_n1054, 
      mult_28_C96_n1053, mult_28_C96_n1052, mult_28_C96_n1051, 
      mult_28_C96_n1050, mult_28_C96_n1049, mult_28_C96_n1048, 
      mult_28_C96_n1047, mult_28_C96_n1046, mult_28_C96_n1045, 
      mult_28_C96_n1044, mult_28_C96_n1043, mult_28_C96_n1042, 
      mult_28_C96_n1041, mult_28_C96_n1040, mult_28_C96_n1039, 
      mult_28_C96_n1038, mult_28_C96_n1037, mult_28_C96_n1036, 
      mult_28_C96_n1035, mult_28_C96_n1034, mult_28_C96_n1033, 
      mult_28_C96_n1032, mult_28_C96_n1031, mult_28_C96_n1030, 
      mult_28_C96_n1029, mult_28_C96_n1028, mult_28_C96_n1027, 
      mult_28_C96_n1026, mult_28_C96_n1025, mult_28_C96_n1024, 
      mult_28_C96_n1023, mult_28_C96_n1022, mult_28_C96_n1021, 
      mult_28_C96_n1020, mult_28_C96_n1019, mult_28_C96_n1018, 
      mult_28_C96_n1017, mult_28_C96_n1016, mult_28_C96_n1015, 
      mult_28_C96_n1014, mult_28_C96_n1013, mult_28_C96_n1012, 
      mult_28_C96_n1011, mult_28_C96_n1010, mult_28_C96_n1009, 
      mult_28_C96_n1008, mult_28_C96_n1007, mult_28_C96_n1006, 
      mult_28_C96_n1005, mult_28_C96_n1004, mult_28_C96_n1003, 
      mult_28_C96_n1002, mult_28_C96_n1001, mult_28_C96_n1000, mult_28_C96_n999
      , mult_28_C96_n998, mult_28_C96_n997, mult_28_C96_n996, mult_28_C96_n995,
      mult_28_C96_n994, mult_28_C96_n993, mult_28_C96_n992, mult_28_C96_n991, 
      mult_28_C96_n990, mult_28_C96_n989, mult_28_C96_n988, mult_28_C96_n987, 
      mult_28_C96_n986, mult_28_C96_n985, mult_28_C96_n984, mult_28_C96_n983, 
      mult_28_C96_n982, mult_28_C96_n981, mult_28_C96_n980, mult_28_C96_n979, 
      mult_28_C96_n978, mult_28_C96_n977, mult_28_C96_n976, mult_28_C96_n975, 
      mult_28_C96_n974, mult_28_C96_n973, mult_28_C96_n972, mult_28_C96_n971, 
      mult_28_C96_n970, mult_28_C96_n969, mult_28_C96_n968, mult_28_C96_n967, 
      mult_28_C96_n966, mult_28_C96_n965, mult_28_C96_n964, mult_28_C96_n963, 
      mult_28_C96_n962, mult_28_C96_n961, mult_28_C96_n960, mult_28_C96_n959, 
      mult_28_C96_n958, mult_28_C96_n957, mult_28_C96_n956, mult_28_C96_n955, 
      mult_28_C96_n954, mult_28_C96_n953, mult_28_C96_n952, mult_28_C96_n951, 
      mult_28_C96_n950, mult_28_C96_n949, mult_28_C96_n948, mult_28_C96_n947, 
      mult_28_C96_n946, mult_28_C96_n945, mult_28_C96_n944, mult_28_C96_n943, 
      mult_28_C96_n942, mult_28_C96_n941, mult_28_C96_n940, mult_28_C96_n939, 
      mult_28_C96_n938, mult_28_C96_n937, mult_28_C96_n936, mult_28_C96_n935, 
      mult_28_C96_n934, mult_28_C96_n933, mult_28_C96_n932, mult_28_C96_n931, 
      mult_28_C96_n930, mult_28_C96_n929, mult_28_C96_n928, mult_28_C96_n927, 
      mult_28_C96_n926, mult_28_C96_n925, mult_28_C96_n924, mult_28_C96_n923, 
      mult_28_C96_n922, mult_28_C96_n921, mult_28_C96_n920, mult_28_C96_n919, 
      mult_28_C96_n918, mult_28_C96_n917, mult_28_C96_n916, mult_28_C96_n915, 
      mult_28_C96_n914, mult_28_C96_n913, mult_28_C96_n912, mult_28_C96_n911, 
      mult_28_C96_n910, mult_28_C96_n909, mult_28_C96_n908, mult_28_C96_n907, 
      mult_28_C96_n906, mult_28_C96_n905, mult_28_C96_n904, mult_28_C96_n903, 
      mult_28_C96_n902, mult_28_C96_n901, mult_28_C96_n900, mult_28_C96_n832, 
      mult_28_C96_n831, mult_28_C96_n830, mult_28_C96_n829, mult_28_C96_n828, 
      mult_28_C96_n827, mult_28_C96_n826, mult_28_C96_n825, mult_28_C96_n824, 
      mult_28_C96_n808, mult_28_C96_n807, mult_28_C96_n806, mult_28_C96_n805, 
      mult_28_C96_n804, mult_28_C96_n803, mult_28_C96_n802, mult_28_C96_n801, 
      mult_28_C96_n784, mult_28_C96_n783, mult_28_C96_n782, mult_28_C96_n781, 
      mult_28_C96_n780, mult_28_C96_n779, mult_28_C96_n778, mult_28_C96_n777, 
      mult_28_C96_n776, mult_28_C96_n775, mult_28_C96_n774, mult_28_C96_n773, 
      mult_28_C96_n772, mult_28_C96_n771, mult_28_C96_n770, mult_28_C96_n769, 
      mult_28_C96_n768, mult_28_C96_n767, mult_28_C96_n766, mult_28_C96_n765, 
      mult_28_C96_n764, mult_28_C96_n763, mult_28_C96_n762, mult_28_C96_n761, 
      mult_28_C96_n760, mult_28_C96_n759, mult_28_C96_n758, mult_28_C96_n757, 
      mult_28_C96_n756, mult_28_C96_n755, mult_28_C96_n754, mult_28_C96_n753, 
      mult_28_C96_n752, mult_28_C96_n751, mult_28_C96_n750, mult_28_C96_n749, 
      mult_28_C96_n748, mult_28_C96_n747, mult_28_C96_n746, mult_28_C96_n745, 
      mult_28_C96_n744, mult_28_C96_n743, mult_28_C96_n742, mult_28_C96_n741, 
      mult_28_C96_n740, mult_28_C96_n738, mult_28_C96_n737, mult_28_C96_n736, 
      mult_28_C96_n735, mult_28_C96_n734, mult_28_C96_n733, mult_28_C96_n732, 
      mult_28_C96_n731, mult_28_C96_n730, mult_28_C96_n729, mult_28_C96_n728, 
      mult_28_C96_n727, mult_28_C96_n726, mult_28_C96_n725, mult_28_C96_n724, 
      mult_28_C96_n723, mult_28_C96_n722, mult_28_C96_n721, mult_28_C96_n720, 
      mult_28_C96_n719, mult_28_C96_n718, mult_28_C96_n717, mult_28_C96_n716, 
      mult_28_C96_n715, mult_28_C96_n714, mult_28_C96_n713, mult_28_C96_n712, 
      mult_28_C96_n711, mult_28_C96_n710, mult_28_C96_n709, mult_28_C96_n708, 
      mult_28_C96_n707, mult_28_C96_n706, mult_28_C96_n705, mult_28_C96_n704, 
      mult_28_C96_n703, mult_28_C96_n702, mult_28_C96_n701, mult_28_C96_n700, 
      mult_28_C96_n699, mult_28_C96_n698, mult_28_C96_n697, mult_28_C96_n696, 
      mult_28_C96_n695, mult_28_C96_n694, mult_28_C96_n693, mult_28_C96_n692, 
      mult_28_C96_n691, mult_28_C96_n690, mult_28_C96_n689, mult_28_C96_n688, 
      mult_28_C96_n687, mult_28_C96_n686, mult_28_C96_n685, mult_28_C96_n684, 
      mult_28_C96_n683, mult_28_C96_n682, mult_28_C96_n681, mult_28_C96_n680, 
      mult_28_C96_n679, mult_28_C96_n678, mult_28_C96_n677, mult_28_C96_n676, 
      mult_28_C96_n675, mult_28_C96_n674, mult_28_C96_n673, mult_28_C96_n672, 
      mult_28_C96_n671, mult_28_C96_n670, mult_28_C96_n669, mult_28_C96_n668, 
      mult_28_C96_n667, mult_28_C96_n666, mult_28_C96_n665, mult_28_C96_n664, 
      mult_28_C96_n663, mult_28_C96_n662, mult_28_C96_n661, mult_28_C96_n660, 
      mult_28_C96_n659, mult_28_C96_n658, mult_28_C96_n657, mult_28_C96_n656, 
      mult_28_C96_n655, mult_28_C96_n654, mult_28_C96_n653, mult_28_C96_n652, 
      mult_28_C96_n651, mult_28_C96_n650, mult_28_C96_n649, mult_28_C96_n648, 
      mult_28_C96_n647, mult_28_C96_n646, mult_28_C96_n645, mult_28_C96_n644, 
      mult_28_C96_n643, mult_28_C96_n642, mult_28_C96_n641, mult_28_C96_n640, 
      mult_28_C96_n639, mult_28_C96_n638, mult_28_C96_n637, mult_28_C96_n636, 
      mult_28_C96_n635, mult_28_C96_n634, mult_28_C96_n633, mult_28_C96_n632, 
      mult_28_C96_n631, mult_28_C96_n630, mult_28_C96_n629, mult_28_C96_n628, 
      mult_28_C96_n627, mult_28_C96_n626, mult_28_C96_n625, mult_28_C96_n624, 
      mult_28_C96_n623, mult_28_C96_n622, mult_28_C96_n621, mult_28_C96_n620, 
      mult_28_C96_n619, mult_28_C96_n618, mult_28_C96_n617, mult_28_C96_n616, 
      mult_28_C96_n615, mult_28_C96_n614, mult_28_C96_n613, mult_28_C96_n612, 
      mult_28_C96_n611, mult_28_C96_n610, mult_28_C96_n609, mult_28_C96_n608, 
      mult_28_C96_n607, mult_28_C96_n606, mult_28_C96_n605, mult_28_C96_n604, 
      mult_28_C96_n603, mult_28_C96_n602, mult_28_C96_n601, mult_28_C96_n600, 
      mult_28_C96_n599, mult_28_C96_n598, mult_28_C96_n597, mult_28_C96_n596, 
      mult_28_C96_n595, mult_28_C96_n594, mult_28_C96_n593, mult_28_C96_n592, 
      mult_28_C96_n591, mult_28_C96_n590, mult_28_C96_n589, mult_28_C96_n588, 
      mult_28_C96_n587, mult_28_C96_n586, mult_28_C96_n585, mult_28_C96_n584, 
      mult_28_C96_n583, mult_28_C96_n582, mult_28_C96_n581, mult_28_C96_n580, 
      mult_28_C96_n579, mult_28_C96_n578, mult_28_C96_n577, mult_28_C96_n576, 
      mult_28_C96_n575, mult_28_C96_n574, mult_28_C96_n573, mult_28_C96_n572, 
      mult_28_C96_n571, mult_28_C96_n570, mult_28_C96_n569, mult_28_C96_n568, 
      mult_28_C96_n567, mult_28_C96_n566, mult_28_C96_n565, mult_28_C96_n564, 
      mult_28_C96_n563, mult_28_C96_n562, mult_28_C96_n561, mult_28_C96_n560, 
      mult_28_C96_n559, mult_28_C96_n558, mult_28_C96_n557, mult_28_C96_n556, 
      mult_28_C96_n555, mult_28_C96_n554, mult_28_C96_n553, mult_28_C96_n552, 
      mult_28_C96_n551, mult_28_C96_n550, mult_28_C96_n549, mult_28_C96_n548, 
      mult_28_C96_n547, mult_28_C96_n546, mult_28_C96_n545, mult_28_C96_n544, 
      mult_28_C96_n543, mult_28_C96_n542, mult_28_C96_n541, mult_28_C96_n540, 
      mult_28_C96_n539, mult_28_C96_n538, mult_28_C96_n537, mult_28_C96_n536, 
      mult_28_C96_n535, mult_28_C96_n534, mult_28_C96_n533, mult_28_C96_n532, 
      mult_28_C96_n531, mult_28_C96_n530, mult_28_C96_n529, mult_28_C96_n528, 
      mult_28_C96_n527, mult_28_C96_n526, mult_28_C96_n525, mult_28_C96_n524, 
      mult_28_C96_n523, mult_28_C96_n522, mult_28_C96_n520, mult_28_C96_n519, 
      mult_28_C96_n518, mult_28_C96_n517, mult_28_C96_n516, mult_28_C96_n515, 
      mult_28_C96_n514, mult_28_C96_n513, mult_28_C96_n512, mult_28_C96_n511, 
      mult_28_C96_n510, mult_28_C96_n509, mult_28_C96_n508, mult_28_C96_n507, 
      mult_28_C96_n506, mult_28_C96_n505, mult_28_C96_n504, mult_28_C96_n503, 
      mult_28_C96_n502, mult_28_C96_n501, mult_28_C96_n500, mult_28_C96_n499, 
      mult_28_C96_n498, mult_28_C96_n497, mult_28_C96_n496, mult_28_C96_n495, 
      mult_28_C96_n494, mult_28_C96_n493, mult_28_C96_n492, mult_28_C96_n491, 
      mult_28_C96_n490, mult_28_C96_n489, mult_28_C96_n488, mult_28_C96_n487, 
      mult_28_C96_n486, mult_28_C96_n485, mult_28_C96_n484, mult_28_C96_n483, 
      mult_28_C96_n482, mult_28_C96_n481, mult_28_C96_n480, mult_28_C96_n479, 
      mult_28_C96_n478, mult_28_C96_n477, mult_28_C96_n476, mult_28_C96_n475, 
      mult_28_C96_n474, mult_28_C96_n473, mult_28_C96_n472, mult_28_C96_n471, 
      mult_28_C96_n470, mult_28_C96_n469, mult_28_C96_n468, mult_28_C96_n467, 
      mult_28_C96_n466, mult_28_C96_n465, mult_28_C96_n464, mult_28_C96_n463, 
      mult_28_C96_n462, mult_28_C96_n461, mult_28_C96_n460, mult_28_C96_n459, 
      mult_28_C96_n458, mult_28_C96_n457, mult_28_C96_n456, mult_28_C96_n455, 
      mult_28_C96_n454, mult_28_C96_n453, mult_28_C96_n452, mult_28_C96_n451, 
      mult_28_C96_n450, mult_28_C96_n449, mult_28_C96_n448, mult_28_C96_n447, 
      mult_28_C96_n446, mult_28_C96_n445, mult_28_C96_n444, mult_28_C96_n443, 
      mult_28_C96_n442, mult_28_C96_n441, mult_28_C96_n440, mult_28_C96_n439, 
      mult_28_C96_n438, mult_28_C96_n437, mult_28_C96_n436, mult_28_C96_n435, 
      mult_28_C96_n434, mult_28_C96_n433, mult_28_C96_n432, mult_28_C96_n431, 
      mult_28_C96_n430, mult_28_C96_n429, mult_28_C96_n428, mult_28_C96_n427, 
      mult_28_C96_n426, mult_28_C96_n425, mult_28_C96_n424, mult_28_C96_n423, 
      mult_28_C96_n422, mult_28_C96_n421, mult_28_C96_n420, mult_28_C96_n419, 
      mult_28_C96_n418, mult_28_C96_n417, mult_28_C96_n416, mult_28_C96_n415, 
      mult_28_C96_n414, mult_28_C96_n413, mult_28_C96_n412, mult_28_C96_n411, 
      mult_28_C96_n410, mult_28_C96_n409, mult_28_C96_n408, mult_28_C96_n407, 
      mult_28_C96_n406, mult_28_C96_n405, mult_28_C96_n404, mult_28_C96_n403, 
      mult_28_C96_n402, mult_28_C96_n401, mult_28_C96_n400, mult_28_C96_n399, 
      mult_28_C96_n398, mult_28_C96_n397, mult_28_C96_n396, mult_28_C96_n395, 
      mult_28_C96_n394, mult_28_C96_n393, mult_28_C96_n392, mult_28_C96_n391, 
      mult_28_C96_n390, mult_28_C96_n389, mult_28_C96_n388, mult_28_C96_n387, 
      mult_28_C96_n386, mult_28_C96_n385, mult_28_C96_n384, mult_28_C96_n383, 
      mult_28_C96_n382, mult_28_C96_n381, mult_28_C96_n380, mult_28_C96_n379, 
      mult_28_C96_n378, mult_28_C96_n377, mult_28_C96_n376, mult_28_C96_n375, 
      mult_28_C96_n374, mult_28_C96_n373, mult_28_C96_n372, mult_28_C96_n371, 
      mult_28_C96_n370, mult_28_C96_n369, mult_28_C96_n368, mult_28_C96_n367, 
      mult_28_C96_n366, mult_28_C96_n365, mult_28_C96_n364, mult_28_C96_n363, 
      mult_28_C96_n362, mult_28_C96_n361, mult_28_C96_n360, mult_28_C96_n359, 
      mult_28_C96_n358, mult_28_C96_n357, mult_28_C96_n356, mult_28_C96_n355, 
      mult_28_C96_n354, mult_28_C96_n353, mult_28_C96_n352, mult_28_C96_n351, 
      mult_28_C96_n350, mult_28_C96_n349, mult_28_C96_n348, mult_28_C96_n347, 
      mult_28_C96_n346, mult_28_C96_n345, mult_28_C96_n344, mult_28_C96_n343, 
      mult_28_C96_n342, mult_28_C96_n341, mult_28_C96_n340, mult_28_C96_n339, 
      mult_28_C96_n338, mult_28_C96_n337, mult_28_C96_n336, mult_28_C96_n335, 
      mult_28_C96_n334, mult_28_C96_n333, mult_28_C96_n332, mult_28_C96_n331, 
      mult_28_C96_n330, mult_28_C96_n329, mult_28_C96_n328, mult_28_C96_n327, 
      mult_28_C96_n326, mult_28_C96_n325, mult_28_C96_n324, mult_28_C96_n323, 
      mult_28_C96_n322, mult_28_C96_n321, mult_28_C96_n320, mult_28_C96_n319, 
      mult_28_C96_n318, mult_28_C96_n317, mult_28_C96_n316, mult_28_C96_n315, 
      mult_28_C96_n314, mult_28_C96_n313, mult_28_C96_n312, mult_28_C96_n311, 
      mult_28_C96_n310, mult_28_C96_n309, mult_28_C96_n308, mult_28_C96_n307, 
      mult_28_C96_n306, mult_28_C96_n305, mult_28_C96_n288, mult_28_C96_n286, 
      mult_28_C96_n285, mult_28_C96_n284, mult_28_C96_n283, mult_28_C96_n282, 
      mult_28_C96_n281, mult_28_C96_n279, mult_28_C96_n278, mult_28_C96_n276, 
      mult_28_C96_n267, mult_28_C96_n266, mult_28_C96_n265, mult_28_C96_n264, 
      mult_28_C96_n259, mult_28_C96_n258, mult_28_C96_n257, mult_28_C96_n256, 
      mult_28_C96_n251, mult_28_C96_n250, mult_28_C96_n249, mult_28_C96_n248, 
      mult_28_C96_n243, mult_28_C96_n232, mult_28_C96_n230, mult_28_C96_n225, 
      mult_28_C96_n223, mult_28_C96_n217, mult_28_C96_n215, mult_28_C96_n214, 
      mult_28_C96_n213, mult_28_C96_n212, mult_28_C96_n211, mult_28_C96_n210, 
      mult_28_C96_n209, mult_28_C96_n208, mult_28_C96_n207, mult_28_C96_n206, 
      mult_28_C96_n205, mult_28_C96_n204, mult_28_C96_n203, mult_28_C96_n202, 
      mult_28_C96_n201, mult_28_C96_n200, mult_28_C96_n199, mult_28_C96_n197, 
      mult_28_C96_n196, mult_28_C96_n195, mult_28_C96_n192, mult_28_C96_n190, 
      mult_28_C96_n189, mult_28_C96_n188, mult_28_C96_n187, mult_28_C96_n184, 
      mult_28_C96_n183, mult_28_C96_n182, mult_28_C96_n180, mult_28_C96_n179, 
      mult_28_C96_n178, mult_28_C96_n177, mult_28_C96_n176, mult_28_C96_n175, 
      mult_28_C96_n173, mult_28_C96_n169, mult_28_C96_n168, mult_28_C96_n167, 
      mult_28_C96_n164, mult_28_C96_n163, mult_28_C96_n162, mult_28_C96_n161, 
      mult_28_C96_n160, mult_28_C96_n155, mult_28_C96_n154, mult_28_C96_n153, 
      mult_28_C96_n152, mult_28_C96_n151, mult_28_C96_n150, mult_28_C96_n149, 
      mult_28_C96_n148, mult_28_C96_n144, mult_28_C96_n143, mult_28_C96_n142, 
      mult_28_C96_n141, mult_28_C96_n140, mult_28_C96_n139, mult_28_C96_n135, 
      mult_28_C96_n134, mult_28_C96_n133, mult_28_C96_n129, mult_28_C96_n128, 
      mult_28_C96_n127, mult_28_C96_n118, mult_28_C96_n117, mult_28_C96_n116, 
      mult_28_C96_n115, mult_28_C96_n114, mult_28_C96_n113, mult_28_C96_n112, 
      mult_28_C96_n109, mult_28_C96_n108, mult_28_C96_n107, mult_28_C96_n106, 
      mult_28_C96_n105, mult_28_C96_n104, mult_28_C96_n103, mult_28_C96_n102, 
      mult_28_C96_n101, mult_28_C96_n100, mult_28_C96_n97, mult_28_C96_n96, 
      mult_28_C96_n95, mult_28_C96_n93, mult_28_C96_n92, mult_28_C96_n87, 
      mult_28_C96_n86, mult_28_C96_n85, mult_28_C96_n84, mult_28_C96_n69, 
      mult_28_C96_n68, mult_28_C96_n67, mult_28_C96_n66, mult_28_C96_n65, 
      mult_28_C96_n63, mult_28_C96_n57, mult_28_C96_n56, mult_28_C96_n54, 
      mult_28_C96_n53, mult_28_C96_n52, mult_28_C96_n51, mult_28_C96_n48, 
      mult_28_C96_n46, mult_28_C96_n42, mult_28_C96_n40, mult_28_C96_n36, 
      mult_28_C96_n34, mult_28_C96_n30, mult_28_C96_n28, mult_28_C96_n24, 
      mult_28_C96_n22, mult_28_C96_n18, mult_28_C96_n16, mult_28_C96_n12, 
      mult_28_C96_n9, mult_28_C96_n6 : std_logic;

begin
   ready <= ready_port;
   
   coeff_memory_reg_2_1 : DFERPQ1 port map( D => data_in(1), CEB => n27, CK => 
                           clk, RB => n52, Q => coeff_memory_33_port);
   coeff_memory_reg_4_1 : DFERPQ1 port map( D => data_in(1), CEB => n26, CK => 
                           clk, RB => n51, Q => coeff_memory_1_port);
   coeff_memory_reg_3_1 : DFERPQ1 port map( D => data_in(1), CEB => n28, CK => 
                           clk, RB => n60, Q => coeff_memory_17_port);
   data_out_reg_15 : DFERPQL port map( D => y_15_port, CEB => n23, CK => clk, 
                           RB => n45, Q => data_out(15));
   z2_reg_5 : DFERPQ1 port map( D => z2_next_5_port, CEB => n23, CK => clk, RB 
                           => n47, Q => z2_5_port);
   coeff_counter_reg_0 : DFFRPQ1 port map( D => n32, CK => clk, RB => n53, Q =>
                           coeff_counter_0_port);
   coeff_counter_reg_2 : DFFRPQ1 port map( D => n30, CK => clk, RB => n60, Q =>
                           coeff_counter_2_port);
   coeff_counter_reg_1 : DFFRPQ1 port map( D => n31, CK => clk, RB => n60, Q =>
                           coeff_counter_1_port);
   z1_reg_5 : DFERPQ1 port map( D => z1_next_5_port, CEB => n23, CK => clk, RB 
                           => n50, Q => z1_5_port);
   z1_reg_4 : DFERPQ1 port map( D => z1_next_4_port, CEB => n23, CK => clk, RB 
                           => n50, Q => z1_4_port);
   z1_reg_2 : DFERPQ1 port map( D => z1_next_2_port, CEB => n23, CK => clk, RB 
                           => n50, Q => z1_2_port);
   z1_reg_3 : DFERPQ1 port map( D => z1_next_3_port, CEB => n23, CK => clk, RB 
                           => n50, Q => z1_3_port);
   z1_reg_1 : DFERPQ1 port map( D => z1_next_1_port, CEB => n23, CK => clk, RB 
                           => n50, Q => z1_1_port);
   z1_reg_0 : DFERPQ1 port map( D => z1_next_0_port, CEB => n23, CK => clk, RB 
                           => n50, Q => z1_0_port);
   ready_reg : DFFRPQ1 port map( D => n22, CK => clk, RB => n53, Q => 
                           ready_port);
   coeff_memory_reg_4_0 : DFERPQ1 port map( D => data_in(0), CEB => n26, CK => 
                           clk, RB => n51, Q => coeff_memory_0_port);
   coeff_memory_reg_3_0 : DFERPQ1 port map( D => data_in(0), CEB => n28, CK => 
                           clk, RB => n60, Q => coeff_memory_16_port);
   coeff_memory_reg_4_2 : DFERPQ1 port map( D => data_in(2), CEB => n26, CK => 
                           clk, RB => n51, Q => coeff_memory_2_port);
   coeff_memory_reg_3_2 : DFERPQ1 port map( D => data_in(2), CEB => n28, CK => 
                           clk, RB => n60, Q => coeff_memory_18_port);
   coeff_memory_reg_4_4 : DFERPQ1 port map( D => data_in(4), CEB => n26, CK => 
                           clk, RB => n51, Q => coeff_memory_4_port);
   coeff_memory_reg_3_4 : DFERPQ1 port map( D => data_in(4), CEB => n28, CK => 
                           clk, RB => n48, Q => coeff_memory_20_port);
   coeff_memory_reg_4_6 : DFERPQ1 port map( D => data_in(6), CEB => n26, CK => 
                           clk, RB => n51, Q => coeff_memory_6_port);
   coeff_memory_reg_3_6 : DFERPQ1 port map( D => data_in(6), CEB => n28, CK => 
                           clk, RB => n48, Q => coeff_memory_22_port);
   coeff_memory_reg_4_8 : DFERPQ1 port map( D => data_in(8), CEB => n26, CK => 
                           clk, RB => n52, Q => coeff_memory_8_port);
   coeff_memory_reg_4_3 : DFERPQ1 port map( D => data_in(3), CEB => n26, CK => 
                           clk, RB => n51, Q => coeff_memory_3_port);
   z2_reg_4 : DFERPQ1 port map( D => z2_next_4_port, CEB => n23, CK => clk, RB 
                           => n47, Q => z2_4_port);
   coeff_memory_reg_3_8 : DFERPQ1 port map( D => data_in(8), CEB => n28, CK => 
                           clk, RB => n48, Q => coeff_memory_24_port);
   coeff_memory_reg_3_3 : DFERPQ1 port map( D => data_in(3), CEB => n28, CK => 
                           clk, RB => n60, Q => coeff_memory_19_port);
   coeff_memory_reg_4_10 : DFERPQ1 port map( D => data_in(10), CEB => n26, CK 
                           => clk, RB => n52, Q => coeff_memory_10_port);
   coeff_memory_reg_3_10 : DFERPQ1 port map( D => data_in(10), CEB => n28, CK 
                           => clk, RB => n48, Q => coeff_memory_26_port);
   coeff_memory_reg_4_15 : DFERPQ1 port map( D => data_in(15), CEB => n26, CK 
                           => clk, RB => n52, Q => coeff_memory_15_port);
   z2_reg_3 : DFERPQ1 port map( D => z2_next_3_port, CEB => n23, CK => clk, RB 
                           => n47, Q => z2_3_port);
   coeff_memory_reg_4_5 : DFERPQ1 port map( D => data_in(5), CEB => n26, CK => 
                           clk, RB => n51, Q => coeff_memory_5_port);
   coeff_memory_reg_4_12 : DFERPQ1 port map( D => data_in(12), CEB => n26, CK 
                           => clk, RB => n52, Q => coeff_memory_12_port);
   coeff_memory_reg_3_15 : DFERPQ1 port map( D => data_in(15), CEB => n28, CK 
                           => clk, RB => n48, Q => coeff_memory_31_port);
   z2_reg_2 : DFERPQ1 port map( D => z2_next_2_port, CEB => n23, CK => clk, RB 
                           => n47, Q => z2_2_port);
   coeff_memory_reg_3_12 : DFERPQ1 port map( D => data_in(12), CEB => n28, CK 
                           => clk, RB => n48, Q => coeff_memory_28_port);
   coeff_memory_reg_3_5 : DFERPQ1 port map( D => data_in(5), CEB => n28, CK => 
                           clk, RB => n48, Q => coeff_memory_21_port);
   coeff_memory_reg_4_14 : DFERPQ1 port map( D => data_in(14), CEB => n26, CK 
                           => clk, RB => n52, Q => coeff_memory_14_port);
   coeff_memory_reg_3_14 : DFERPQ1 port map( D => data_in(14), CEB => n28, CK 
                           => clk, RB => n48, Q => coeff_memory_30_port);
   coeff_memory_reg_3_7 : DFERPQ1 port map( D => data_in(7), CEB => n28, CK => 
                           clk, RB => n48, Q => coeff_memory_23_port);
   z2_reg_1 : DFERPQ1 port map( D => z2_next_1_port, CEB => n23, CK => clk, RB 
                           => n47, Q => z2_1_port);
   coeff_memory_reg_4_9 : DFERPQ1 port map( D => data_in(9), CEB => n26, CK => 
                           clk, RB => n52, Q => coeff_memory_9_port);
   coeff_memory_reg_3_9 : DFERPQ1 port map( D => data_in(9), CEB => n28, CK => 
                           clk, RB => n48, Q => coeff_memory_25_port);
   z2_reg_0 : DFERPQ1 port map( D => z2_next_0_port, CEB => n23, CK => clk, RB 
                           => n47, Q => z2_0_port);
   coeff_memory_reg_4_11 : DFERPQ1 port map( D => data_in(11), CEB => n26, CK 
                           => clk, RB => n52, Q => coeff_memory_11_port);
   coeff_memory_reg_2_15 : DFERPQ1 port map( D => data_in(15), CEB => n27, CK 
                           => clk, RB => n53, Q => coeff_memory_47_port);
   coeff_memory_reg_3_11 : DFERPQ1 port map( D => data_in(11), CEB => n28, CK 
                           => clk, RB => n48, Q => coeff_memory_27_port);
   coeff_memory_reg_4_13 : DFERPQ1 port map( D => data_in(13), CEB => n26, CK 
                           => clk, RB => n52, Q => coeff_memory_13_port);
   coeff_memory_reg_3_13 : DFERPQ1 port map( D => data_in(13), CEB => n28, CK 
                           => clk, RB => n48, Q => coeff_memory_29_port);
   coeff_memory_reg_2_0 : DFERPQ1 port map( D => data_in(0), CEB => n27, CK => 
                           clk, RB => n52, Q => coeff_memory_32_port);
   coeff_memory_reg_2_14 : DFERPQ1 port map( D => data_in(14), CEB => n27, CK 
                           => clk, RB => n53, Q => coeff_memory_46_port);
   coeff_memory_reg_2_12 : DFERPQ1 port map( D => data_in(12), CEB => n27, CK 
                           => clk, RB => n53, Q => coeff_memory_44_port);
   coeff_memory_reg_2_4 : DFERPQ1 port map( D => data_in(4), CEB => n27, CK => 
                           clk, RB => n52, Q => coeff_memory_36_port);
   coeff_memory_reg_2_13 : DFERPQ1 port map( D => data_in(13), CEB => n27, CK 
                           => clk, RB => n53, Q => coeff_memory_45_port);
   coeff_memory_reg_2_11 : DFERPQ1 port map( D => data_in(11), CEB => n27, CK 
                           => clk, RB => n53, Q => coeff_memory_43_port);
   coeff_memory_reg_2_8 : DFERPQ1 port map( D => data_in(8), CEB => n27, CK => 
                           clk, RB => n53, Q => coeff_memory_40_port);
   coeff_memory_reg_2_2 : DFERPQ1 port map( D => data_in(2), CEB => n27, CK => 
                           clk, RB => n52, Q => coeff_memory_34_port);
   coeff_memory_reg_2_10 : DFERPQ1 port map( D => data_in(10), CEB => n27, CK 
                           => clk, RB => n53, Q => coeff_memory_42_port);
   coeff_memory_reg_2_6 : DFERPQ1 port map( D => data_in(6), CEB => n27, CK => 
                           clk, RB => n53, Q => coeff_memory_38_port);
   coeff_memory_reg_2_7 : DFERPQ1 port map( D => data_in(7), CEB => n27, CK => 
                           clk, RB => n53, Q => coeff_memory_39_port);
   coeff_memory_reg_2_3 : DFERPQ1 port map( D => data_in(3), CEB => n27, CK => 
                           clk, RB => n52, Q => coeff_memory_35_port);
   coeff_memory_reg_2_9 : DFERPQ1 port map( D => data_in(9), CEB => n27, CK => 
                           clk, RB => n53, Q => coeff_memory_41_port);
   coeff_memory_reg_2_5 : DFERPQ1 port map( D => data_in(5), CEB => n27, CK => 
                           clk, RB => n53, Q => coeff_memory_37_port);
   coeff_memory_reg_1_15 : DFERPQ1 port map( D => data_in(15), CEB => n29, CK 
                           => clk, RB => n50, Q => coeff_memory_63_port);
   coeff_memory_reg_1_0 : DFERPQ1 port map( D => data_in(0), CEB => n29, CK => 
                           clk, RB => n48, Q => coeff_memory_48_port);
   coeff_memory_reg_1_14 : DFERPQ1 port map( D => data_in(14), CEB => n29, CK 
                           => clk, RB => n50, Q => coeff_memory_62_port);
   coeff_memory_reg_1_12 : DFERPQ1 port map( D => data_in(12), CEB => n29, CK 
                           => clk, RB => n49, Q => coeff_memory_60_port);
   coeff_memory_reg_1_4 : DFERPQ1 port map( D => data_in(4), CEB => n29, CK => 
                           clk, RB => n49, Q => coeff_memory_52_port);
   coeff_memory_reg_1_13 : DFERPQ1 port map( D => data_in(13), CEB => n29, CK 
                           => clk, RB => n49, Q => coeff_memory_61_port);
   coeff_memory_reg_1_11 : DFERPQ1 port map( D => data_in(11), CEB => n29, CK 
                           => clk, RB => n49, Q => coeff_memory_59_port);
   coeff_memory_reg_1_8 : DFERPQ1 port map( D => data_in(8), CEB => n29, CK => 
                           clk, RB => n49, Q => coeff_memory_56_port);
   coeff_memory_reg_1_2 : DFERPQ1 port map( D => data_in(2), CEB => n29, CK => 
                           clk, RB => n49, Q => coeff_memory_50_port);
   coeff_memory_reg_1_10 : DFERPQ1 port map( D => data_in(10), CEB => n29, CK 
                           => clk, RB => n49, Q => coeff_memory_58_port);
   coeff_memory_reg_1_6 : DFERPQ1 port map( D => data_in(6), CEB => n29, CK => 
                           clk, RB => n49, Q => coeff_memory_54_port);
   coeff_memory_reg_1_7 : DFERPQ1 port map( D => data_in(7), CEB => n29, CK => 
                           clk, RB => n49, Q => coeff_memory_55_port);
   coeff_memory_reg_1_1 : DFERPQ1 port map( D => data_in(1), CEB => n29, CK => 
                           clk, RB => n49, Q => coeff_memory_49_port);
   coeff_memory_reg_1_3 : DFERPQ1 port map( D => data_in(3), CEB => n29, CK => 
                           clk, RB => n49, Q => coeff_memory_51_port);
   coeff_memory_reg_1_9 : DFERPQ1 port map( D => data_in(9), CEB => n29, CK => 
                           clk, RB => n49, Q => coeff_memory_57_port);
   coeff_memory_reg_1_5 : DFERPQ1 port map( D => data_in(5), CEB => n29, CK => 
                           clk, RB => n49, Q => coeff_memory_53_port);
   coeff_memory_reg_0_0 : DFERPQ1 port map( D => data_in(0), CEB => n25, CK => 
                           clk, RB => n46, Q => coeff_memory_64_port);
   coeff_memory_reg_0_14 : DFERPQ1 port map( D => data_in(14), CEB => n25, CK 
                           => clk, RB => n47, Q => coeff_memory_78_port);
   coeff_memory_reg_0_10 : DFERPQ1 port map( D => data_in(10), CEB => n25, CK 
                           => clk, RB => n47, Q => coeff_memory_74_port);
   coeff_memory_reg_0_8 : DFERPQ1 port map( D => data_in(8), CEB => n25, CK => 
                           clk, RB => n46, Q => coeff_memory_72_port);
   coeff_memory_reg_0_6 : DFERPQ1 port map( D => data_in(6), CEB => n25, CK => 
                           clk, RB => n46, Q => coeff_memory_70_port);
   coeff_memory_reg_0_4 : DFERPQ1 port map( D => data_in(4), CEB => n25, CK => 
                           clk, RB => n46, Q => coeff_memory_68_port);
   coeff_memory_reg_0_2 : DFERPQ1 port map( D => data_in(2), CEB => n25, CK => 
                           clk, RB => n46, Q => coeff_memory_66_port);
   coeff_memory_reg_0_12 : DFERPQ1 port map( D => data_in(12), CEB => n25, CK 
                           => clk, RB => n47, Q => coeff_memory_76_port);
   data_out_reg_14 : DFERPQL port map( D => y_14_port, CEB => n23, CK => clk, 
                           RB => n45, Q => data_out(14));
   data_out_reg_13 : DFERPQL port map( D => y_13_port, CEB => n23, CK => clk, 
                           RB => n45, Q => data_out(13));
   data_out_reg_12 : DFERPQL port map( D => y_12_port, CEB => n23, CK => clk, 
                           RB => n45, Q => data_out(12));
   data_out_reg_11 : DFERPQL port map( D => y_11_port, CEB => n23, CK => clk, 
                           RB => n45, Q => data_out(11));
   data_out_reg_10 : DFERPQL port map( D => n42, CEB => n23, CK => clk, RB => 
                           n45, Q => data_out(10));
   data_out_reg_9 : DFERPQL port map( D => y_9_port, CEB => n23, CK => clk, RB 
                           => n45, Q => data_out(9));
   data_out_reg_8 : DFERPQL port map( D => y_8_port, CEB => n23, CK => clk, RB 
                           => n45, Q => data_out(8));
   data_out_reg_7 : DFERPQL port map( D => y_7_port, CEB => n23, CK => clk, RB 
                           => n45, Q => data_out(7));
   data_out_reg_6 : DFERPQL port map( D => y_6_port, CEB => n23, CK => clk, RB 
                           => n45, Q => data_out(6));
   data_out_reg_5 : DFERPQL port map( D => n38, CEB => n23, CK => clk, RB => 
                           n45, Q => data_out(5));
   data_out_reg_3 : DFERPQL port map( D => y_3_port, CEB => n23, CK => clk, RB 
                           => n45, Q => data_out(3));
   data_out_reg_1 : DFERPQL port map( D => n36, CEB => n23, CK => clk, RB => 
                           n46, Q => data_out(1));
   data_out_reg_0 : DFERPQ1 port map( D => n39, CEB => n23, CK => clk, RB => 
                           n46, Q => data_out(0));
   data_out_reg_4 : DFERPQ1 port map( D => n44, CEB => n23, CK => clk, RB => 
                           n45, Q => data_out(4));
   data_out_reg_2 : DFERPQL port map( D => n43, CEB => n23, CK => clk, RB => 
                           n46, Q => data_out(2));
   z1_reg_15 : DFERPQ1 port map( D => z1_next_15_port, CEB => n23, CK => clk, 
                           RB => n60, Q => z1_15_port);
   z1_reg_14 : DFERPQ1 port map( D => z1_next_14_port, CEB => n23, CK => clk, 
                           RB => n60, Q => z1_14_port);
   z1_reg_13 : DFERPQ1 port map( D => z1_next_13_port, CEB => n23, CK => clk, 
                           RB => n60, Q => z1_13_port);
   z1_reg_12 : DFERPQ1 port map( D => z1_next_12_port, CEB => n23, CK => clk, 
                           RB => n60, Q => z1_12_port);
   z1_reg_8 : DFERPQ1 port map( D => z1_next_8_port, CEB => n23, CK => clk, RB 
                           => n60, Q => z1_8_port);
   z1_reg_11 : DFERPQ1 port map( D => z1_next_11_port, CEB => n23, CK => clk, 
                           RB => n60, Q => z1_11_port);
   z1_reg_10 : DFERPQ1 port map( D => z1_next_10_port, CEB => n23, CK => clk, 
                           RB => n60, Q => z1_10_port);
   z1_reg_9 : DFERPQ1 port map( D => z1_next_9_port, CEB => n23, CK => clk, RB 
                           => n60, Q => z1_9_port);
   z1_reg_7 : DFERPQ1 port map( D => z1_next_7_port, CEB => n23, CK => clk, RB 
                           => n60, Q => z1_7_port);
   z1_reg_6 : DFERPQ1 port map( D => z1_next_6_port, CEB => n23, CK => clk, RB 
                           => n60, Q => z1_6_port);
   z2_reg_15 : DFERPQ1 port map( D => z2_next_15_port, CEB => n23, CK => clk, 
                           RB => n60, Q => z2_15_port);
   z2_reg_14 : DFERPQ1 port map( D => z2_next_14_port, CEB => n23, CK => clk, 
                           RB => n60, Q => z2_14_port);
   z2_reg_10 : DFERPQ1 port map( D => z2_next_10_port, CEB => n23, CK => clk, 
                           RB => n60, Q => z2_10_port);
   z2_reg_12 : DFERPQ1 port map( D => z2_next_12_port, CEB => n23, CK => clk, 
                           RB => n60, Q => z2_12_port);
   z2_reg_11 : DFERPQ1 port map( D => z2_next_11_port, CEB => n23, CK => clk, 
                           RB => n60, Q => z2_11_port);
   z2_reg_13 : DFERPQ1 port map( D => z2_next_13_port, CEB => n23, CK => clk, 
                           RB => n60, Q => z2_13_port);
   z2_reg_8 : DFERPQ1 port map( D => z2_next_8_port, CEB => n23, CK => clk, RB 
                           => n60, Q => z2_8_port);
   z2_reg_7 : DFERPQ1 port map( D => z2_next_7_port, CEB => n23, CK => clk, RB 
                           => n60, Q => z2_7_port);
   z2_reg_9 : DFERPQ1 port map( D => z2_next_9_port, CEB => n23, CK => clk, RB 
                           => n60, Q => z2_9_port);
   z2_reg_6 : DFERPQ1 port map( D => z2_next_6_port, CEB => n23, CK => clk, RB 
                           => n60, Q => z2_6_port);
   coeff_memory_reg_0_1 : DFERPQ4 port map( D => data_in(1), CEB => n25, CK => 
                           clk, RB => n46, Q => coeff_memory_65_port);
   coeff_memory_reg_0_11 : DFERPQ2 port map( D => data_in(11), CEB => n25, CK 
                           => clk, RB => n47, Q => coeff_memory_75_port);
   coeff_memory_reg_0_5 : DFERPQ4 port map( D => data_in(5), CEB => n25, CK => 
                           clk, RB => n46, Q => coeff_memory_69_port);
   coeff_memory_reg_0_7 : DFERPQ4 port map( D => data_in(7), CEB => n25, CK => 
                           clk, RB => n46, Q => coeff_memory_71_port);
   coeff_memory_reg_0_3 : DFERPQ4 port map( D => data_in(3), CEB => n25, CK => 
                           clk, RB => n46, Q => coeff_memory_67_port);
   coeff_memory_reg_0_13 : DFERPQ2 port map( D => data_in(13), CEB => n25, CK 
                           => clk, RB => n47, Q => coeff_memory_77_port);
   coeff_memory_reg_4_7 : DFERPQL port map( D => data_in(7), CEB => n26, CK => 
                           clk, RB => n60, Q => coeff_memory_7_port);
   coeff_memory_reg_0_9 : DFERPQ4 port map( D => data_in(9), CEB => n25, CK => 
                           clk, RB => n46, Q => coeff_memory_73_port);
   coeff_memory_reg_0_15 : DFERPQ1 port map( D => data_in(15), CEB => n25, CK 
                           => clk, RB => n60, Q => coeff_memory_79_port);
   U21 : INVD4 port map( A => n35, Z => n36);
   U22 : INVD4 port map( A => n35, Z => n34);
   U23 : INVD4 port map( A => n37, Z => n33);
   U24 : INVBD4 port map( A => y_5_port, Z => n37);
   U25 : INVD4 port map( A => y_1_port, Z => n35);
   U26 : BUFD4 port map( A => y_10_port, Z => n42);
   U27 : INVD4 port map( A => n37, Z => n38);
   U28 : BUFD8 port map( A => y_0_port, Z => n39);
   U29 : INVD1 port map( A => n56, Z => n59);
   U30 : INVD1 port map( A => reset, Z => n46);
   U31 : INVD1 port map( A => reset, Z => n52);
   U32 : INVD1 port map( A => n54, Z => n48);
   U33 : INVD1 port map( A => reset, Z => n49);
   U34 : INVD1 port map( A => n54, Z => n53);
   U35 : INVD1 port map( A => n54, Z => n45);
   U36 : INVD1 port map( A => n54, Z => n47);
   U37 : INVD1 port map( A => n54, Z => n51);
   U38 : INVD1 port map( A => reset, Z => n50);
   U39 : NAN3D1 port map( A1 => n59, A2 => n58, A3 => n57, Z => n25);
   U40 : OA21D1 port map( A1 => n57, A2 => n58, B => n23, Z => n40);
   U41 : NAN2D1 port map( A1 => n41, A2 => n58, Z => n29);
   U42 : INVD1 port map( A => n60, Z => n54);
   U43 : INVD1 port map( A => coeff_counter_1_port, Z => n58);
   U44 : NAN2D1 port map( A1 => coeff_counter_2_port, A2 => n59, Z => n26);
   U45 : NAN2D1 port map( A1 => coeff_counter_1_port, A2 => n59, Z => n27);
   U46 : NAN2D1 port map( A1 => n41, A2 => coeff_counter_1_port, Z => n28);
   U47 : AND2D1 port map( A1 => n40, A2 => coeff_counter_0_port, Z => n41);
   U48 : INVD1 port map( A => coeff_counter_2_port, Z => n57);
   U49 : NAN2M1D1 port map( A1 => ready_port, A2 => n23, Z => n22);
   U50 : INVD1 port map( A => coeff_counter_0_port, Z => n55);
   U51 : INVD1 port map( A => reset, Z => n60);
   U52 : TIEHI port map( Z => req);
   U53 : TIELO port map( Z => n61);
   U54 : BUFD4 port map( A => y_2_port, Z => n43);
   U55 : BUFDL port map( A => y_4_port, Z => n44);
   U56 : NAN3D1 port map( A1 => coeff_counter_2_port, A2 => 
                           coeff_counter_0_port, A3 => n58, Z => n23);
   U57 : OAI21D1 port map( A1 => n41, A2 => n58, B => n29, Z => n31);
   U58 : NAN2D1 port map( A1 => n57, A2 => n28, Z => n30);
   U59 : NAN2D1 port map( A1 => n40, A2 => n55, Z => n56);
   U60 : OAI21D1 port map( A1 => n40, A2 => n55, B => n56, Z => n32);
   mult_28_C94_U1004 : BUFD1 port map( A => coeff_memory_47_port, Z => 
                           mult_28_C94_n43);
   mult_28_C94_U1003 : BUFD1 port map( A => coeff_memory_45_port, Z => 
                           mult_28_C94_n37);
   mult_28_C94_U1002 : BUFD1 port map( A => coeff_memory_35_port, Z => 
                           mult_28_C94_n7);
   mult_28_C94_U1001 : BUFD1 port map( A => coeff_memory_41_port, Z => 
                           mult_28_C94_n25);
   mult_28_C94_U1000 : BUFD1 port map( A => coeff_memory_37_port, Z => 
                           mult_28_C94_n13);
   mult_28_C94_U999 : BUFD1 port map( A => coeff_memory_43_port, Z => 
                           mult_28_C94_n31);
   mult_28_C94_U998 : BUFD1 port map( A => coeff_memory_39_port, Z => 
                           mult_28_C94_n19);
   mult_28_C94_U997 : BUFD1 port map( A => coeff_memory_33_port, Z => 
                           mult_28_C94_n1);
   mult_28_C94_U996 : INVD1 port map( A => coeff_memory_32_port, Z => 
                           mult_28_C94_n834);
   mult_28_C94_U995 : NAN2D1 port map( A1 => mult_28_C94_n818, A2 => 
                           mult_28_C94_n834, Z => mult_28_C94_n826);
   mult_28_C94_U994 : NAN2D1 port map( A1 => mult_28_C94_n811, A2 => 
                           mult_28_C94_n827, Z => mult_28_C94_n819);
   mult_28_C94_U993 : NAN2D1 port map( A1 => mult_28_C94_n812, A2 => 
                           mult_28_C94_n828, Z => mult_28_C94_n820);
   mult_28_C94_U992 : NAN2D1 port map( A1 => mult_28_C94_n814, A2 => 
                           mult_28_C94_n830, Z => mult_28_C94_n822);
   mult_28_C94_U991 : NAN2D1 port map( A1 => mult_28_C94_n816, A2 => 
                           mult_28_C94_n832, Z => mult_28_C94_n824);
   mult_28_C94_U990 : NAN2D1 port map( A1 => mult_28_C94_n813, A2 => 
                           mult_28_C94_n829, Z => mult_28_C94_n821);
   mult_28_C94_U989 : NAN2D1 port map( A1 => mult_28_C94_n815, A2 => 
                           mult_28_C94_n831, Z => mult_28_C94_n823);
   mult_28_C94_U988 : NAN2D1 port map( A1 => mult_28_C94_n817, A2 => 
                           mult_28_C94_n833, Z => mult_28_C94_n825);
   mult_28_C94_U987 : OAI22M10D1 port map( A1 => mult_28_C94_n7, A2 => 
                           mult_28_C94_n12, B1 => mult_28_C94_n10, B2 => 
                           mult_28_C94_n777, Z => mult_28_C94_n529);
   mult_28_C94_U986 : ADHALFDL port map( A => mult_28_C94_n641, B => 
                           mult_28_C94_n656, CO => mult_28_C94_n521, S => 
                           mult_28_C94_n522);
   mult_28_C94_U985 : BUFD1 port map( A => data_in(13), Z => mult_28_C94_n797);
   mult_28_C94_U984 : BUFD1 port map( A => data_in(12), Z => mult_28_C94_n798);
   mult_28_C94_U983 : BUFD1 port map( A => data_in(14), Z => mult_28_C94_n796);
   mult_28_C94_U982 : BUFD1 port map( A => data_in(15), Z => mult_28_C94_n795);
   mult_28_C94_U981 : BUFD1 port map( A => data_in(11), Z => mult_28_C94_n799);
   mult_28_C94_U980 : BUFD1 port map( A => data_in(3), Z => mult_28_C94_n807);
   mult_28_C94_U979 : BUFD1 port map( A => data_in(2), Z => mult_28_C94_n808);
   mult_28_C94_U978 : BUFD1 port map( A => data_in(8), Z => mult_28_C94_n802);
   mult_28_C94_U977 : BUFD1 port map( A => data_in(7), Z => mult_28_C94_n803);
   mult_28_C94_U976 : BUFD1 port map( A => data_in(4), Z => mult_28_C94_n806);
   mult_28_C94_U975 : BUFD1 port map( A => data_in(1), Z => mult_28_C94_n809);
   mult_28_C94_U974 : INVD1 port map( A => mult_28_C94_n1, Z => 
                           mult_28_C94_n842);
   mult_28_C94_U973 : BUFD1 port map( A => mult_28_C94_n834, Z => 
                           mult_28_C94_n3);
   mult_28_C94_U972 : BUFD1 port map( A => mult_28_C94_n834, Z => 
                           mult_28_C94_n4);
   mult_28_C94_U971 : BUFD1 port map( A => mult_28_C94_n832, Z => 
                           mult_28_C94_n16);
   mult_28_C94_U970 : OA22D1 port map( A1 => mult_28_C94_n46, A2 => 
                           mult_28_C94_n659, B1 => mult_28_C94_n48, B2 => 
                           mult_28_C94_n660, Z => mult_28_C94_n940);
   mult_28_C94_U969 : BUFD1 port map( A => mult_28_C94_n827, Z => 
                           mult_28_C94_n46);
   mult_28_C94_U968 : BUFD1 port map( A => mult_28_C94_n828, Z => 
                           mult_28_C94_n40);
   mult_28_C94_U967 : BUFD1 port map( A => mult_28_C94_n827, Z => 
                           mult_28_C94_n45);
   mult_28_C94_U966 : BUFD1 port map( A => mult_28_C94_n828, Z => 
                           mult_28_C94_n39);
   mult_28_C94_U965 : BUFD1 port map( A => mult_28_C94_n826, Z => 
                           mult_28_C94_n5);
   mult_28_C94_U964 : BUFD1 port map( A => mult_28_C94_n826, Z => 
                           mult_28_C94_n6);
   mult_28_C94_U963 : BUFD1 port map( A => mult_28_C94_n829, Z => 
                           mult_28_C94_n34);
   mult_28_C94_U962 : BUFD1 port map( A => mult_28_C94_n830, Z => 
                           mult_28_C94_n28);
   mult_28_C94_U961 : BUFD1 port map( A => mult_28_C94_n831, Z => 
                           mult_28_C94_n22);
   mult_28_C94_U960 : BUFD1 port map( A => mult_28_C94_n830, Z => 
                           mult_28_C94_n27);
   mult_28_C94_U959 : BUFD1 port map( A => mult_28_C94_n832, Z => 
                           mult_28_C94_n15);
   mult_28_C94_U958 : BUFD1 port map( A => mult_28_C94_n829, Z => 
                           mult_28_C94_n33);
   mult_28_C94_U957 : BUFD1 port map( A => mult_28_C94_n833, Z => 
                           mult_28_C94_n9);
   mult_28_C94_U956 : BUFD1 port map( A => mult_28_C94_n831, Z => 
                           mult_28_C94_n21);
   mult_28_C94_U955 : BUFD1 port map( A => mult_28_C94_n833, Z => 
                           mult_28_C94_n10);
   mult_28_C94_U954 : BUFD1 port map( A => mult_28_C94_n824, Z => 
                           mult_28_C94_n18);
   mult_28_C94_U953 : BUFD1 port map( A => mult_28_C94_n820, Z => 
                           mult_28_C94_n42);
   mult_28_C94_U952 : BUFD1 port map( A => mult_28_C94_n819, Z => 
                           mult_28_C94_n47);
   mult_28_C94_U951 : BUFD1 port map( A => mult_28_C94_n819, Z => 
                           mult_28_C94_n48);
   mult_28_C94_U950 : BUFD1 port map( A => mult_28_C94_n820, Z => 
                           mult_28_C94_n41);
   mult_28_C94_U949 : BUFD1 port map( A => mult_28_C94_n821, Z => 
                           mult_28_C94_n36);
   mult_28_C94_U948 : BUFD1 port map( A => mult_28_C94_n822, Z => 
                           mult_28_C94_n30);
   mult_28_C94_U947 : BUFD1 port map( A => mult_28_C94_n822, Z => 
                           mult_28_C94_n29);
   mult_28_C94_U946 : BUFD1 port map( A => mult_28_C94_n823, Z => 
                           mult_28_C94_n24);
   mult_28_C94_U945 : BUFD1 port map( A => mult_28_C94_n824, Z => 
                           mult_28_C94_n17);
   mult_28_C94_U944 : BUFD1 port map( A => mult_28_C94_n821, Z => 
                           mult_28_C94_n35);
   mult_28_C94_U943 : BUFD1 port map( A => mult_28_C94_n825, Z => 
                           mult_28_C94_n11);
   mult_28_C94_U942 : BUFD1 port map( A => mult_28_C94_n823, Z => 
                           mult_28_C94_n23);
   mult_28_C94_U941 : BUFD1 port map( A => mult_28_C94_n825, Z => 
                           mult_28_C94_n12);
   mult_28_C94_U940 : AND2D1 port map( A1 => mult_28_C94_n658, A2 => 
                           mult_28_C94_n530, Z => mult_28_C94_n939);
   mult_28_C94_U939 : AND2DL port map( A1 => mult_28_C94_n657, A2 => 
                           mult_28_C94_n642, Z => mult_28_C94_n938);
   mult_28_C94_U938 : OR2D1 port map( A1 => mult_28_C94_n657, A2 => 
                           mult_28_C94_n642, Z => mult_28_C94_n937);
   mult_28_C94_U937 : NOR2D1 port map( A1 => mult_28_C94_n522, A2 => 
                           mult_28_C94_n529, Z => mult_28_C94_n275);
   mult_28_C94_U936 : OAI22M10D1 port map( A1 => mult_28_C94_n37, A2 => 
                           mult_28_C94_n42, B1 => mult_28_C94_n40, B2 => 
                           mult_28_C94_n692, Z => mult_28_C94_n524);
   mult_28_C94_U935 : INVD1 port map( A => mult_28_C94_n13, Z => 
                           mult_28_C94_n840);
   mult_28_C94_U934 : ADHALFDL port map( A => mult_28_C94_n528, B => 
                           mult_28_C94_n654, CO => mult_28_C94_n517, S => 
                           mult_28_C94_n518);
   mult_28_C94_U933 : AND2DL port map( A1 => mult_28_C94_n520, A2 => 
                           mult_28_C94_n521, Z => mult_28_C94_n936);
   mult_28_C94_U932 : OAI22M10D1 port map( A1 => mult_28_C94_n43, A2 => 
                           mult_28_C94_n48, B1 => mult_28_C94_n46, B2 => 
                           mult_28_C94_n675, Z => mult_28_C94_n523);
   mult_28_C94_U931 : OR2D1 port map( A1 => mult_28_C94_n520, A2 => 
                           mult_28_C94_n521, Z => mult_28_C94_n935);
   mult_28_C94_U930 : NAN2DL port map( A1 => mult_28_C94_n516, A2 => 
                           mult_28_C94_n519, Z => mult_28_C94_n268);
   mult_28_C94_U929 : INVD1 port map( A => mult_28_C94_n31, Z => 
                           mult_28_C94_n837);
   mult_28_C94_U928 : ADHALFDL port map( A => mult_28_C94_n525, B => 
                           mult_28_C94_n648, CO => mult_28_C94_n481, S => 
                           mult_28_C94_n482);
   mult_28_C94_U927 : INVD1 port map( A => mult_28_C94_n25, Z => 
                           mult_28_C94_n838);
   mult_28_C94_U926 : ADHALFDL port map( A => mult_28_C94_n526, B => 
                           mult_28_C94_n650, CO => mult_28_C94_n497, S => 
                           mult_28_C94_n498);
   mult_28_C94_U925 : OR2D1 port map( A1 => mult_28_C94_n512, A2 => 
                           mult_28_C94_n515, Z => mult_28_C94_n933);
   mult_28_C94_U924 : INVD1 port map( A => mult_28_C94_n19, Z => 
                           mult_28_C94_n839);
   mult_28_C94_U923 : ADHALFDL port map( A => mult_28_C94_n527, B => 
                           mult_28_C94_n652, CO => mult_28_C94_n509, S => 
                           mult_28_C94_n510);
   mult_28_C94_U922 : OR2D1 port map( A1 => mult_28_C94_n315, A2 => 
                           mult_28_C94_n940, Z => mult_28_C94_n932);
   mult_28_C94_U921 : AO21D1 port map( A1 => mult_28_C94_n42, A2 => 
                           mult_28_C94_n40, B => mult_28_C94_n676, Z => 
                           mult_28_C94_n547);
   mult_28_C94_U920 : INVD1 port map( A => mult_28_C94_n319, Z => 
                           mult_28_C94_n320);
   mult_28_C94_U919 : AO21D1 port map( A1 => mult_28_C94_n36, A2 => 
                           mult_28_C94_n34, B => mult_28_C94_n693, Z => 
                           mult_28_C94_n563);
   mult_28_C94_U918 : AO21D1 port map( A1 => mult_28_C94_n30, A2 => 
                           mult_28_C94_n28, B => mult_28_C94_n710, Z => 
                           mult_28_C94_n579);
   mult_28_C94_U917 : INVDL port map( A => mult_28_C94_n329, Z => 
                           mult_28_C94_n330);
   mult_28_C94_U916 : INVDL port map( A => mult_28_C94_n361, Z => 
                           mult_28_C94_n362);
   mult_28_C94_U915 : AO21D1 port map( A1 => mult_28_C94_n24, A2 => 
                           mult_28_C94_n22, B => mult_28_C94_n727, Z => 
                           mult_28_C94_n595);
   mult_28_C94_U914 : NAN2D1 port map( A1 => mult_28_C94_n315, A2 => 
                           mult_28_C94_n940, Z => mult_28_C94_n84);
   mult_28_C94_U913 : NAN2D1 port map( A1 => mult_28_C94_n932, A2 => 
                           mult_28_C94_n84, Z => mult_28_C94_n54);
   mult_28_C94_U912 : AO21D1 port map( A1 => mult_28_C94_n18, A2 => 
                           mult_28_C94_n16, B => mult_28_C94_n744, Z => 
                           mult_28_C94_n611);
   mult_28_C94_U911 : AO21D1 port map( A1 => mult_28_C94_n6, A2 => 
                           mult_28_C94_n4, B => mult_28_C94_n778, Z => 
                           mult_28_C94_n643);
   mult_28_C94_U910 : EXNOR2D1 port map( A1 => mult_28_C94_n600, A2 => 
                           mult_28_C94_n558, Z => mult_28_C94_n424);
   mult_28_C94_U909 : AO21D1 port map( A1 => mult_28_C94_n12, A2 => 
                           mult_28_C94_n10, B => mult_28_C94_n761, Z => 
                           mult_28_C94_n627);
   mult_28_C94_U908 : INVDL port map( A => mult_28_C94_n383, Z => 
                           mult_28_C94_n384);
   mult_28_C94_U907 : AND2DL port map( A1 => mult_28_C94_n492, A2 => 
                           mult_28_C94_n499, Z => mult_28_C94_n931);
   mult_28_C94_U906 : OR2D1 port map( A1 => mult_28_C94_n506, A2 => 
                           mult_28_C94_n511, Z => mult_28_C94_n930);
   mult_28_C94_U905 : AND2D1 port map( A1 => mult_28_C94_n506, A2 => 
                           mult_28_C94_n511, Z => mult_28_C94_n929);
   mult_28_C94_U904 : OR2D1 port map( A1 => mult_28_C94_n492, A2 => 
                           mult_28_C94_n499, Z => mult_28_C94_n928);
   mult_28_C94_U903 : AND2DL port map( A1 => mult_28_C94_n500, A2 => 
                           mult_28_C94_n505, Z => mult_28_C94_n927);
   mult_28_C94_U902 : OR2D1 port map( A1 => mult_28_C94_n500, A2 => 
                           mult_28_C94_n505, Z => mult_28_C94_n926);
   mult_28_C94_U901 : NAN2D1 port map( A1 => mult_28_C94_n926, A2 => 
                           mult_28_C94_n930, Z => mult_28_C94_n249);
   mult_28_C94_U900 : NAN2D1 port map( A1 => mult_28_C94_n317, A2 => 
                           mult_28_C94_n316, Z => mult_28_C94_n93);
   mult_28_C94_U899 : NOR2D1 port map( A1 => mult_28_C94_n317, A2 => 
                           mult_28_C94_n316, Z => mult_28_C94_n92);
   mult_28_C94_U898 : NAN2D1 port map( A1 => mult_28_C94_n318, A2 => 
                           mult_28_C94_n321, Z => mult_28_C94_n104);
   mult_28_C94_U897 : NOR2D1 port map( A1 => mult_28_C94_n318, A2 => 
                           mult_28_C94_n321, Z => mult_28_C94_n103);
   mult_28_C94_U896 : NAN2D1 port map( A1 => mult_28_C94_n325, A2 => 
                           mult_28_C94_n322, Z => mult_28_C94_n113);
   mult_28_C94_U895 : NOR2D1 port map( A1 => mult_28_C94_n325, A2 => 
                           mult_28_C94_n322, Z => mult_28_C94_n112);
   mult_28_C94_U894 : INVDL port map( A => mult_28_C94_n343, Z => 
                           mult_28_C94_n344);
   mult_28_C94_U893 : NAN2D1 port map( A1 => mult_28_C94_n925, A2 => 
                           mult_28_C94_n918, Z => mult_28_C94_n216);
   mult_28_C94_U892 : OR2D1 port map( A1 => mult_28_C94_n452, A2 => 
                           mult_28_C94_n463, Z => mult_28_C94_n925);
   mult_28_C94_U891 : AND2DL port map( A1 => mult_28_C94_n474, A2 => 
                           mult_28_C94_n483, Z => mult_28_C94_n924);
   mult_28_C94_U890 : OR2D1 port map( A1 => mult_28_C94_n484, A2 => 
                           mult_28_C94_n491, Z => mult_28_C94_n922);
   mult_28_C94_U889 : OR2D1 port map( A1 => mult_28_C94_n474, A2 => 
                           mult_28_C94_n483, Z => mult_28_C94_n921);
   mult_28_C94_U888 : INVD1 port map( A => mult_28_C94_n112, Z => 
                           mult_28_C94_n110);
   mult_28_C94_U887 : NOR2D1 port map( A1 => mult_28_C94_n112, A2 => 
                           mult_28_C94_n103, Z => mult_28_C94_n101);
   mult_28_C94_U886 : NAN2DL port map( A1 => mult_28_C94_n326, A2 => 
                           mult_28_C94_n331, Z => mult_28_C94_n126);
   mult_28_C94_U885 : OR2D1 port map( A1 => mult_28_C94_n99, A2 => 
                           mult_28_C94_n92, Z => mult_28_C94_n920);
   mult_28_C94_U884 : NOR2D1 port map( A1 => mult_28_C94_n326, A2 => 
                           mult_28_C94_n331, Z => mult_28_C94_n125);
   mult_28_C94_U883 : NAN2D1 port map( A1 => mult_28_C94_n332, A2 => 
                           mult_28_C94_n337, Z => mult_28_C94_n133);
   mult_28_C94_U882 : INVDL port map( A => mult_28_C94_n208, Z => 
                           mult_28_C94_n206);
   mult_28_C94_U881 : INVDL port map( A => mult_28_C94_n207, Z => 
                           mult_28_C94_n205);
   mult_28_C94_U880 : NAN2DL port map( A1 => mult_28_C94_n386, A2 => 
                           mult_28_C94_n397, Z => mult_28_C94_n187);
   mult_28_C94_U879 : INVDL port map( A => mult_28_C94_n230, Z => 
                           mult_28_C94_n229);
   mult_28_C94_U878 : NAN2D1 port map( A1 => mult_28_C94_n346, A2 => 
                           mult_28_C94_n353, Z => mult_28_C94_n157);
   mult_28_C94_U877 : NAN2D1 port map( A1 => mult_28_C94_n354, A2 => 
                           mult_28_C94_n363, Z => mult_28_C94_n166);
   mult_28_C94_U876 : OA21D1 port map( A1 => mult_28_C94_n100, A2 => 
                           mult_28_C94_n92, B => mult_28_C94_n93, Z => 
                           mult_28_C94_n919);
   mult_28_C94_U875 : NAN2DL port map( A1 => mult_28_C94_n364, A2 => 
                           mult_28_C94_n373, Z => mult_28_C94_n175);
   mult_28_C94_U874 : OA21M20D1 port map( A1 => mult_28_C94_n124, A2 => 
                           mult_28_C94_n110, B => mult_28_C94_n113, Z => 
                           mult_28_C94_n109);
   mult_28_C94_U873 : NAN2D1 port map( A1 => mult_28_C94_n123, A2 => 
                           mult_28_C94_n101, Z => mult_28_C94_n99);
   mult_28_C94_U872 : NAN2D1 port map( A1 => mult_28_C94_n123, A2 => 
                           mult_28_C94_n110, Z => mult_28_C94_n108);
   mult_28_C94_U871 : NOR2D1 port map( A1 => mult_28_C94_n132, A2 => 
                           mult_28_C94_n125, Z => mult_28_C94_n123);
   mult_28_C94_U870 : INVDL port map( A => mult_28_C94_n165, Z => 
                           mult_28_C94_n163);
   mult_28_C94_U869 : INVDL port map( A => mult_28_C94_n193, Z => 
                           mult_28_C94_n192);
   mult_28_C94_U868 : INVD1 port map( A => mult_28_C94_n192, Z => 
                           mult_28_C94_n191);
   mult_28_C94_U867 : NOR2DL port map( A1 => mult_28_C94_n911, A2 => 
                           mult_28_C94_n920, Z => mult_28_C94_n86);
   mult_28_C94_U866 : INVD1 port map( A => mult_28_C94_n146, Z => 
                           mult_28_C94_n144);
   mult_28_C94_U865 : INVDL port map( A => mult_28_C94_n201, Z => 
                           mult_28_C94_n199);
   mult_28_C94_U864 : INVD1 port map( A => mult_28_C94_n157, Z => 
                           mult_28_C94_n155);
   mult_28_C94_U863 : NOR2D1 port map( A1 => mult_28_C94_n179, A2 => 
                           mult_28_C94_n174, Z => mult_28_C94_n172);
   mult_28_C94_U862 : NOR2D1 port map( A1 => mult_28_C94_n374, A2 => 
                           mult_28_C94_n385, Z => mult_28_C94_n179);
   mult_28_C94_U861 : NOR2D1 port map( A1 => mult_28_C94_n141, A2 => 
                           mult_28_C94_n165, Z => mult_28_C94_n139);
   mult_28_C94_U860 : INVD1 port map( A => mult_28_C94_n210, Z => 
                           mult_28_C94_n209);
   mult_28_C94_U859 : NAN2DL port map( A1 => mult_28_C94_n200, A2 => 
                           mult_28_C94_n184, Z => mult_28_C94_n182);
   mult_28_C94_U858 : BUFD4 port map( A => mult_28_C94_n181, Z => 
                           mult_28_C94_n51);
   mult_28_C94_U857 : INVDL port map( A => mult_28_C94_n180, Z => 
                           mult_28_C94_n178);
   mult_28_C94_U856 : INVD1 port map( A => mult_28_C94_n123, Z => 
                           mult_28_C94_n121);
   mult_28_C94_U855 : INVD1 port map( A => mult_28_C94_n163, Z => 
                           mult_28_C94_n161);
   mult_28_C94_U854 : INVD1 port map( A => mult_28_C94_n156, Z => 
                           mult_28_C94_n152);
   mult_28_C94_U853 : NAN2D1 port map( A1 => mult_28_C94_n163, A2 => 
                           mult_28_C94_n152, Z => mult_28_C94_n150);
   mult_28_C94_U852 : INVD1 port map( A => mult_28_C94_n164, Z => 
                           mult_28_C94_n162);
   mult_28_C94_U851 : NOR2DL port map( A1 => mult_28_C94_n911, A2 => 
                           mult_28_C94_n108, Z => mult_28_C94_n106);
   mult_28_C94_U850 : NOR2D1 port map( A1 => mult_28_C94_n911, A2 => 
                           mult_28_C94_n132, Z => mult_28_C94_n128);
   mult_28_C94_U849 : NAN2D1 port map( A1 => mult_28_C94_n154, A2 => 
                           mult_28_C94_n143, Z => mult_28_C94_n141);
   mult_28_C94_U848 : INVD1 port map( A => mult_28_C94_n913, Z => 
                           mult_28_C94_n136);
   mult_28_C94_U847 : AO21M20D1 port map( A1 => mult_28_C94_n913, A2 => 
                           mult_28_C94_n121, B => mult_28_C94_n124, Z => 
                           mult_28_C94_n116);
   mult_28_C94_U846 : NOR2D1 port map( A1 => mult_28_C94_n911, A2 => 
                           mult_28_C94_n99, Z => mult_28_C94_n95);
   mult_28_C94_U845 : INVD1 port map( A => mult_28_C94_n170, Z => 
                           mult_28_C94_n168);
   mult_28_C94_U844 : NOR2D1 port map( A1 => mult_28_C94_n170, A2 => 
                           mult_28_C94_n161, Z => mult_28_C94_n159);
   mult_28_C94_U843 : NOR2D1 port map( A1 => mult_28_C94_n170, A2 => 
                           mult_28_C94_n150, Z => mult_28_C94_n148);
   mult_28_C94_U842 : INVD1 port map( A => mult_28_C94_n911, Z => 
                           mult_28_C94_n135);
   mult_28_C94_U841 : NOR2D1 port map( A1 => mult_28_C94_n911, A2 => 
                           mult_28_C94_n121, Z => mult_28_C94_n115);
   mult_28_C94_U840 : NAN2DL port map( A1 => mult_28_C94_n522, A2 => 
                           mult_28_C94_n529, Z => mult_28_C94_n276);
   mult_28_C94_U839 : NOR2D1 port map( A1 => mult_28_C94_n516, A2 => 
                           mult_28_C94_n519, Z => mult_28_C94_n267);
   mult_28_C94_U838 : OAI22DL port map( A1 => mult_28_C94_n778, A2 => 
                           mult_28_C94_n4, B1 => mult_28_C94_n6, B2 => 
                           mult_28_C94_n779, Z => mult_28_C94_n644);
   mult_28_C94_U837 : OR2DL port map( A1 => mult_28_C94_n600, A2 => 
                           mult_28_C94_n558, Z => mult_28_C94_n423);
   mult_28_C94_U836 : AND2D1 port map( A1 => mult_28_C94_n484, A2 => 
                           mult_28_C94_n491, Z => mult_28_C94_n923);
   mult_28_C94_U835 : NAN2DL port map( A1 => mult_28_C94_n921, A2 => 
                           mult_28_C94_n922, Z => mult_28_C94_n231);
   mult_28_C94_U834 : OR2D1 port map( A1 => mult_28_C94_n464, A2 => 
                           mult_28_C94_n473, Z => mult_28_C94_n918);
   mult_28_C94_U833 : AND2DL port map( A1 => mult_28_C94_n452, A2 => 
                           mult_28_C94_n463, Z => mult_28_C94_n917);
   mult_28_C94_U832 : NAN2DL port map( A1 => mult_28_C94_n338, A2 => 
                           mult_28_C94_n345, Z => mult_28_C94_n146);
   mult_28_C94_U831 : NAN2M1D1 port map( A1 => mult_28_C94_n92, A2 => 
                           mult_28_C94_n93, Z => mult_28_C94_n55);
   mult_28_C94_U830 : NAN2M1DL port map( A1 => mult_28_C94_n213, A2 => 
                           mult_28_C94_n214, Z => mult_28_C94_n69);
   mult_28_C94_U829 : NAN2M1D1 port map( A1 => mult_28_C94_n103, A2 => 
                           mult_28_C94_n104, Z => mult_28_C94_n56);
   mult_28_C94_U828 : NAN2M1D1 port map( A1 => mult_28_C94_n112, A2 => 
                           mult_28_C94_n113, Z => mult_28_C94_n57);
   mult_28_C94_U827 : NAN2M1DL port map( A1 => mult_28_C94_n207, A2 => 
                           mult_28_C94_n208, Z => mult_28_C94_n68);
   mult_28_C94_U826 : NAN2D1 port map( A1 => mult_28_C94_n398, A2 => 
                           mult_28_C94_n411, Z => mult_28_C94_n194);
   mult_28_C94_U825 : OAI21D1 port map( A1 => mult_28_C94_n217, A2 => 
                           mult_28_C94_n213, B => mult_28_C94_n214, Z => 
                           mult_28_C94_n916);
   mult_28_C94_U824 : NOR2DL port map( A1 => mult_28_C94_n216, A2 => 
                           mult_28_C94_n213, Z => mult_28_C94_n915);
   mult_28_C94_U823 : AOI21D1 port map( A1 => mult_28_C94_n915, A2 => 
                           mult_28_C94_n230, B => mult_28_C94_n916, Z => 
                           mult_28_C94_n210);
   mult_28_C94_U822 : INVDL port map( A => mult_28_C94_n166, Z => 
                           mult_28_C94_n164);
   mult_28_C94_U821 : INVDL port map( A => mult_28_C94_n200, Z => 
                           mult_28_C94_n198);
   mult_28_C94_U820 : OAI21DL port map( A1 => mult_28_C94_n141, A2 => 
                           mult_28_C94_n166, B => mult_28_C94_n142, Z => 
                           mult_28_C94_n914);
   mult_28_C94_U819 : AOI21D1 port map( A1 => mult_28_C94_n173, A2 => 
                           mult_28_C94_n139, B => mult_28_C94_n914, Z => 
                           mult_28_C94_n913);
   mult_28_C94_U818 : NAN2M1DL port map( A1 => mult_28_C94_n186, A2 => 
                           mult_28_C94_n187, Z => mult_28_C94_n65);
   mult_28_C94_U817 : NAN2M1DL port map( A1 => mult_28_C94_n193, A2 => 
                           mult_28_C94_n194, Z => mult_28_C94_n66);
   mult_28_C94_U816 : NAN2M1D1 port map( A1 => mult_28_C94_n125, A2 => 
                           mult_28_C94_n126, Z => mult_28_C94_n58);
   mult_28_C94_U815 : NAN2M1D1 port map( A1 => mult_28_C94_n132, A2 => 
                           mult_28_C94_n133, Z => mult_28_C94_n59);
   mult_28_C94_U814 : NAN2M1DL port map( A1 => mult_28_C94_n156, A2 => 
                           mult_28_C94_n157, Z => mult_28_C94_n61);
   mult_28_C94_U813 : NAN2M1DL port map( A1 => mult_28_C94_n165, A2 => 
                           mult_28_C94_n166, Z => mult_28_C94_n62);
   mult_28_C94_U812 : NAN2DL port map( A1 => mult_28_C94_n294, A2 => 
                           mult_28_C94_n175, Z => mult_28_C94_n912);
   mult_28_C94_U811 : NAN2M1DL port map( A1 => mult_28_C94_n202, A2 => 
                           mult_28_C94_n203, Z => mult_28_C94_n67);
   mult_28_C94_U810 : INVDL port map( A => mult_28_C94_n179, Z => 
                           mult_28_C94_n177);
   mult_28_C94_U809 : NOR2DL port map( A1 => mult_28_C94_n198, A2 => 
                           mult_28_C94_n191, Z => mult_28_C94_n189);
   mult_28_C94_U808 : INVDL port map( A => mult_28_C94_n199, Z => 
                           mult_28_C94_n197);
   mult_28_C94_U807 : NAN2M1DL port map( A1 => mult_28_C94_n179, A2 => 
                           mult_28_C94_n180, Z => mult_28_C94_n64);
   mult_28_C94_U806 : AND2DL port map( A1 => mult_28_C94_n512, A2 => 
                           mult_28_C94_n515, Z => mult_28_C94_n934);
   mult_28_C94_U805 : INVDL port map( A => mult_28_C94_n409, Z => 
                           mult_28_C94_n410);
   mult_28_C94_U804 : NAN2DL port map( A1 => mult_28_C94_n440, A2 => 
                           mult_28_C94_n451, Z => mult_28_C94_n214);
   mult_28_C94_U803 : AOI21DL port map( A1 => mult_28_C94_n51, A2 => 
                           mult_28_C94_n95, B => mult_28_C94_n96, Z => 
                           mult_28_C94_n94);
   mult_28_C94_U802 : OAI21DL port map( A1 => mult_28_C94_n229, A2 => 
                           mult_28_C94_n216, B => mult_28_C94_n217, Z => 
                           mult_28_C94_n215);
   mult_28_C94_U801 : AOI21DL port map( A1 => mult_28_C94_n51, A2 => 
                           mult_28_C94_n106, B => mult_28_C94_n107, Z => 
                           mult_28_C94_n105);
   mult_28_C94_U800 : AOI21DL port map( A1 => mult_28_C94_n51, A2 => 
                           mult_28_C94_n115, B => mult_28_C94_n116, Z => 
                           mult_28_C94_n114);
   mult_28_C94_U799 : NAN2DL port map( A1 => mult_28_C94_n412, A2 => 
                           mult_28_C94_n425, Z => mult_28_C94_n203);
   mult_28_C94_U798 : INVD2 port map( A => mult_28_C94_n145, Z => 
                           mult_28_C94_n143);
   mult_28_C94_U797 : AOI21DL port map( A1 => mult_28_C94_n189, A2 => 
                           mult_28_C94_n209, B => mult_28_C94_n190, Z => 
                           mult_28_C94_n188);
   mult_28_C94_U796 : AOI21DL port map( A1 => mult_28_C94_n209, A2 => 
                           mult_28_C94_n200, B => mult_28_C94_n197, Z => 
                           mult_28_C94_n195);
   mult_28_C94_U795 : AOI21DL port map( A1 => mult_28_C94_n51, A2 => 
                           mult_28_C94_n135, B => mult_28_C94_n136, Z => 
                           mult_28_C94_n134);
   mult_28_C94_U794 : AOI21DL port map( A1 => mult_28_C94_n51, A2 => 
                           mult_28_C94_n128, B => mult_28_C94_n129, Z => 
                           mult_28_C94_n127);
   mult_28_C94_U793 : AOI21DL port map( A1 => mult_28_C94_n51, A2 => 
                           mult_28_C94_n148, B => mult_28_C94_n149, Z => 
                           mult_28_C94_n147);
   mult_28_C94_U792 : NAN2M1DL port map( A1 => mult_28_C94_n145, A2 => 
                           mult_28_C94_n146, Z => mult_28_C94_n60);
   mult_28_C94_U791 : NAN2D1 port map( A1 => mult_28_C94_n172, A2 => 
                           mult_28_C94_n139, Z => mult_28_C94_n911);
   mult_28_C94_U790 : AOI21D1 port map( A1 => mult_28_C94_n51, A2 => 
                           mult_28_C94_n159, B => mult_28_C94_n160, Z => 
                           mult_28_C94_n158);
   mult_28_C94_U789 : INVD1 port map( A => mult_28_C94_n172, Z => 
                           mult_28_C94_n170);
   mult_28_C94_U788 : EXOR2D1 port map( A1 => mult_28_C94_n176, A2 => 
                           mult_28_C94_n912, Z => m4_6);
   mult_28_C94_U787 : BUFD20 port map( A => data_in(9), Z => mult_28_C94_n801);
   mult_28_C94_U786 : BUFD20 port map( A => data_in(5), Z => mult_28_C94_n805);
   mult_28_C94_U785 : NOR2D1 port map( A1 => mult_28_C94_n332, A2 => 
                           mult_28_C94_n337, Z => mult_28_C94_n132);
   mult_28_C94_U784 : INVD1 port map( A => mult_28_C94_n173, Z => 
                           mult_28_C94_n171);
   mult_28_C94_U783 : NOR2D1 port map( A1 => mult_28_C94_n202, A2 => 
                           mult_28_C94_n207, Z => mult_28_C94_n200);
   mult_28_C94_U782 : NOR2D1 port map( A1 => mult_28_C94_n346, A2 => 
                           mult_28_C94_n353, Z => mult_28_C94_n156);
   mult_28_C94_U781 : INVDL port map( A => mult_28_C94_n156, Z => 
                           mult_28_C94_n154);
   mult_28_C94_U780 : AND2D1 port map( A1 => mult_28_C94_n464, A2 => 
                           mult_28_C94_n473, Z => mult_28_C94_n910);
   mult_28_C94_U779 : INVDL port map( A => mult_28_C94_n174, Z => 
                           mult_28_C94_n294);
   mult_28_C94_U778 : NOR2D1 port map( A1 => mult_28_C94_n193, A2 => 
                           mult_28_C94_n186, Z => mult_28_C94_n184);
   mult_28_C94_U777 : BUFD20 port map( A => data_in(10), Z => mult_28_C94_n800)
                           ;
   mult_28_C94_U773 : EXOR2D1 port map( A1 => coeff_memory_32_port, A2 => 
                           coeff_memory_33_port, Z => mult_28_C94_n818);
   mult_28_C94_U771 : EXNOR2D1 port map( A1 => coeff_memory_34_port, A2 => 
                           coeff_memory_33_port, Z => mult_28_C94_n833);
   mult_28_C94_U770 : EXOR2D1 port map( A1 => coeff_memory_34_port, A2 => 
                           coeff_memory_35_port, Z => mult_28_C94_n817);
   mult_28_C94_U768 : EXNOR2D1 port map( A1 => coeff_memory_36_port, A2 => 
                           coeff_memory_35_port, Z => mult_28_C94_n832);
   mult_28_C94_U767 : EXOR2D1 port map( A1 => coeff_memory_36_port, A2 => 
                           coeff_memory_37_port, Z => mult_28_C94_n816);
   mult_28_C94_U765 : EXNOR2D1 port map( A1 => coeff_memory_38_port, A2 => 
                           coeff_memory_37_port, Z => mult_28_C94_n831);
   mult_28_C94_U764 : EXOR2D1 port map( A1 => coeff_memory_38_port, A2 => 
                           coeff_memory_39_port, Z => mult_28_C94_n815);
   mult_28_C94_U762 : EXNOR2D1 port map( A1 => coeff_memory_40_port, A2 => 
                           coeff_memory_39_port, Z => mult_28_C94_n830);
   mult_28_C94_U761 : EXOR2D1 port map( A1 => coeff_memory_40_port, A2 => 
                           coeff_memory_41_port, Z => mult_28_C94_n814);
   mult_28_C94_U759 : EXNOR2D1 port map( A1 => coeff_memory_42_port, A2 => 
                           coeff_memory_41_port, Z => mult_28_C94_n829);
   mult_28_C94_U758 : EXOR2D1 port map( A1 => coeff_memory_42_port, A2 => 
                           coeff_memory_43_port, Z => mult_28_C94_n813);
   mult_28_C94_U756 : EXNOR2D1 port map( A1 => coeff_memory_44_port, A2 => 
                           coeff_memory_43_port, Z => mult_28_C94_n828);
   mult_28_C94_U755 : EXOR2D1 port map( A1 => coeff_memory_44_port, A2 => 
                           coeff_memory_45_port, Z => mult_28_C94_n812);
   mult_28_C94_U753 : EXNOR2D1 port map( A1 => coeff_memory_46_port, A2 => 
                           coeff_memory_45_port, Z => mult_28_C94_n827);
   mult_28_C94_U752 : EXOR2D1 port map( A1 => coeff_memory_46_port, A2 => 
                           coeff_memory_47_port, Z => mult_28_C94_n811);
   mult_28_C94_U727 : NAN2M1D1 port map( A1 => data_in(0), A2 => mult_28_C94_n1
                           , Z => mult_28_C94_n794);
   mult_28_C94_U726 : EXNOR2D1 port map( A1 => mult_28_C94_n1, A2 => data_in(0)
                           , Z => mult_28_C94_n793);
   mult_28_C94_U725 : EXNOR2D1 port map( A1 => mult_28_C94_n1, A2 => 
                           mult_28_C94_n809, Z => mult_28_C94_n792);
   mult_28_C94_U724 : EXNOR2D1 port map( A1 => mult_28_C94_n1, A2 => 
                           mult_28_C94_n808, Z => mult_28_C94_n791);
   mult_28_C94_U723 : EXNOR2D1 port map( A1 => mult_28_C94_n1, A2 => 
                           mult_28_C94_n807, Z => mult_28_C94_n790);
   mult_28_C94_U722 : EXNOR2D1 port map( A1 => mult_28_C94_n1, A2 => 
                           mult_28_C94_n806, Z => mult_28_C94_n789);
   mult_28_C94_U721 : EXNOR2D1 port map( A1 => mult_28_C94_n1, A2 => 
                           mult_28_C94_n805, Z => mult_28_C94_n788);
   mult_28_C94_U720 : EXNOR2D1 port map( A1 => mult_28_C94_n1, A2 => data_in(6)
                           , Z => mult_28_C94_n787);
   mult_28_C94_U719 : EXNOR2D1 port map( A1 => mult_28_C94_n1, A2 => 
                           mult_28_C94_n803, Z => mult_28_C94_n786);
   mult_28_C94_U718 : EXNOR2D1 port map( A1 => mult_28_C94_n1, A2 => 
                           mult_28_C94_n802, Z => mult_28_C94_n785);
   mult_28_C94_U717 : EXNOR2D1 port map( A1 => mult_28_C94_n1, A2 => 
                           mult_28_C94_n801, Z => mult_28_C94_n784);
   mult_28_C94_U716 : EXNOR2D1 port map( A1 => mult_28_C94_n1, A2 => 
                           mult_28_C94_n800, Z => mult_28_C94_n783);
   mult_28_C94_U715 : EXNOR2D1 port map( A1 => mult_28_C94_n1, A2 => 
                           mult_28_C94_n799, Z => mult_28_C94_n782);
   mult_28_C94_U714 : EXNOR2D1 port map( A1 => mult_28_C94_n1, A2 => 
                           mult_28_C94_n798, Z => mult_28_C94_n781);
   mult_28_C94_U713 : EXNOR2D1 port map( A1 => mult_28_C94_n1, A2 => 
                           mult_28_C94_n797, Z => mult_28_C94_n780);
   mult_28_C94_U712 : EXNOR2D1 port map( A1 => mult_28_C94_n1, A2 => 
                           mult_28_C94_n796, Z => mult_28_C94_n779);
   mult_28_C94_U711 : EXNOR2D1 port map( A1 => mult_28_C94_n1, A2 => 
                           mult_28_C94_n795, Z => mult_28_C94_n778);
   mult_28_C94_U709 : OAI22D1 port map( A1 => mult_28_C94_n792, A2 => 
                           mult_28_C94_n3, B1 => mult_28_C94_n5, B2 => 
                           mult_28_C94_n793, Z => mult_28_C94_n658);
   mult_28_C94_U708 : OAI22D1 port map( A1 => mult_28_C94_n791, A2 => 
                           mult_28_C94_n3, B1 => mult_28_C94_n5, B2 => 
                           mult_28_C94_n792, Z => mult_28_C94_n657);
   mult_28_C94_U707 : OAI22D1 port map( A1 => mult_28_C94_n790, A2 => 
                           mult_28_C94_n3, B1 => mult_28_C94_n5, B2 => 
                           mult_28_C94_n791, Z => mult_28_C94_n656);
   mult_28_C94_U706 : OAI22D1 port map( A1 => mult_28_C94_n789, A2 => 
                           mult_28_C94_n3, B1 => mult_28_C94_n5, B2 => 
                           mult_28_C94_n790, Z => mult_28_C94_n655);
   mult_28_C94_U705 : OAI22D1 port map( A1 => mult_28_C94_n788, A2 => 
                           mult_28_C94_n3, B1 => mult_28_C94_n5, B2 => 
                           mult_28_C94_n789, Z => mult_28_C94_n654);
   mult_28_C94_U704 : OAI22D1 port map( A1 => mult_28_C94_n787, A2 => 
                           mult_28_C94_n3, B1 => mult_28_C94_n5, B2 => 
                           mult_28_C94_n788, Z => mult_28_C94_n653);
   mult_28_C94_U703 : OAI22D1 port map( A1 => mult_28_C94_n786, A2 => 
                           mult_28_C94_n3, B1 => mult_28_C94_n5, B2 => 
                           mult_28_C94_n787, Z => mult_28_C94_n652);
   mult_28_C94_U702 : OAI22D1 port map( A1 => mult_28_C94_n785, A2 => 
                           mult_28_C94_n3, B1 => mult_28_C94_n5, B2 => 
                           mult_28_C94_n786, Z => mult_28_C94_n651);
   mult_28_C94_U701 : OAI22D1 port map( A1 => mult_28_C94_n784, A2 => 
                           mult_28_C94_n4, B1 => mult_28_C94_n6, B2 => 
                           mult_28_C94_n785, Z => mult_28_C94_n650);
   mult_28_C94_U700 : OAI22D1 port map( A1 => mult_28_C94_n783, A2 => 
                           mult_28_C94_n4, B1 => mult_28_C94_n6, B2 => 
                           mult_28_C94_n784, Z => mult_28_C94_n649);
   mult_28_C94_U699 : OAI22D1 port map( A1 => mult_28_C94_n782, A2 => 
                           mult_28_C94_n4, B1 => mult_28_C94_n6, B2 => 
                           mult_28_C94_n783, Z => mult_28_C94_n648);
   mult_28_C94_U698 : OAI22D1 port map( A1 => mult_28_C94_n781, A2 => 
                           mult_28_C94_n4, B1 => mult_28_C94_n6, B2 => 
                           mult_28_C94_n782, Z => mult_28_C94_n647);
   mult_28_C94_U697 : OAI22D1 port map( A1 => mult_28_C94_n780, A2 => 
                           mult_28_C94_n4, B1 => mult_28_C94_n6, B2 => 
                           mult_28_C94_n781, Z => mult_28_C94_n646);
   mult_28_C94_U696 : OAI22D1 port map( A1 => mult_28_C94_n779, A2 => 
                           mult_28_C94_n4, B1 => mult_28_C94_n6, B2 => 
                           mult_28_C94_n780, Z => mult_28_C94_n645);
   mult_28_C94_U693 : OAI22D1 port map( A1 => mult_28_C94_n794, A2 => 
                           mult_28_C94_n4, B1 => mult_28_C94_n6, B2 => 
                           mult_28_C94_n842, Z => mult_28_C94_n530);
   mult_28_C94_U692 : NAN2M1D1 port map( A1 => data_in(0), A2 => mult_28_C94_n7
                           , Z => mult_28_C94_n777);
   mult_28_C94_U691 : EXNOR2D1 port map( A1 => mult_28_C94_n7, A2 => data_in(0)
                           , Z => mult_28_C94_n776);
   mult_28_C94_U690 : EXNOR2D1 port map( A1 => mult_28_C94_n7, A2 => 
                           mult_28_C94_n809, Z => mult_28_C94_n775);
   mult_28_C94_U689 : EXNOR2D1 port map( A1 => mult_28_C94_n7, A2 => 
                           mult_28_C94_n808, Z => mult_28_C94_n774);
   mult_28_C94_U688 : EXNOR2D1 port map( A1 => mult_28_C94_n7, A2 => 
                           mult_28_C94_n807, Z => mult_28_C94_n773);
   mult_28_C94_U687 : EXNOR2D1 port map( A1 => mult_28_C94_n7, A2 => 
                           mult_28_C94_n806, Z => mult_28_C94_n772);
   mult_28_C94_U686 : EXNOR2D1 port map( A1 => mult_28_C94_n7, A2 => 
                           mult_28_C94_n805, Z => mult_28_C94_n771);
   mult_28_C94_U685 : EXNOR2D1 port map( A1 => mult_28_C94_n7, A2 => data_in(6)
                           , Z => mult_28_C94_n770);
   mult_28_C94_U684 : EXNOR2D1 port map( A1 => mult_28_C94_n7, A2 => 
                           mult_28_C94_n803, Z => mult_28_C94_n769);
   mult_28_C94_U683 : EXNOR2D1 port map( A1 => mult_28_C94_n7, A2 => 
                           mult_28_C94_n802, Z => mult_28_C94_n768);
   mult_28_C94_U682 : EXNOR2D1 port map( A1 => mult_28_C94_n7, A2 => 
                           mult_28_C94_n801, Z => mult_28_C94_n767);
   mult_28_C94_U681 : EXNOR2D1 port map( A1 => mult_28_C94_n7, A2 => 
                           mult_28_C94_n800, Z => mult_28_C94_n766);
   mult_28_C94_U680 : EXNOR2D1 port map( A1 => mult_28_C94_n7, A2 => 
                           mult_28_C94_n799, Z => mult_28_C94_n765);
   mult_28_C94_U679 : EXNOR2D1 port map( A1 => mult_28_C94_n7, A2 => 
                           mult_28_C94_n798, Z => mult_28_C94_n764);
   mult_28_C94_U678 : EXNOR2D1 port map( A1 => mult_28_C94_n7, A2 => 
                           mult_28_C94_n797, Z => mult_28_C94_n763);
   mult_28_C94_U677 : EXNOR2D1 port map( A1 => mult_28_C94_n7, A2 => 
                           mult_28_C94_n796, Z => mult_28_C94_n762);
   mult_28_C94_U676 : EXNOR2D1 port map( A1 => mult_28_C94_n7, A2 => 
                           mult_28_C94_n795, Z => mult_28_C94_n761);
   mult_28_C94_U675 : NOR2M1D1 port map( A1 => data_in(0), A2 => mult_28_C94_n9
                           , Z => mult_28_C94_n642);
   mult_28_C94_U674 : OAI22D1 port map( A1 => mult_28_C94_n9, A2 => 
                           mult_28_C94_n775, B1 => mult_28_C94_n11, B2 => 
                           mult_28_C94_n776, Z => mult_28_C94_n641);
   mult_28_C94_U673 : OAI22D1 port map( A1 => mult_28_C94_n9, A2 => 
                           mult_28_C94_n774, B1 => mult_28_C94_n11, B2 => 
                           mult_28_C94_n775, Z => mult_28_C94_n640);
   mult_28_C94_U672 : OAI22D1 port map( A1 => mult_28_C94_n9, A2 => 
                           mult_28_C94_n773, B1 => mult_28_C94_n11, B2 => 
                           mult_28_C94_n774, Z => mult_28_C94_n639);
   mult_28_C94_U671 : OAI22D1 port map( A1 => mult_28_C94_n9, A2 => 
                           mult_28_C94_n772, B1 => mult_28_C94_n11, B2 => 
                           mult_28_C94_n773, Z => mult_28_C94_n638);
   mult_28_C94_U670 : OAI22D1 port map( A1 => mult_28_C94_n9, A2 => 
                           mult_28_C94_n771, B1 => mult_28_C94_n11, B2 => 
                           mult_28_C94_n772, Z => mult_28_C94_n637);
   mult_28_C94_U669 : OAI22D1 port map( A1 => mult_28_C94_n9, A2 => 
                           mult_28_C94_n770, B1 => mult_28_C94_n11, B2 => 
                           mult_28_C94_n771, Z => mult_28_C94_n636);
   mult_28_C94_U668 : OAI22D1 port map( A1 => mult_28_C94_n9, A2 => 
                           mult_28_C94_n769, B1 => mult_28_C94_n11, B2 => 
                           mult_28_C94_n770, Z => mult_28_C94_n635);
   mult_28_C94_U667 : OAI22D1 port map( A1 => mult_28_C94_n9, A2 => 
                           mult_28_C94_n768, B1 => mult_28_C94_n11, B2 => 
                           mult_28_C94_n769, Z => mult_28_C94_n634);
   mult_28_C94_U666 : OAI22D1 port map( A1 => mult_28_C94_n10, A2 => 
                           mult_28_C94_n767, B1 => mult_28_C94_n12, B2 => 
                           mult_28_C94_n768, Z => mult_28_C94_n633);
   mult_28_C94_U665 : OAI22D1 port map( A1 => mult_28_C94_n10, A2 => 
                           mult_28_C94_n766, B1 => mult_28_C94_n12, B2 => 
                           mult_28_C94_n767, Z => mult_28_C94_n632);
   mult_28_C94_U664 : OAI22D1 port map( A1 => mult_28_C94_n10, A2 => 
                           mult_28_C94_n765, B1 => mult_28_C94_n12, B2 => 
                           mult_28_C94_n766, Z => mult_28_C94_n631);
   mult_28_C94_U663 : OAI22D1 port map( A1 => mult_28_C94_n10, A2 => 
                           mult_28_C94_n764, B1 => mult_28_C94_n12, B2 => 
                           mult_28_C94_n765, Z => mult_28_C94_n630);
   mult_28_C94_U662 : OAI22D1 port map( A1 => mult_28_C94_n10, A2 => 
                           mult_28_C94_n763, B1 => mult_28_C94_n12, B2 => 
                           mult_28_C94_n764, Z => mult_28_C94_n629);
   mult_28_C94_U661 : OAI22D1 port map( A1 => mult_28_C94_n10, A2 => 
                           mult_28_C94_n762, B1 => mult_28_C94_n12, B2 => 
                           mult_28_C94_n763, Z => mult_28_C94_n628);
   mult_28_C94_U660 : OAI22D1 port map( A1 => mult_28_C94_n10, A2 => 
                           mult_28_C94_n761, B1 => mult_28_C94_n12, B2 => 
                           mult_28_C94_n762, Z => mult_28_C94_n409);
   mult_28_C94_U657 : NAN2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C94_n13, Z => mult_28_C94_n760);
   mult_28_C94_U656 : EXNOR2D1 port map( A1 => mult_28_C94_n13, A2 => 
                           data_in(0), Z => mult_28_C94_n759);
   mult_28_C94_U655 : EXNOR2D1 port map( A1 => mult_28_C94_n13, A2 => 
                           mult_28_C94_n809, Z => mult_28_C94_n758);
   mult_28_C94_U654 : EXNOR2D1 port map( A1 => mult_28_C94_n13, A2 => 
                           mult_28_C94_n808, Z => mult_28_C94_n757);
   mult_28_C94_U653 : EXNOR2D1 port map( A1 => mult_28_C94_n13, A2 => 
                           mult_28_C94_n807, Z => mult_28_C94_n756);
   mult_28_C94_U652 : EXNOR2D1 port map( A1 => mult_28_C94_n13, A2 => 
                           mult_28_C94_n806, Z => mult_28_C94_n755);
   mult_28_C94_U651 : EXNOR2D1 port map( A1 => mult_28_C94_n13, A2 => 
                           mult_28_C94_n805, Z => mult_28_C94_n754);
   mult_28_C94_U650 : EXNOR2D1 port map( A1 => mult_28_C94_n13, A2 => 
                           data_in(6), Z => mult_28_C94_n753);
   mult_28_C94_U649 : EXNOR2D1 port map( A1 => mult_28_C94_n13, A2 => 
                           mult_28_C94_n803, Z => mult_28_C94_n752);
   mult_28_C94_U648 : EXNOR2D1 port map( A1 => mult_28_C94_n13, A2 => 
                           mult_28_C94_n802, Z => mult_28_C94_n751);
   mult_28_C94_U647 : EXNOR2D1 port map( A1 => mult_28_C94_n13, A2 => 
                           mult_28_C94_n801, Z => mult_28_C94_n750);
   mult_28_C94_U646 : EXNOR2D1 port map( A1 => mult_28_C94_n13, A2 => 
                           mult_28_C94_n800, Z => mult_28_C94_n749);
   mult_28_C94_U645 : EXNOR2D1 port map( A1 => mult_28_C94_n13, A2 => 
                           mult_28_C94_n799, Z => mult_28_C94_n748);
   mult_28_C94_U644 : EXNOR2D1 port map( A1 => mult_28_C94_n13, A2 => 
                           mult_28_C94_n798, Z => mult_28_C94_n747);
   mult_28_C94_U643 : EXNOR2D1 port map( A1 => mult_28_C94_n13, A2 => 
                           mult_28_C94_n797, Z => mult_28_C94_n746);
   mult_28_C94_U642 : EXNOR2D1 port map( A1 => mult_28_C94_n13, A2 => 
                           mult_28_C94_n796, Z => mult_28_C94_n745);
   mult_28_C94_U641 : EXNOR2D1 port map( A1 => mult_28_C94_n13, A2 => 
                           mult_28_C94_n795, Z => mult_28_C94_n744);
   mult_28_C94_U640 : NOR2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C94_n15, Z => mult_28_C94_n626);
   mult_28_C94_U639 : OAI22D1 port map( A1 => mult_28_C94_n15, A2 => 
                           mult_28_C94_n758, B1 => mult_28_C94_n17, B2 => 
                           mult_28_C94_n759, Z => mult_28_C94_n625);
   mult_28_C94_U638 : OAI22D1 port map( A1 => mult_28_C94_n15, A2 => 
                           mult_28_C94_n757, B1 => mult_28_C94_n17, B2 => 
                           mult_28_C94_n758, Z => mult_28_C94_n624);
   mult_28_C94_U637 : OAI22D1 port map( A1 => mult_28_C94_n15, A2 => 
                           mult_28_C94_n756, B1 => mult_28_C94_n17, B2 => 
                           mult_28_C94_n757, Z => mult_28_C94_n623);
   mult_28_C94_U636 : OAI22D1 port map( A1 => mult_28_C94_n15, A2 => 
                           mult_28_C94_n755, B1 => mult_28_C94_n17, B2 => 
                           mult_28_C94_n756, Z => mult_28_C94_n622);
   mult_28_C94_U635 : OAI22D1 port map( A1 => mult_28_C94_n15, A2 => 
                           mult_28_C94_n754, B1 => mult_28_C94_n17, B2 => 
                           mult_28_C94_n755, Z => mult_28_C94_n621);
   mult_28_C94_U634 : OAI22D1 port map( A1 => mult_28_C94_n15, A2 => 
                           mult_28_C94_n753, B1 => mult_28_C94_n17, B2 => 
                           mult_28_C94_n754, Z => mult_28_C94_n620);
   mult_28_C94_U633 : OAI22D1 port map( A1 => mult_28_C94_n15, A2 => 
                           mult_28_C94_n752, B1 => mult_28_C94_n17, B2 => 
                           mult_28_C94_n753, Z => mult_28_C94_n619);
   mult_28_C94_U632 : OAI22D1 port map( A1 => mult_28_C94_n15, A2 => 
                           mult_28_C94_n751, B1 => mult_28_C94_n17, B2 => 
                           mult_28_C94_n752, Z => mult_28_C94_n618);
   mult_28_C94_U631 : OAI22D1 port map( A1 => mult_28_C94_n16, A2 => 
                           mult_28_C94_n750, B1 => mult_28_C94_n18, B2 => 
                           mult_28_C94_n751, Z => mult_28_C94_n617);
   mult_28_C94_U630 : OAI22D1 port map( A1 => mult_28_C94_n16, A2 => 
                           mult_28_C94_n749, B1 => mult_28_C94_n18, B2 => 
                           mult_28_C94_n750, Z => mult_28_C94_n616);
   mult_28_C94_U629 : OAI22D1 port map( A1 => mult_28_C94_n16, A2 => 
                           mult_28_C94_n748, B1 => mult_28_C94_n18, B2 => 
                           mult_28_C94_n749, Z => mult_28_C94_n615);
   mult_28_C94_U628 : OAI22D1 port map( A1 => mult_28_C94_n16, A2 => 
                           mult_28_C94_n747, B1 => mult_28_C94_n18, B2 => 
                           mult_28_C94_n748, Z => mult_28_C94_n614);
   mult_28_C94_U627 : OAI22D1 port map( A1 => mult_28_C94_n16, A2 => 
                           mult_28_C94_n746, B1 => mult_28_C94_n18, B2 => 
                           mult_28_C94_n747, Z => mult_28_C94_n613);
   mult_28_C94_U626 : OAI22D1 port map( A1 => mult_28_C94_n16, A2 => 
                           mult_28_C94_n745, B1 => mult_28_C94_n18, B2 => 
                           mult_28_C94_n746, Z => mult_28_C94_n612);
   mult_28_C94_U625 : OAI22D1 port map( A1 => mult_28_C94_n16, A2 => 
                           mult_28_C94_n744, B1 => mult_28_C94_n18, B2 => 
                           mult_28_C94_n745, Z => mult_28_C94_n383);
   mult_28_C94_U623 : OAI22D1 port map( A1 => mult_28_C94_n16, A2 => 
                           mult_28_C94_n760, B1 => mult_28_C94_n18, B2 => 
                           mult_28_C94_n840, Z => mult_28_C94_n528);
   mult_28_C94_U622 : NAN2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C94_n19, Z => mult_28_C94_n743);
   mult_28_C94_U621 : EXNOR2D1 port map( A1 => mult_28_C94_n19, A2 => 
                           data_in(0), Z => mult_28_C94_n742);
   mult_28_C94_U620 : EXNOR2D1 port map( A1 => mult_28_C94_n19, A2 => 
                           mult_28_C94_n809, Z => mult_28_C94_n741);
   mult_28_C94_U619 : EXNOR2D1 port map( A1 => mult_28_C94_n19, A2 => 
                           mult_28_C94_n808, Z => mult_28_C94_n740);
   mult_28_C94_U618 : EXNOR2D1 port map( A1 => mult_28_C94_n19, A2 => 
                           mult_28_C94_n807, Z => mult_28_C94_n739);
   mult_28_C94_U617 : EXNOR2D1 port map( A1 => mult_28_C94_n19, A2 => 
                           mult_28_C94_n806, Z => mult_28_C94_n738);
   mult_28_C94_U616 : EXNOR2D1 port map( A1 => mult_28_C94_n19, A2 => 
                           mult_28_C94_n805, Z => mult_28_C94_n737);
   mult_28_C94_U615 : EXNOR2D1 port map( A1 => mult_28_C94_n19, A2 => 
                           data_in(6), Z => mult_28_C94_n736);
   mult_28_C94_U614 : EXNOR2D1 port map( A1 => mult_28_C94_n19, A2 => 
                           mult_28_C94_n803, Z => mult_28_C94_n735);
   mult_28_C94_U613 : EXNOR2D1 port map( A1 => mult_28_C94_n19, A2 => 
                           mult_28_C94_n802, Z => mult_28_C94_n734);
   mult_28_C94_U612 : EXNOR2D1 port map( A1 => mult_28_C94_n19, A2 => 
                           mult_28_C94_n801, Z => mult_28_C94_n733);
   mult_28_C94_U611 : EXNOR2D1 port map( A1 => mult_28_C94_n19, A2 => 
                           mult_28_C94_n800, Z => mult_28_C94_n732);
   mult_28_C94_U610 : EXNOR2D1 port map( A1 => mult_28_C94_n19, A2 => 
                           mult_28_C94_n799, Z => mult_28_C94_n731);
   mult_28_C94_U609 : EXNOR2D1 port map( A1 => mult_28_C94_n19, A2 => 
                           mult_28_C94_n798, Z => mult_28_C94_n730);
   mult_28_C94_U608 : EXNOR2D1 port map( A1 => mult_28_C94_n19, A2 => 
                           mult_28_C94_n797, Z => mult_28_C94_n729);
   mult_28_C94_U607 : EXNOR2D1 port map( A1 => mult_28_C94_n19, A2 => 
                           mult_28_C94_n796, Z => mult_28_C94_n728);
   mult_28_C94_U606 : EXNOR2D1 port map( A1 => mult_28_C94_n19, A2 => 
                           mult_28_C94_n795, Z => mult_28_C94_n727);
   mult_28_C94_U605 : NOR2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C94_n21, Z => mult_28_C94_n610);
   mult_28_C94_U604 : OAI22D1 port map( A1 => mult_28_C94_n21, A2 => 
                           mult_28_C94_n741, B1 => mult_28_C94_n23, B2 => 
                           mult_28_C94_n742, Z => mult_28_C94_n609);
   mult_28_C94_U603 : OAI22D1 port map( A1 => mult_28_C94_n21, A2 => 
                           mult_28_C94_n740, B1 => mult_28_C94_n23, B2 => 
                           mult_28_C94_n741, Z => mult_28_C94_n608);
   mult_28_C94_U602 : OAI22D1 port map( A1 => mult_28_C94_n21, A2 => 
                           mult_28_C94_n739, B1 => mult_28_C94_n23, B2 => 
                           mult_28_C94_n740, Z => mult_28_C94_n607);
   mult_28_C94_U601 : OAI22D1 port map( A1 => mult_28_C94_n21, A2 => 
                           mult_28_C94_n738, B1 => mult_28_C94_n23, B2 => 
                           mult_28_C94_n739, Z => mult_28_C94_n606);
   mult_28_C94_U600 : OAI22D1 port map( A1 => mult_28_C94_n21, A2 => 
                           mult_28_C94_n737, B1 => mult_28_C94_n23, B2 => 
                           mult_28_C94_n738, Z => mult_28_C94_n605);
   mult_28_C94_U599 : OAI22D1 port map( A1 => mult_28_C94_n21, A2 => 
                           mult_28_C94_n736, B1 => mult_28_C94_n23, B2 => 
                           mult_28_C94_n737, Z => mult_28_C94_n604);
   mult_28_C94_U598 : OAI22D1 port map( A1 => mult_28_C94_n21, A2 => 
                           mult_28_C94_n735, B1 => mult_28_C94_n23, B2 => 
                           mult_28_C94_n736, Z => mult_28_C94_n603);
   mult_28_C94_U597 : OAI22D1 port map( A1 => mult_28_C94_n21, A2 => 
                           mult_28_C94_n734, B1 => mult_28_C94_n23, B2 => 
                           mult_28_C94_n735, Z => mult_28_C94_n602);
   mult_28_C94_U596 : OAI22D1 port map( A1 => mult_28_C94_n22, A2 => 
                           mult_28_C94_n733, B1 => mult_28_C94_n24, B2 => 
                           mult_28_C94_n734, Z => mult_28_C94_n601);
   mult_28_C94_U595 : OAI22D1 port map( A1 => mult_28_C94_n22, A2 => 
                           mult_28_C94_n732, B1 => mult_28_C94_n24, B2 => 
                           mult_28_C94_n733, Z => mult_28_C94_n600);
   mult_28_C94_U594 : OAI22D1 port map( A1 => mult_28_C94_n22, A2 => 
                           mult_28_C94_n731, B1 => mult_28_C94_n24, B2 => 
                           mult_28_C94_n732, Z => mult_28_C94_n599);
   mult_28_C94_U593 : OAI22D1 port map( A1 => mult_28_C94_n22, A2 => 
                           mult_28_C94_n730, B1 => mult_28_C94_n24, B2 => 
                           mult_28_C94_n731, Z => mult_28_C94_n598);
   mult_28_C94_U592 : OAI22D1 port map( A1 => mult_28_C94_n22, A2 => 
                           mult_28_C94_n729, B1 => mult_28_C94_n24, B2 => 
                           mult_28_C94_n730, Z => mult_28_C94_n597);
   mult_28_C94_U591 : OAI22D1 port map( A1 => mult_28_C94_n22, A2 => 
                           mult_28_C94_n728, B1 => mult_28_C94_n24, B2 => 
                           mult_28_C94_n729, Z => mult_28_C94_n596);
   mult_28_C94_U590 : OAI22D1 port map( A1 => mult_28_C94_n22, A2 => 
                           mult_28_C94_n727, B1 => mult_28_C94_n24, B2 => 
                           mult_28_C94_n728, Z => mult_28_C94_n361);
   mult_28_C94_U588 : OAI22D1 port map( A1 => mult_28_C94_n22, A2 => 
                           mult_28_C94_n743, B1 => mult_28_C94_n24, B2 => 
                           mult_28_C94_n839, Z => mult_28_C94_n527);
   mult_28_C94_U587 : NAN2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C94_n25, Z => mult_28_C94_n726);
   mult_28_C94_U586 : EXNOR2D1 port map( A1 => mult_28_C94_n25, A2 => 
                           data_in(0), Z => mult_28_C94_n725);
   mult_28_C94_U585 : EXNOR2D1 port map( A1 => mult_28_C94_n25, A2 => 
                           mult_28_C94_n809, Z => mult_28_C94_n724);
   mult_28_C94_U584 : EXNOR2D1 port map( A1 => mult_28_C94_n25, A2 => 
                           mult_28_C94_n808, Z => mult_28_C94_n723);
   mult_28_C94_U583 : EXNOR2D1 port map( A1 => mult_28_C94_n25, A2 => 
                           mult_28_C94_n807, Z => mult_28_C94_n722);
   mult_28_C94_U582 : EXNOR2D1 port map( A1 => mult_28_C94_n25, A2 => 
                           mult_28_C94_n806, Z => mult_28_C94_n721);
   mult_28_C94_U581 : EXNOR2D1 port map( A1 => mult_28_C94_n25, A2 => 
                           mult_28_C94_n805, Z => mult_28_C94_n720);
   mult_28_C94_U580 : EXNOR2D1 port map( A1 => mult_28_C94_n25, A2 => 
                           data_in(6), Z => mult_28_C94_n719);
   mult_28_C94_U579 : EXNOR2D1 port map( A1 => mult_28_C94_n25, A2 => 
                           mult_28_C94_n803, Z => mult_28_C94_n718);
   mult_28_C94_U578 : EXNOR2D1 port map( A1 => mult_28_C94_n25, A2 => 
                           mult_28_C94_n802, Z => mult_28_C94_n717);
   mult_28_C94_U577 : EXNOR2D1 port map( A1 => mult_28_C94_n25, A2 => 
                           mult_28_C94_n801, Z => mult_28_C94_n716);
   mult_28_C94_U576 : EXNOR2D1 port map( A1 => mult_28_C94_n25, A2 => 
                           mult_28_C94_n800, Z => mult_28_C94_n715);
   mult_28_C94_U575 : EXNOR2D1 port map( A1 => mult_28_C94_n25, A2 => 
                           mult_28_C94_n799, Z => mult_28_C94_n714);
   mult_28_C94_U574 : EXNOR2D1 port map( A1 => mult_28_C94_n25, A2 => 
                           mult_28_C94_n798, Z => mult_28_C94_n713);
   mult_28_C94_U573 : EXNOR2D1 port map( A1 => mult_28_C94_n25, A2 => 
                           mult_28_C94_n797, Z => mult_28_C94_n712);
   mult_28_C94_U572 : EXNOR2D1 port map( A1 => mult_28_C94_n25, A2 => 
                           mult_28_C94_n796, Z => mult_28_C94_n711);
   mult_28_C94_U571 : EXNOR2D1 port map( A1 => mult_28_C94_n25, A2 => 
                           mult_28_C94_n795, Z => mult_28_C94_n710);
   mult_28_C94_U570 : NOR2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C94_n27, Z => mult_28_C94_n594);
   mult_28_C94_U569 : OAI22D1 port map( A1 => mult_28_C94_n27, A2 => 
                           mult_28_C94_n724, B1 => mult_28_C94_n29, B2 => 
                           mult_28_C94_n725, Z => mult_28_C94_n593);
   mult_28_C94_U568 : OAI22D1 port map( A1 => mult_28_C94_n27, A2 => 
                           mult_28_C94_n723, B1 => mult_28_C94_n29, B2 => 
                           mult_28_C94_n724, Z => mult_28_C94_n592);
   mult_28_C94_U567 : OAI22D1 port map( A1 => mult_28_C94_n27, A2 => 
                           mult_28_C94_n722, B1 => mult_28_C94_n29, B2 => 
                           mult_28_C94_n723, Z => mult_28_C94_n591);
   mult_28_C94_U566 : OAI22D1 port map( A1 => mult_28_C94_n27, A2 => 
                           mult_28_C94_n721, B1 => mult_28_C94_n29, B2 => 
                           mult_28_C94_n722, Z => mult_28_C94_n590);
   mult_28_C94_U565 : OAI22D1 port map( A1 => mult_28_C94_n27, A2 => 
                           mult_28_C94_n720, B1 => mult_28_C94_n29, B2 => 
                           mult_28_C94_n721, Z => mult_28_C94_n589);
   mult_28_C94_U564 : OAI22D1 port map( A1 => mult_28_C94_n27, A2 => 
                           mult_28_C94_n719, B1 => mult_28_C94_n29, B2 => 
                           mult_28_C94_n720, Z => mult_28_C94_n588);
   mult_28_C94_U563 : OAI22D1 port map( A1 => mult_28_C94_n27, A2 => 
                           mult_28_C94_n718, B1 => mult_28_C94_n29, B2 => 
                           mult_28_C94_n719, Z => mult_28_C94_n587);
   mult_28_C94_U562 : OAI22D1 port map( A1 => mult_28_C94_n27, A2 => 
                           mult_28_C94_n717, B1 => mult_28_C94_n29, B2 => 
                           mult_28_C94_n718, Z => mult_28_C94_n586);
   mult_28_C94_U561 : OAI22D1 port map( A1 => mult_28_C94_n28, A2 => 
                           mult_28_C94_n716, B1 => mult_28_C94_n30, B2 => 
                           mult_28_C94_n717, Z => mult_28_C94_n585);
   mult_28_C94_U560 : OAI22D1 port map( A1 => mult_28_C94_n28, A2 => 
                           mult_28_C94_n715, B1 => mult_28_C94_n30, B2 => 
                           mult_28_C94_n716, Z => mult_28_C94_n584);
   mult_28_C94_U559 : OAI22D1 port map( A1 => mult_28_C94_n28, A2 => 
                           mult_28_C94_n714, B1 => mult_28_C94_n30, B2 => 
                           mult_28_C94_n715, Z => mult_28_C94_n583);
   mult_28_C94_U558 : OAI22D1 port map( A1 => mult_28_C94_n28, A2 => 
                           mult_28_C94_n713, B1 => mult_28_C94_n30, B2 => 
                           mult_28_C94_n714, Z => mult_28_C94_n582);
   mult_28_C94_U557 : OAI22D1 port map( A1 => mult_28_C94_n28, A2 => 
                           mult_28_C94_n712, B1 => mult_28_C94_n30, B2 => 
                           mult_28_C94_n713, Z => mult_28_C94_n581);
   mult_28_C94_U556 : OAI22D1 port map( A1 => mult_28_C94_n28, A2 => 
                           mult_28_C94_n711, B1 => mult_28_C94_n30, B2 => 
                           mult_28_C94_n712, Z => mult_28_C94_n580);
   mult_28_C94_U555 : OAI22D1 port map( A1 => mult_28_C94_n28, A2 => 
                           mult_28_C94_n710, B1 => mult_28_C94_n30, B2 => 
                           mult_28_C94_n711, Z => mult_28_C94_n343);
   mult_28_C94_U553 : OAI22D1 port map( A1 => mult_28_C94_n28, A2 => 
                           mult_28_C94_n726, B1 => mult_28_C94_n30, B2 => 
                           mult_28_C94_n838, Z => mult_28_C94_n526);
   mult_28_C94_U552 : NAN2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C94_n31, Z => mult_28_C94_n709);
   mult_28_C94_U551 : EXNOR2D1 port map( A1 => mult_28_C94_n31, A2 => 
                           data_in(0), Z => mult_28_C94_n708);
   mult_28_C94_U550 : EXNOR2D1 port map( A1 => mult_28_C94_n31, A2 => 
                           mult_28_C94_n809, Z => mult_28_C94_n707);
   mult_28_C94_U549 : EXNOR2D1 port map( A1 => mult_28_C94_n31, A2 => 
                           mult_28_C94_n808, Z => mult_28_C94_n706);
   mult_28_C94_U548 : EXNOR2D1 port map( A1 => mult_28_C94_n31, A2 => 
                           mult_28_C94_n807, Z => mult_28_C94_n705);
   mult_28_C94_U547 : EXNOR2D1 port map( A1 => mult_28_C94_n31, A2 => 
                           mult_28_C94_n806, Z => mult_28_C94_n704);
   mult_28_C94_U546 : EXNOR2D1 port map( A1 => mult_28_C94_n31, A2 => 
                           mult_28_C94_n805, Z => mult_28_C94_n703);
   mult_28_C94_U545 : EXNOR2D1 port map( A1 => mult_28_C94_n31, A2 => 
                           data_in(6), Z => mult_28_C94_n702);
   mult_28_C94_U544 : EXNOR2D1 port map( A1 => mult_28_C94_n31, A2 => 
                           mult_28_C94_n803, Z => mult_28_C94_n701);
   mult_28_C94_U543 : EXNOR2D1 port map( A1 => mult_28_C94_n31, A2 => 
                           mult_28_C94_n802, Z => mult_28_C94_n700);
   mult_28_C94_U542 : EXNOR2D1 port map( A1 => mult_28_C94_n31, A2 => 
                           mult_28_C94_n801, Z => mult_28_C94_n699);
   mult_28_C94_U541 : EXNOR2D1 port map( A1 => mult_28_C94_n31, A2 => 
                           mult_28_C94_n800, Z => mult_28_C94_n698);
   mult_28_C94_U540 : EXNOR2D1 port map( A1 => mult_28_C94_n31, A2 => 
                           mult_28_C94_n799, Z => mult_28_C94_n697);
   mult_28_C94_U539 : EXNOR2D1 port map( A1 => mult_28_C94_n31, A2 => 
                           mult_28_C94_n798, Z => mult_28_C94_n696);
   mult_28_C94_U538 : EXNOR2D1 port map( A1 => mult_28_C94_n31, A2 => 
                           mult_28_C94_n797, Z => mult_28_C94_n695);
   mult_28_C94_U537 : EXNOR2D1 port map( A1 => mult_28_C94_n31, A2 => 
                           mult_28_C94_n796, Z => mult_28_C94_n694);
   mult_28_C94_U536 : EXNOR2D1 port map( A1 => mult_28_C94_n31, A2 => 
                           mult_28_C94_n795, Z => mult_28_C94_n693);
   mult_28_C94_U535 : NOR2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C94_n33, Z => mult_28_C94_n578);
   mult_28_C94_U534 : OAI22D1 port map( A1 => mult_28_C94_n33, A2 => 
                           mult_28_C94_n707, B1 => mult_28_C94_n35, B2 => 
                           mult_28_C94_n708, Z => mult_28_C94_n577);
   mult_28_C94_U533 : OAI22D1 port map( A1 => mult_28_C94_n33, A2 => 
                           mult_28_C94_n706, B1 => mult_28_C94_n35, B2 => 
                           mult_28_C94_n707, Z => mult_28_C94_n576);
   mult_28_C94_U532 : OAI22D1 port map( A1 => mult_28_C94_n33, A2 => 
                           mult_28_C94_n705, B1 => mult_28_C94_n35, B2 => 
                           mult_28_C94_n706, Z => mult_28_C94_n575);
   mult_28_C94_U531 : OAI22D1 port map( A1 => mult_28_C94_n33, A2 => 
                           mult_28_C94_n704, B1 => mult_28_C94_n35, B2 => 
                           mult_28_C94_n705, Z => mult_28_C94_n574);
   mult_28_C94_U530 : OAI22D1 port map( A1 => mult_28_C94_n33, A2 => 
                           mult_28_C94_n703, B1 => mult_28_C94_n35, B2 => 
                           mult_28_C94_n704, Z => mult_28_C94_n573);
   mult_28_C94_U529 : OAI22D1 port map( A1 => mult_28_C94_n33, A2 => 
                           mult_28_C94_n702, B1 => mult_28_C94_n35, B2 => 
                           mult_28_C94_n703, Z => mult_28_C94_n572);
   mult_28_C94_U528 : OAI22D1 port map( A1 => mult_28_C94_n33, A2 => 
                           mult_28_C94_n701, B1 => mult_28_C94_n35, B2 => 
                           mult_28_C94_n702, Z => mult_28_C94_n571);
   mult_28_C94_U527 : OAI22D1 port map( A1 => mult_28_C94_n33, A2 => 
                           mult_28_C94_n700, B1 => mult_28_C94_n35, B2 => 
                           mult_28_C94_n701, Z => mult_28_C94_n570);
   mult_28_C94_U526 : OAI22D1 port map( A1 => mult_28_C94_n34, A2 => 
                           mult_28_C94_n699, B1 => mult_28_C94_n36, B2 => 
                           mult_28_C94_n700, Z => mult_28_C94_n569);
   mult_28_C94_U525 : OAI22D1 port map( A1 => mult_28_C94_n34, A2 => 
                           mult_28_C94_n698, B1 => mult_28_C94_n36, B2 => 
                           mult_28_C94_n699, Z => mult_28_C94_n568);
   mult_28_C94_U524 : OAI22D1 port map( A1 => mult_28_C94_n34, A2 => 
                           mult_28_C94_n697, B1 => mult_28_C94_n36, B2 => 
                           mult_28_C94_n698, Z => mult_28_C94_n567);
   mult_28_C94_U523 : OAI22D1 port map( A1 => mult_28_C94_n34, A2 => 
                           mult_28_C94_n696, B1 => mult_28_C94_n36, B2 => 
                           mult_28_C94_n697, Z => mult_28_C94_n566);
   mult_28_C94_U522 : OAI22D1 port map( A1 => mult_28_C94_n34, A2 => 
                           mult_28_C94_n695, B1 => mult_28_C94_n36, B2 => 
                           mult_28_C94_n696, Z => mult_28_C94_n565);
   mult_28_C94_U521 : OAI22D1 port map( A1 => mult_28_C94_n34, A2 => 
                           mult_28_C94_n694, B1 => mult_28_C94_n36, B2 => 
                           mult_28_C94_n695, Z => mult_28_C94_n564);
   mult_28_C94_U520 : OAI22D1 port map( A1 => mult_28_C94_n34, A2 => 
                           mult_28_C94_n693, B1 => mult_28_C94_n36, B2 => 
                           mult_28_C94_n694, Z => mult_28_C94_n329);
   mult_28_C94_U518 : OAI22D1 port map( A1 => mult_28_C94_n34, A2 => 
                           mult_28_C94_n709, B1 => mult_28_C94_n36, B2 => 
                           mult_28_C94_n837, Z => mult_28_C94_n525);
   mult_28_C94_U517 : NAN2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C94_n37, Z => mult_28_C94_n692);
   mult_28_C94_U516 : EXNOR2D1 port map( A1 => mult_28_C94_n37, A2 => 
                           data_in(0), Z => mult_28_C94_n691);
   mult_28_C94_U515 : EXNOR2D1 port map( A1 => mult_28_C94_n37, A2 => 
                           mult_28_C94_n809, Z => mult_28_C94_n690);
   mult_28_C94_U514 : EXNOR2D1 port map( A1 => mult_28_C94_n37, A2 => 
                           mult_28_C94_n808, Z => mult_28_C94_n689);
   mult_28_C94_U513 : EXNOR2D1 port map( A1 => mult_28_C94_n37, A2 => 
                           mult_28_C94_n807, Z => mult_28_C94_n688);
   mult_28_C94_U512 : EXNOR2D1 port map( A1 => mult_28_C94_n37, A2 => 
                           mult_28_C94_n806, Z => mult_28_C94_n687);
   mult_28_C94_U511 : EXNOR2D1 port map( A1 => mult_28_C94_n37, A2 => 
                           mult_28_C94_n805, Z => mult_28_C94_n686);
   mult_28_C94_U510 : EXNOR2D1 port map( A1 => mult_28_C94_n37, A2 => 
                           data_in(6), Z => mult_28_C94_n685);
   mult_28_C94_U509 : EXNOR2D1 port map( A1 => mult_28_C94_n37, A2 => 
                           mult_28_C94_n803, Z => mult_28_C94_n684);
   mult_28_C94_U508 : EXNOR2D1 port map( A1 => mult_28_C94_n37, A2 => 
                           mult_28_C94_n802, Z => mult_28_C94_n683);
   mult_28_C94_U507 : EXNOR2D1 port map( A1 => mult_28_C94_n37, A2 => 
                           mult_28_C94_n801, Z => mult_28_C94_n682);
   mult_28_C94_U506 : EXNOR2D1 port map( A1 => mult_28_C94_n37, A2 => 
                           mult_28_C94_n800, Z => mult_28_C94_n681);
   mult_28_C94_U505 : EXNOR2D1 port map( A1 => mult_28_C94_n37, A2 => 
                           mult_28_C94_n799, Z => mult_28_C94_n680);
   mult_28_C94_U504 : EXNOR2D1 port map( A1 => mult_28_C94_n37, A2 => 
                           mult_28_C94_n798, Z => mult_28_C94_n679);
   mult_28_C94_U503 : EXNOR2D1 port map( A1 => mult_28_C94_n37, A2 => 
                           mult_28_C94_n797, Z => mult_28_C94_n678);
   mult_28_C94_U502 : EXNOR2D1 port map( A1 => mult_28_C94_n37, A2 => 
                           mult_28_C94_n796, Z => mult_28_C94_n677);
   mult_28_C94_U501 : EXNOR2D1 port map( A1 => mult_28_C94_n37, A2 => 
                           mult_28_C94_n795, Z => mult_28_C94_n676);
   mult_28_C94_U500 : NOR2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C94_n39, Z => mult_28_C94_n562);
   mult_28_C94_U499 : OAI22D1 port map( A1 => mult_28_C94_n39, A2 => 
                           mult_28_C94_n690, B1 => mult_28_C94_n41, B2 => 
                           mult_28_C94_n691, Z => mult_28_C94_n561);
   mult_28_C94_U498 : OAI22D1 port map( A1 => mult_28_C94_n39, A2 => 
                           mult_28_C94_n689, B1 => mult_28_C94_n41, B2 => 
                           mult_28_C94_n690, Z => mult_28_C94_n560);
   mult_28_C94_U497 : OAI22D1 port map( A1 => mult_28_C94_n39, A2 => 
                           mult_28_C94_n688, B1 => mult_28_C94_n41, B2 => 
                           mult_28_C94_n689, Z => mult_28_C94_n559);
   mult_28_C94_U496 : OAI22D1 port map( A1 => mult_28_C94_n39, A2 => 
                           mult_28_C94_n687, B1 => mult_28_C94_n41, B2 => 
                           mult_28_C94_n688, Z => mult_28_C94_n558);
   mult_28_C94_U495 : OAI22D1 port map( A1 => mult_28_C94_n39, A2 => 
                           mult_28_C94_n686, B1 => mult_28_C94_n41, B2 => 
                           mult_28_C94_n687, Z => mult_28_C94_n557);
   mult_28_C94_U494 : OAI22D1 port map( A1 => mult_28_C94_n39, A2 => 
                           mult_28_C94_n685, B1 => mult_28_C94_n41, B2 => 
                           mult_28_C94_n686, Z => mult_28_C94_n556);
   mult_28_C94_U493 : OAI22D1 port map( A1 => mult_28_C94_n39, A2 => 
                           mult_28_C94_n684, B1 => mult_28_C94_n41, B2 => 
                           mult_28_C94_n685, Z => mult_28_C94_n555);
   mult_28_C94_U492 : OAI22D1 port map( A1 => mult_28_C94_n39, A2 => 
                           mult_28_C94_n683, B1 => mult_28_C94_n41, B2 => 
                           mult_28_C94_n684, Z => mult_28_C94_n554);
   mult_28_C94_U491 : OAI22D1 port map( A1 => mult_28_C94_n40, A2 => 
                           mult_28_C94_n682, B1 => mult_28_C94_n42, B2 => 
                           mult_28_C94_n683, Z => mult_28_C94_n553);
   mult_28_C94_U490 : OAI22D1 port map( A1 => mult_28_C94_n40, A2 => 
                           mult_28_C94_n681, B1 => mult_28_C94_n42, B2 => 
                           mult_28_C94_n682, Z => mult_28_C94_n552);
   mult_28_C94_U489 : OAI22D1 port map( A1 => mult_28_C94_n40, A2 => 
                           mult_28_C94_n680, B1 => mult_28_C94_n42, B2 => 
                           mult_28_C94_n681, Z => mult_28_C94_n551);
   mult_28_C94_U488 : OAI22D1 port map( A1 => mult_28_C94_n40, A2 => 
                           mult_28_C94_n679, B1 => mult_28_C94_n42, B2 => 
                           mult_28_C94_n680, Z => mult_28_C94_n550);
   mult_28_C94_U487 : OAI22D1 port map( A1 => mult_28_C94_n40, A2 => 
                           mult_28_C94_n678, B1 => mult_28_C94_n42, B2 => 
                           mult_28_C94_n679, Z => mult_28_C94_n549);
   mult_28_C94_U486 : OAI22D1 port map( A1 => mult_28_C94_n40, A2 => 
                           mult_28_C94_n677, B1 => mult_28_C94_n42, B2 => 
                           mult_28_C94_n678, Z => mult_28_C94_n548);
   mult_28_C94_U485 : OAI22D1 port map( A1 => mult_28_C94_n40, A2 => 
                           mult_28_C94_n676, B1 => mult_28_C94_n42, B2 => 
                           mult_28_C94_n677, Z => mult_28_C94_n319);
   mult_28_C94_U482 : NAN2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C94_n43, Z => mult_28_C94_n675);
   mult_28_C94_U481 : EXNOR2D1 port map( A1 => mult_28_C94_n43, A2 => 
                           data_in(0), Z => mult_28_C94_n674);
   mult_28_C94_U480 : EXNOR2D1 port map( A1 => mult_28_C94_n43, A2 => 
                           mult_28_C94_n809, Z => mult_28_C94_n673);
   mult_28_C94_U479 : EXNOR2D1 port map( A1 => mult_28_C94_n43, A2 => 
                           mult_28_C94_n808, Z => mult_28_C94_n672);
   mult_28_C94_U478 : EXNOR2D1 port map( A1 => mult_28_C94_n43, A2 => 
                           mult_28_C94_n807, Z => mult_28_C94_n671);
   mult_28_C94_U477 : EXNOR2D1 port map( A1 => mult_28_C94_n43, A2 => 
                           mult_28_C94_n806, Z => mult_28_C94_n670);
   mult_28_C94_U476 : EXNOR2D1 port map( A1 => mult_28_C94_n43, A2 => 
                           mult_28_C94_n805, Z => mult_28_C94_n669);
   mult_28_C94_U475 : EXNOR2D1 port map( A1 => mult_28_C94_n43, A2 => 
                           data_in(6), Z => mult_28_C94_n668);
   mult_28_C94_U474 : EXNOR2D1 port map( A1 => mult_28_C94_n43, A2 => 
                           mult_28_C94_n803, Z => mult_28_C94_n667);
   mult_28_C94_U473 : EXNOR2D1 port map( A1 => mult_28_C94_n43, A2 => 
                           mult_28_C94_n802, Z => mult_28_C94_n666);
   mult_28_C94_U472 : EXNOR2D1 port map( A1 => mult_28_C94_n43, A2 => 
                           mult_28_C94_n801, Z => mult_28_C94_n665);
   mult_28_C94_U471 : EXNOR2D1 port map( A1 => mult_28_C94_n43, A2 => 
                           mult_28_C94_n800, Z => mult_28_C94_n664);
   mult_28_C94_U470 : EXNOR2D1 port map( A1 => mult_28_C94_n43, A2 => 
                           mult_28_C94_n799, Z => mult_28_C94_n663);
   mult_28_C94_U469 : EXNOR2D1 port map( A1 => mult_28_C94_n43, A2 => 
                           mult_28_C94_n798, Z => mult_28_C94_n662);
   mult_28_C94_U468 : EXNOR2D1 port map( A1 => mult_28_C94_n43, A2 => 
                           mult_28_C94_n797, Z => mult_28_C94_n661);
   mult_28_C94_U467 : EXNOR2D1 port map( A1 => mult_28_C94_n43, A2 => 
                           mult_28_C94_n796, Z => mult_28_C94_n660);
   mult_28_C94_U466 : EXNOR2D1 port map( A1 => mult_28_C94_n43, A2 => 
                           mult_28_C94_n795, Z => mult_28_C94_n659);
   mult_28_C94_U465 : NOR2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C94_n45, Z => mult_28_C94_n546);
   mult_28_C94_U464 : OAI22D1 port map( A1 => mult_28_C94_n45, A2 => 
                           mult_28_C94_n673, B1 => mult_28_C94_n47, B2 => 
                           mult_28_C94_n674, Z => mult_28_C94_n545);
   mult_28_C94_U463 : OAI22D1 port map( A1 => mult_28_C94_n45, A2 => 
                           mult_28_C94_n672, B1 => mult_28_C94_n47, B2 => 
                           mult_28_C94_n673, Z => mult_28_C94_n544);
   mult_28_C94_U462 : OAI22D1 port map( A1 => mult_28_C94_n45, A2 => 
                           mult_28_C94_n671, B1 => mult_28_C94_n47, B2 => 
                           mult_28_C94_n672, Z => mult_28_C94_n543);
   mult_28_C94_U461 : OAI22D1 port map( A1 => mult_28_C94_n45, A2 => 
                           mult_28_C94_n670, B1 => mult_28_C94_n47, B2 => 
                           mult_28_C94_n671, Z => mult_28_C94_n542);
   mult_28_C94_U460 : OAI22D1 port map( A1 => mult_28_C94_n45, A2 => 
                           mult_28_C94_n669, B1 => mult_28_C94_n47, B2 => 
                           mult_28_C94_n670, Z => mult_28_C94_n541);
   mult_28_C94_U459 : OAI22D1 port map( A1 => mult_28_C94_n45, A2 => 
                           mult_28_C94_n668, B1 => mult_28_C94_n47, B2 => 
                           mult_28_C94_n669, Z => mult_28_C94_n540);
   mult_28_C94_U458 : OAI22D1 port map( A1 => mult_28_C94_n45, A2 => 
                           mult_28_C94_n667, B1 => mult_28_C94_n47, B2 => 
                           mult_28_C94_n668, Z => mult_28_C94_n539);
   mult_28_C94_U457 : OAI22D1 port map( A1 => mult_28_C94_n45, A2 => 
                           mult_28_C94_n666, B1 => mult_28_C94_n47, B2 => 
                           mult_28_C94_n667, Z => mult_28_C94_n538);
   mult_28_C94_U456 : OAI22D1 port map( A1 => mult_28_C94_n46, A2 => 
                           mult_28_C94_n665, B1 => mult_28_C94_n48, B2 => 
                           mult_28_C94_n666, Z => mult_28_C94_n537);
   mult_28_C94_U455 : OAI22D1 port map( A1 => mult_28_C94_n46, A2 => 
                           mult_28_C94_n664, B1 => mult_28_C94_n48, B2 => 
                           mult_28_C94_n665, Z => mult_28_C94_n536);
   mult_28_C94_U454 : OAI22D1 port map( A1 => mult_28_C94_n46, A2 => 
                           mult_28_C94_n663, B1 => mult_28_C94_n48, B2 => 
                           mult_28_C94_n664, Z => mult_28_C94_n535);
   mult_28_C94_U453 : OAI22D1 port map( A1 => mult_28_C94_n46, A2 => 
                           mult_28_C94_n662, B1 => mult_28_C94_n48, B2 => 
                           mult_28_C94_n663, Z => mult_28_C94_n534);
   mult_28_C94_U452 : OAI22D1 port map( A1 => mult_28_C94_n46, A2 => 
                           mult_28_C94_n661, B1 => mult_28_C94_n48, B2 => 
                           mult_28_C94_n662, Z => mult_28_C94_n533);
   mult_28_C94_U451 : OAI22D1 port map( A1 => mult_28_C94_n46, A2 => 
                           mult_28_C94_n660, B1 => mult_28_C94_n48, B2 => 
                           mult_28_C94_n661, Z => mult_28_C94_n532);
   mult_28_C94_U447 : ADFULD1 port map( A => mult_28_C94_n655, B => 
                           mult_28_C94_n626, CI => mult_28_C94_n640, CO => 
                           mult_28_C94_n519, S => mult_28_C94_n520);
   mult_28_C94_U445 : ADFULD1 port map( A => mult_28_C94_n625, B => 
                           mult_28_C94_n639, CI => mult_28_C94_n518, CO => 
                           mult_28_C94_n515, S => mult_28_C94_n516);
   mult_28_C94_U444 : ADFULD1 port map( A => mult_28_C94_n653, B => 
                           mult_28_C94_n610, CI => mult_28_C94_n638, CO => 
                           mult_28_C94_n513, S => mult_28_C94_n514);
   mult_28_C94_U443 : ADFULD1 port map( A => mult_28_C94_n517, B => 
                           mult_28_C94_n624, CI => mult_28_C94_n514, CO => 
                           mult_28_C94_n511, S => mult_28_C94_n512);
   mult_28_C94_U441 : ADFULD1 port map( A => mult_28_C94_n609, B => 
                           mult_28_C94_n637, CI => mult_28_C94_n623, CO => 
                           mult_28_C94_n507, S => mult_28_C94_n508);
   mult_28_C94_U440 : ADFULD1 port map( A => mult_28_C94_n513, B => 
                           mult_28_C94_n510, CI => mult_28_C94_n508, CO => 
                           mult_28_C94_n505, S => mult_28_C94_n506);
   mult_28_C94_U439 : ADFULD1 port map( A => mult_28_C94_n651, B => 
                           mult_28_C94_n594, CI => mult_28_C94_n636, CO => 
                           mult_28_C94_n503, S => mult_28_C94_n504);
   mult_28_C94_U438 : ADFULD1 port map( A => mult_28_C94_n608, B => 
                           mult_28_C94_n622, CI => mult_28_C94_n509, CO => 
                           mult_28_C94_n501, S => mult_28_C94_n502);
   mult_28_C94_U437 : ADFULD1 port map( A => mult_28_C94_n504, B => 
                           mult_28_C94_n507, CI => mult_28_C94_n502, CO => 
                           mult_28_C94_n499, S => mult_28_C94_n500);
   mult_28_C94_U435 : ADFULD1 port map( A => mult_28_C94_n593, B => 
                           mult_28_C94_n607, CI => mult_28_C94_n621, CO => 
                           mult_28_C94_n495, S => mult_28_C94_n496);
   mult_28_C94_U434 : ADFULD1 port map( A => mult_28_C94_n498, B => 
                           mult_28_C94_n635, CI => mult_28_C94_n503, CO => 
                           mult_28_C94_n493, S => mult_28_C94_n494);
   mult_28_C94_U433 : ADFULD1 port map( A => mult_28_C94_n496, B => 
                           mult_28_C94_n501, CI => mult_28_C94_n494, CO => 
                           mult_28_C94_n491, S => mult_28_C94_n492);
   mult_28_C94_U432 : ADFULD1 port map( A => mult_28_C94_n649, B => 
                           mult_28_C94_n578, CI => mult_28_C94_n634, CO => 
                           mult_28_C94_n489, S => mult_28_C94_n490);
   mult_28_C94_U431 : ADFULD1 port map( A => mult_28_C94_n592, B => 
                           mult_28_C94_n620, CI => mult_28_C94_n606, CO => 
                           mult_28_C94_n487, S => mult_28_C94_n488);
   mult_28_C94_U430 : ADFULD1 port map( A => mult_28_C94_n495, B => 
                           mult_28_C94_n497, CI => mult_28_C94_n490, CO => 
                           mult_28_C94_n485, S => mult_28_C94_n486);
   mult_28_C94_U429 : ADFULD1 port map( A => mult_28_C94_n493, B => 
                           mult_28_C94_n488, CI => mult_28_C94_n486, CO => 
                           mult_28_C94_n483, S => mult_28_C94_n484);
   mult_28_C94_U427 : ADFULD1 port map( A => mult_28_C94_n577, B => 
                           mult_28_C94_n605, CI => mult_28_C94_n633, CO => 
                           mult_28_C94_n479, S => mult_28_C94_n480);
   mult_28_C94_U426 : ADFULD1 port map( A => mult_28_C94_n591, B => 
                           mult_28_C94_n619, CI => mult_28_C94_n482, CO => 
                           mult_28_C94_n477, S => mult_28_C94_n478);
   mult_28_C94_U425 : ADFULD1 port map( A => mult_28_C94_n487, B => 
                           mult_28_C94_n489, CI => mult_28_C94_n480, CO => 
                           mult_28_C94_n475, S => mult_28_C94_n476);
   mult_28_C94_U424 : ADFULD1 port map( A => mult_28_C94_n485, B => 
                           mult_28_C94_n478, CI => mult_28_C94_n476, CO => 
                           mult_28_C94_n473, S => mult_28_C94_n474);
   mult_28_C94_U423 : ADFULD1 port map( A => mult_28_C94_n647, B => 
                           mult_28_C94_n562, CI => mult_28_C94_n632, CO => 
                           mult_28_C94_n471, S => mult_28_C94_n472);
   mult_28_C94_U422 : ADFULD1 port map( A => mult_28_C94_n576, B => 
                           mult_28_C94_n618, CI => mult_28_C94_n590, CO => 
                           mult_28_C94_n469, S => mult_28_C94_n470);
   mult_28_C94_U421 : ADFULD1 port map( A => mult_28_C94_n481, B => 
                           mult_28_C94_n604, CI => mult_28_C94_n479, CO => 
                           mult_28_C94_n467, S => mult_28_C94_n468);
   mult_28_C94_U420 : ADFULD1 port map( A => mult_28_C94_n470, B => 
                           mult_28_C94_n472, CI => mult_28_C94_n477, CO => 
                           mult_28_C94_n465, S => mult_28_C94_n466);
   mult_28_C94_U419 : ADFULD1 port map( A => mult_28_C94_n468, B => 
                           mult_28_C94_n475, CI => mult_28_C94_n466, CO => 
                           mult_28_C94_n463, S => mult_28_C94_n464);
   mult_28_C94_U418 : ADHALFD1 port map( A => mult_28_C94_n524, B => 
                           mult_28_C94_n646, CO => mult_28_C94_n461, S => 
                           mult_28_C94_n462);
   mult_28_C94_U417 : ADFULD1 port map( A => mult_28_C94_n631, B => 
                           mult_28_C94_n589, CI => mult_28_C94_n617, CO => 
                           mult_28_C94_n459, S => mult_28_C94_n460);
   mult_28_C94_U416 : ADFULD1 port map( A => mult_28_C94_n561, B => 
                           mult_28_C94_n603, CI => mult_28_C94_n575, CO => 
                           mult_28_C94_n457, S => mult_28_C94_n458);
   mult_28_C94_U415 : ADFULD1 port map( A => mult_28_C94_n471, B => 
                           mult_28_C94_n462, CI => mult_28_C94_n469, CO => 
                           mult_28_C94_n455, S => mult_28_C94_n456);
   mult_28_C94_U414 : ADFULD1 port map( A => mult_28_C94_n460, B => 
                           mult_28_C94_n458, CI => mult_28_C94_n467, CO => 
                           mult_28_C94_n453, S => mult_28_C94_n454);
   mult_28_C94_U413 : ADFULD1 port map( A => mult_28_C94_n465, B => 
                           mult_28_C94_n456, CI => mult_28_C94_n454, CO => 
                           mult_28_C94_n451, S => mult_28_C94_n452);
   mult_28_C94_U412 : ADFULD1 port map( A => mult_28_C94_n645, B => 
                           mult_28_C94_n546, CI => mult_28_C94_n630, CO => 
                           mult_28_C94_n449, S => mult_28_C94_n450);
   mult_28_C94_U411 : ADFULD1 port map( A => mult_28_C94_n560, B => 
                           mult_28_C94_n616, CI => mult_28_C94_n574, CO => 
                           mult_28_C94_n447, S => mult_28_C94_n448);
   mult_28_C94_U410 : ADFULD1 port map( A => mult_28_C94_n588, B => 
                           mult_28_C94_n602, CI => mult_28_C94_n461, CO => 
                           mult_28_C94_n445, S => mult_28_C94_n446);
   mult_28_C94_U409 : ADFULD1 port map( A => mult_28_C94_n457, B => 
                           mult_28_C94_n459, CI => mult_28_C94_n450, CO => 
                           mult_28_C94_n443, S => mult_28_C94_n444);
   mult_28_C94_U408 : ADFULD1 port map( A => mult_28_C94_n446, B => 
                           mult_28_C94_n448, CI => mult_28_C94_n455, CO => 
                           mult_28_C94_n441, S => mult_28_C94_n442);
   mult_28_C94_U407 : ADFULD1 port map( A => mult_28_C94_n453, B => 
                           mult_28_C94_n444, CI => mult_28_C94_n442, CO => 
                           mult_28_C94_n439, S => mult_28_C94_n440);
   mult_28_C94_U406 : ADHALFD1 port map( A => mult_28_C94_n523, B => 
                           mult_28_C94_n644, CO => mult_28_C94_n437, S => 
                           mult_28_C94_n438);
   mult_28_C94_U405 : ADFULD1 port map( A => mult_28_C94_n545, B => 
                           mult_28_C94_n587, CI => mult_28_C94_n559, CO => 
                           mult_28_C94_n435, S => mult_28_C94_n436);
   mult_28_C94_U404 : ADFULD1 port map( A => mult_28_C94_n629, B => 
                           mult_28_C94_n573, CI => mult_28_C94_n601, CO => 
                           mult_28_C94_n433, S => mult_28_C94_n434);
   mult_28_C94_U403 : ADFULD1 port map( A => mult_28_C94_n438, B => 
                           mult_28_C94_n615, CI => mult_28_C94_n449, CO => 
                           mult_28_C94_n431, S => mult_28_C94_n432);
   mult_28_C94_U402 : ADFULD1 port map( A => mult_28_C94_n445, B => 
                           mult_28_C94_n447, CI => mult_28_C94_n434, CO => 
                           mult_28_C94_n429, S => mult_28_C94_n430);
   mult_28_C94_U401 : ADFULD1 port map( A => mult_28_C94_n443, B => 
                           mult_28_C94_n436, CI => mult_28_C94_n432, CO => 
                           mult_28_C94_n427, S => mult_28_C94_n428);
   mult_28_C94_U400 : ADFULD1 port map( A => mult_28_C94_n441, B => 
                           mult_28_C94_n430, CI => mult_28_C94_n428, CO => 
                           mult_28_C94_n425, S => mult_28_C94_n426);
   mult_28_C94_U397 : ADFULD1 port map( A => mult_28_C94_n544, B => 
                           mult_28_C94_n586, CI => mult_28_C94_n572, CO => 
                           mult_28_C94_n421, S => mult_28_C94_n422);
   mult_28_C94_U396 : ADFULD1 port map( A => mult_28_C94_n614, B => 
                           mult_28_C94_n628, CI => mult_28_C94_n643, CO => 
                           mult_28_C94_n419, S => mult_28_C94_n420);
   mult_28_C94_U395 : ADFULD1 port map( A => mult_28_C94_n424, B => 
                           mult_28_C94_n437, CI => mult_28_C94_n435, CO => 
                           mult_28_C94_n417, S => mult_28_C94_n418);
   mult_28_C94_U394 : ADFULD1 port map( A => mult_28_C94_n422, B => 
                           mult_28_C94_n433, CI => mult_28_C94_n420, CO => 
                           mult_28_C94_n415, S => mult_28_C94_n416);
   mult_28_C94_U393 : ADFULD1 port map( A => mult_28_C94_n429, B => 
                           mult_28_C94_n431, CI => mult_28_C94_n418, CO => 
                           mult_28_C94_n413, S => mult_28_C94_n414);
   mult_28_C94_U392 : ADFULD1 port map( A => mult_28_C94_n427, B => 
                           mult_28_C94_n416, CI => mult_28_C94_n414, CO => 
                           mult_28_C94_n411, S => mult_28_C94_n412);
   mult_28_C94_U390 : ADFULD1 port map( A => mult_28_C94_n543, B => 
                           mult_28_C94_n571, CI => mult_28_C94_n613, CO => 
                           mult_28_C94_n407, S => mult_28_C94_n408);
   mult_28_C94_U389 : ADFULD1 port map( A => mult_28_C94_n557, B => 
                           mult_28_C94_n599, CI => mult_28_C94_n585, CO => 
                           mult_28_C94_n405, S => mult_28_C94_n406);
   mult_28_C94_U388 : ADFULD1 port map( A => mult_28_C94_n423, B => 
                           mult_28_C94_n410, CI => mult_28_C94_n421, CO => 
                           mult_28_C94_n403, S => mult_28_C94_n404);
   mult_28_C94_U387 : ADFULD1 port map( A => mult_28_C94_n406, B => 
                           mult_28_C94_n419, CI => mult_28_C94_n408, CO => 
                           mult_28_C94_n401, S => mult_28_C94_n402);
   mult_28_C94_U386 : ADFULD1 port map( A => mult_28_C94_n404, B => 
                           mult_28_C94_n417, CI => mult_28_C94_n415, CO => 
                           mult_28_C94_n399, S => mult_28_C94_n400);
   mult_28_C94_U385 : ADFULD1 port map( A => mult_28_C94_n413, B => 
                           mult_28_C94_n402, CI => mult_28_C94_n400, CO => 
                           mult_28_C94_n397, S => mult_28_C94_n398);
   mult_28_C94_U384 : ADFULD1 port map( A => mult_28_C94_n409, B => 
                           mult_28_C94_n542, CI => mult_28_C94_n556, CO => 
                           mult_28_C94_n395, S => mult_28_C94_n396);
   mult_28_C94_U383 : ADFULD1 port map( A => mult_28_C94_n570, B => 
                           mult_28_C94_n598, CI => mult_28_C94_n612, CO => 
                           mult_28_C94_n393, S => mult_28_C94_n394);
   mult_28_C94_U382 : ADFULD1 port map( A => mult_28_C94_n627, B => 
                           mult_28_C94_n584, CI => mult_28_C94_n407, CO => 
                           mult_28_C94_n391, S => mult_28_C94_n392);
   mult_28_C94_U381 : ADFULD1 port map( A => mult_28_C94_n394, B => 
                           mult_28_C94_n405, CI => mult_28_C94_n396, CO => 
                           mult_28_C94_n389, S => mult_28_C94_n390);
   mult_28_C94_U380 : ADFULD1 port map( A => mult_28_C94_n392, B => 
                           mult_28_C94_n403, CI => mult_28_C94_n401, CO => 
                           mult_28_C94_n387, S => mult_28_C94_n388);
   mult_28_C94_U379 : ADFULD1 port map( A => mult_28_C94_n399, B => 
                           mult_28_C94_n390, CI => mult_28_C94_n388, CO => 
                           mult_28_C94_n385, S => mult_28_C94_n386);
   mult_28_C94_U377 : ADFULD1 port map( A => mult_28_C94_n597, B => 
                           mult_28_C94_n569, CI => mult_28_C94_n583, CO => 
                           mult_28_C94_n381, S => mult_28_C94_n382);
   mult_28_C94_U376 : ADFULD1 port map( A => mult_28_C94_n541, B => 
                           mult_28_C94_n555, CI => mult_28_C94_n384, CO => 
                           mult_28_C94_n379, S => mult_28_C94_n380);
   mult_28_C94_U375 : ADFULD1 port map( A => mult_28_C94_n393, B => 
                           mult_28_C94_n395, CI => mult_28_C94_n382, CO => 
                           mult_28_C94_n377, S => mult_28_C94_n378);
   mult_28_C94_U374 : ADFULD1 port map( A => mult_28_C94_n391, B => 
                           mult_28_C94_n380, CI => mult_28_C94_n389, CO => 
                           mult_28_C94_n375, S => mult_28_C94_n376);
   mult_28_C94_U373 : ADFULD1 port map( A => mult_28_C94_n387, B => 
                           mult_28_C94_n378, CI => mult_28_C94_n376, CO => 
                           mult_28_C94_n373, S => mult_28_C94_n374);
   mult_28_C94_U372 : ADFULD1 port map( A => mult_28_C94_n383, B => 
                           mult_28_C94_n540, CI => mult_28_C94_n568, CO => 
                           mult_28_C94_n371, S => mult_28_C94_n372);
   mult_28_C94_U371 : ADFULD1 port map( A => mult_28_C94_n554, B => 
                           mult_28_C94_n582, CI => mult_28_C94_n596, CO => 
                           mult_28_C94_n369, S => mult_28_C94_n370);
   mult_28_C94_U370 : ADFULD1 port map( A => mult_28_C94_n381, B => 
                           mult_28_C94_n611, CI => mult_28_C94_n379, CO => 
                           mult_28_C94_n367, S => mult_28_C94_n368);
   mult_28_C94_U369 : ADFULD1 port map( A => mult_28_C94_n372, B => 
                           mult_28_C94_n370, CI => mult_28_C94_n377, CO => 
                           mult_28_C94_n365, S => mult_28_C94_n366);
   mult_28_C94_U368 : ADFULD1 port map( A => mult_28_C94_n375, B => 
                           mult_28_C94_n368, CI => mult_28_C94_n366, CO => 
                           mult_28_C94_n363, S => mult_28_C94_n364);
   mult_28_C94_U366 : ADFULD1 port map( A => mult_28_C94_n581, B => 
                           mult_28_C94_n553, CI => mult_28_C94_n539, CO => 
                           mult_28_C94_n359, S => mult_28_C94_n360);
   mult_28_C94_U365 : ADFULD1 port map( A => mult_28_C94_n362, B => 
                           mult_28_C94_n567, CI => mult_28_C94_n371, CO => 
                           mult_28_C94_n357, S => mult_28_C94_n358);
   mult_28_C94_U364 : ADFULD1 port map( A => mult_28_C94_n360, B => 
                           mult_28_C94_n369, CI => mult_28_C94_n367, CO => 
                           mult_28_C94_n355, S => mult_28_C94_n356);
   mult_28_C94_U363 : ADFULD1 port map( A => mult_28_C94_n365, B => 
                           mult_28_C94_n358, CI => mult_28_C94_n356, CO => 
                           mult_28_C94_n353, S => mult_28_C94_n354);
   mult_28_C94_U362 : ADFULD1 port map( A => mult_28_C94_n580, B => 
                           mult_28_C94_n538, CI => mult_28_C94_n361, CO => 
                           mult_28_C94_n351, S => mult_28_C94_n352);
   mult_28_C94_U361 : ADFULD1 port map( A => mult_28_C94_n566, B => 
                           mult_28_C94_n552, CI => mult_28_C94_n595, CO => 
                           mult_28_C94_n349, S => mult_28_C94_n350);
   mult_28_C94_U360 : ADFULD1 port map( A => mult_28_C94_n352, B => 
                           mult_28_C94_n359, CI => mult_28_C94_n350, CO => 
                           mult_28_C94_n347, S => mult_28_C94_n348);
   mult_28_C94_U359 : ADFULD1 port map( A => mult_28_C94_n348, B => 
                           mult_28_C94_n357, CI => mult_28_C94_n355, CO => 
                           mult_28_C94_n345, S => mult_28_C94_n346);
   mult_28_C94_U357 : ADFULD1 port map( A => mult_28_C94_n551, B => 
                           mult_28_C94_n537, CI => mult_28_C94_n565, CO => 
                           mult_28_C94_n341, S => mult_28_C94_n342);
   mult_28_C94_U356 : ADFULD1 port map( A => mult_28_C94_n351, B => 
                           mult_28_C94_n344, CI => mult_28_C94_n349, CO => 
                           mult_28_C94_n339, S => mult_28_C94_n340);
   mult_28_C94_U355 : ADFULD1 port map( A => mult_28_C94_n347, B => 
                           mult_28_C94_n342, CI => mult_28_C94_n340, CO => 
                           mult_28_C94_n337, S => mult_28_C94_n338);
   mult_28_C94_U354 : ADFULD1 port map( A => mult_28_C94_n550, B => 
                           mult_28_C94_n536, CI => mult_28_C94_n343, CO => 
                           mult_28_C94_n335, S => mult_28_C94_n336);
   mult_28_C94_U353 : ADFULD1 port map( A => mult_28_C94_n579, B => 
                           mult_28_C94_n564, CI => mult_28_C94_n341, CO => 
                           mult_28_C94_n333, S => mult_28_C94_n334);
   mult_28_C94_U352 : ADFULD1 port map( A => mult_28_C94_n339, B => 
                           mult_28_C94_n336, CI => mult_28_C94_n334, CO => 
                           mult_28_C94_n331, S => mult_28_C94_n332);
   mult_28_C94_U350 : ADFULD1 port map( A => mult_28_C94_n535, B => 
                           mult_28_C94_n549, CI => mult_28_C94_n330, CO => 
                           mult_28_C94_n327, S => mult_28_C94_n328);
   mult_28_C94_U349 : ADFULD1 port map( A => mult_28_C94_n328, B => 
                           mult_28_C94_n335, CI => mult_28_C94_n333, CO => 
                           mult_28_C94_n325, S => mult_28_C94_n326);
   mult_28_C94_U348 : ADFULD1 port map( A => mult_28_C94_n548, B => 
                           mult_28_C94_n329, CI => mult_28_C94_n534, CO => 
                           mult_28_C94_n323, S => mult_28_C94_n324);
   mult_28_C94_U347 : ADFULD1 port map( A => mult_28_C94_n327, B => 
                           mult_28_C94_n563, CI => mult_28_C94_n324, CO => 
                           mult_28_C94_n321, S => mult_28_C94_n322);
   mult_28_C94_U345 : ADFULD1 port map( A => mult_28_C94_n320, B => 
                           mult_28_C94_n533, CI => mult_28_C94_n323, CO => 
                           mult_28_C94_n317, S => mult_28_C94_n318);
   mult_28_C94_U344 : ADFULD1 port map( A => mult_28_C94_n532, B => 
                           mult_28_C94_n319, CI => mult_28_C94_n547, CO => 
                           mult_28_C94_n315, S => mult_28_C94_n316);
   mult_28_C94_U330 : AOI21D1 port map( A1 => mult_28_C94_n937, A2 => 
                           mult_28_C94_n939, B => mult_28_C94_n938, Z => 
                           mult_28_C94_n277);
   mult_28_C94_U324 : OAI21D1 port map( A1 => mult_28_C94_n275, A2 => 
                           mult_28_C94_n277, B => mult_28_C94_n276, Z => 
                           mult_28_C94_n274);
   mult_28_C94_U316 : AOI21D1 port map( A1 => mult_28_C94_n274, A2 => 
                           mult_28_C94_n935, B => mult_28_C94_n936, Z => 
                           mult_28_C94_n269);
   mult_28_C94_U310 : OAI21D1 port map( A1 => mult_28_C94_n267, A2 => 
                           mult_28_C94_n269, B => mult_28_C94_n268, Z => 
                           mult_28_C94_n266);
   mult_28_C94_U302 : AOI21D1 port map( A1 => mult_28_C94_n266, A2 => 
                           mult_28_C94_n933, B => mult_28_C94_n934, Z => 
                           mult_28_C94_n261);
   mult_28_C94_U285 : AOI21D1 port map( A1 => mult_28_C94_n926, A2 => 
                           mult_28_C94_n929, B => mult_28_C94_n927, Z => 
                           mult_28_C94_n250);
   mult_28_C94_U283 : OAI21D1 port map( A1 => mult_28_C94_n249, A2 => 
                           mult_28_C94_n261, B => mult_28_C94_n250, Z => 
                           mult_28_C94_n248);
   mult_28_C94_U275 : AOI21D1 port map( A1 => mult_28_C94_n248, A2 => 
                           mult_28_C94_n928, B => mult_28_C94_n931, Z => 
                           mult_28_C94_n243);
   mult_28_C94_U258 : AOI21D1 port map( A1 => mult_28_C94_n921, A2 => 
                           mult_28_C94_n923, B => mult_28_C94_n924, Z => 
                           mult_28_C94_n232);
   mult_28_C94_U256 : OAI21D1 port map( A1 => mult_28_C94_n243, A2 => 
                           mult_28_C94_n231, B => mult_28_C94_n232, Z => 
                           mult_28_C94_n230);
   mult_28_C94_U237 : AOI21D1 port map( A1 => mult_28_C94_n925, A2 => 
                           mult_28_C94_n910, B => mult_28_C94_n917, Z => 
                           mult_28_C94_n217);
   mult_28_C94_U232 : NOR2D2 port map( A1 => mult_28_C94_n440, A2 => 
                           mult_28_C94_n451, Z => mult_28_C94_n213);
   mult_28_C94_U225 : EXNOR2D1 port map( A1 => mult_28_C94_n215, A2 => 
                           mult_28_C94_n69, Z => m4_0);
   mult_28_C94_U224 : NAN2D2 port map( A1 => mult_28_C94_n426, A2 => 
                           mult_28_C94_n439, Z => mult_28_C94_n208);
   mult_28_C94_U223 : NOR2D2 port map( A1 => mult_28_C94_n426, A2 => 
                           mult_28_C94_n439, Z => mult_28_C94_n207);
   mult_28_C94_U218 : AOI21D1 port map( A1 => mult_28_C94_n209, A2 => 
                           mult_28_C94_n205, B => mult_28_C94_n206, Z => 
                           mult_28_C94_n204);
   mult_28_C94_U217 : EXNOR2D1 port map( A1 => mult_28_C94_n209, A2 => 
                           mult_28_C94_n68, Z => m4_1);
   mult_28_C94_U215 : NOR2D2 port map( A1 => mult_28_C94_n412, A2 => 
                           mult_28_C94_n425, Z => mult_28_C94_n202);
   mult_28_C94_U212 : OAI21D1 port map( A1 => mult_28_C94_n202, A2 => 
                           mult_28_C94_n208, B => mult_28_C94_n203, Z => 
                           mult_28_C94_n201);
   mult_28_C94_U205 : EXOR2D1 port map( A1 => mult_28_C94_n204, A2 => 
                           mult_28_C94_n67, Z => m4_2);
   mult_28_C94_U203 : NOR2D2 port map( A1 => mult_28_C94_n398, A2 => 
                           mult_28_C94_n411, Z => mult_28_C94_n193);
   mult_28_C94_U198 : OAI21D1 port map( A1 => mult_28_C94_n199, A2 => 
                           mult_28_C94_n191, B => mult_28_C94_n194, Z => 
                           mult_28_C94_n190);
   mult_28_C94_U195 : EXOR2D1 port map( A1 => mult_28_C94_n195, A2 => 
                           mult_28_C94_n66, Z => m4_3);
   mult_28_C94_U193 : NOR2D2 port map( A1 => mult_28_C94_n386, A2 => 
                           mult_28_C94_n397, Z => mult_28_C94_n186);
   mult_28_C94_U190 : OAI21D1 port map( A1 => mult_28_C94_n186, A2 => 
                           mult_28_C94_n194, B => mult_28_C94_n187, Z => 
                           mult_28_C94_n185);
   mult_28_C94_U188 : AOI21D1 port map( A1 => mult_28_C94_n201, A2 => 
                           mult_28_C94_n184, B => mult_28_C94_n185, Z => 
                           mult_28_C94_n183);
   mult_28_C94_U186 : OAI21D1 port map( A1 => mult_28_C94_n182, A2 => 
                           mult_28_C94_n210, B => mult_28_C94_n183, Z => 
                           mult_28_C94_n181);
   mult_28_C94_U185 : EXOR2D1 port map( A1 => mult_28_C94_n188, A2 => 
                           mult_28_C94_n65, Z => m4_4);
   mult_28_C94_U184 : NAN2D2 port map( A1 => mult_28_C94_n374, A2 => 
                           mult_28_C94_n385, Z => mult_28_C94_n180);
   mult_28_C94_U178 : AOI21D1 port map( A1 => mult_28_C94_n51, A2 => 
                           mult_28_C94_n177, B => mult_28_C94_n178, Z => 
                           mult_28_C94_n176);
   mult_28_C94_U177 : EXNOR2D1 port map( A1 => mult_28_C94_n51, A2 => 
                           mult_28_C94_n64, Z => m4_5);
   mult_28_C94_U175 : NOR2D2 port map( A1 => mult_28_C94_n364, A2 => 
                           mult_28_C94_n373, Z => mult_28_C94_n174);
   mult_28_C94_U172 : OAI21D1 port map( A1 => mult_28_C94_n174, A2 => 
                           mult_28_C94_n180, B => mult_28_C94_n175, Z => 
                           mult_28_C94_n173);
   mult_28_C94_U166 : AOI21D1 port map( A1 => mult_28_C94_n51, A2 => 
                           mult_28_C94_n168, B => mult_28_C94_n173, Z => 
                           mult_28_C94_n167);
   mult_28_C94_U163 : NOR2D2 port map( A1 => mult_28_C94_n354, A2 => 
                           mult_28_C94_n363, Z => mult_28_C94_n165);
   mult_28_C94_U156 : OAI21D1 port map( A1 => mult_28_C94_n171, A2 => 
                           mult_28_C94_n161, B => mult_28_C94_n162, Z => 
                           mult_28_C94_n160);
   mult_28_C94_U153 : EXOR2D1 port map( A1 => mult_28_C94_n167, A2 => 
                           mult_28_C94_n62, Z => m4_7);
   mult_28_C94_U144 : AOI21D1 port map( A1 => mult_28_C94_n164, A2 => 
                           mult_28_C94_n152, B => mult_28_C94_n155, Z => 
                           mult_28_C94_n151);
   mult_28_C94_U142 : OAI21D1 port map( A1 => mult_28_C94_n171, A2 => 
                           mult_28_C94_n150, B => mult_28_C94_n151, Z => 
                           mult_28_C94_n149);
   mult_28_C94_U139 : EXOR2D1 port map( A1 => mult_28_C94_n158, A2 => 
                           mult_28_C94_n61, Z => m4_8);
   mult_28_C94_U137 : NOR2D2 port map( A1 => mult_28_C94_n338, A2 => 
                           mult_28_C94_n345, Z => mult_28_C94_n145);
   mult_28_C94_U132 : AOI21D1 port map( A1 => mult_28_C94_n155, A2 => 
                           mult_28_C94_n143, B => mult_28_C94_n144, Z => 
                           mult_28_C94_n142);
   mult_28_C94_U123 : EXOR2D1 port map( A1 => mult_28_C94_n147, A2 => 
                           mult_28_C94_n60, Z => m4_9);
   mult_28_C94_U116 : OAI21D1 port map( A1 => mult_28_C94_n913, A2 => 
                           mult_28_C94_n132, B => mult_28_C94_n133, Z => 
                           mult_28_C94_n129);
   mult_28_C94_U113 : EXOR2D1 port map( A1 => mult_28_C94_n134, A2 => 
                           mult_28_C94_n59, Z => m4_10);
   mult_28_C94_U108 : OAI21D1 port map( A1 => mult_28_C94_n133, A2 => 
                           mult_28_C94_n125, B => mult_28_C94_n126, Z => 
                           mult_28_C94_n124);
   mult_28_C94_U97 : EXOR2D1 port map( A1 => mult_28_C94_n127, A2 => 
                           mult_28_C94_n58, Z => m4_11);
   mult_28_C94_U88 : OAI21D1 port map( A1 => mult_28_C94_n913, A2 => 
                           mult_28_C94_n108, B => mult_28_C94_n109, Z => 
                           mult_28_C94_n107);
   mult_28_C94_U85 : EXOR2D1 port map( A1 => mult_28_C94_n114, A2 => 
                           mult_28_C94_n57, Z => m4_12);
   mult_28_C94_U80 : OAI21D1 port map( A1 => mult_28_C94_n113, A2 => 
                           mult_28_C94_n103, B => mult_28_C94_n104, Z => 
                           mult_28_C94_n102);
   mult_28_C94_U78 : AOI21D1 port map( A1 => mult_28_C94_n124, A2 => 
                           mult_28_C94_n101, B => mult_28_C94_n102, Z => 
                           mult_28_C94_n100);
   mult_28_C94_U74 : OAI21D1 port map( A1 => mult_28_C94_n913, A2 => 
                           mult_28_C94_n99, B => mult_28_C94_n100, Z => 
                           mult_28_C94_n96);
   mult_28_C94_U71 : EXOR2D1 port map( A1 => mult_28_C94_n105, A2 => 
                           mult_28_C94_n56, Z => m4_13);
   mult_28_C94_U62 : OAI21D1 port map( A1 => mult_28_C94_n913, A2 => 
                           mult_28_C94_n920, B => mult_28_C94_n919, Z => 
                           mult_28_C94_n87);
   mult_28_C94_U60 : AOI21D1 port map( A1 => mult_28_C94_n51, A2 => 
                           mult_28_C94_n86, B => mult_28_C94_n87, Z => 
                           mult_28_C94_n85);
   mult_28_C94_U59 : EXOR2D1 port map( A1 => mult_28_C94_n94, A2 => 
                           mult_28_C94_n55, Z => m4_14);
   mult_28_C94_U54 : EXOR2D1 port map( A1 => mult_28_C94_n85, A2 => 
                           mult_28_C94_n54, Z => m4_15);
   mult_28_C93_U1012 : BUFD1 port map( A => coeff_memory_63_port, Z => 
                           mult_28_C93_n43);
   mult_28_C93_U1011 : BUFD1 port map( A => coeff_memory_61_port, Z => 
                           mult_28_C93_n37);
   mult_28_C93_U1010 : BUFD1 port map( A => coeff_memory_51_port, Z => 
                           mult_28_C93_n7);
   mult_28_C93_U1009 : BUFD1 port map( A => coeff_memory_49_port, Z => 
                           mult_28_C93_n1);
   mult_28_C93_U1008 : BUFD1 port map( A => coeff_memory_57_port, Z => 
                           mult_28_C93_n25);
   mult_28_C93_U1007 : BUFD1 port map( A => coeff_memory_53_port, Z => 
                           mult_28_C93_n13);
   mult_28_C93_U1006 : BUFD1 port map( A => coeff_memory_59_port, Z => 
                           mult_28_C93_n31);
   mult_28_C93_U1005 : BUFD1 port map( A => coeff_memory_55_port, Z => 
                           mult_28_C93_n19);
   mult_28_C93_U1004 : INVD1 port map( A => coeff_memory_48_port, Z => 
                           mult_28_C93_n834);
   mult_28_C93_U1003 : NAN2D1 port map( A1 => mult_28_C93_n818, A2 => 
                           mult_28_C93_n834, Z => mult_28_C93_n826);
   mult_28_C93_U1002 : OAI22M10D1 port map( A1 => mult_28_C93_n7, A2 => 
                           mult_28_C93_n12, B1 => mult_28_C93_n10, B2 => 
                           mult_28_C93_n777, Z => mult_28_C93_n529);
   mult_28_C93_U1001 : ADHALFDL port map( A => mult_28_C93_n641, B => 
                           mult_28_C93_n656, CO => mult_28_C93_n521, S => 
                           mult_28_C93_n522);
   mult_28_C93_U1000 : BUFD1 port map( A => data_in(15), Z => mult_28_C93_n795)
                           ;
   mult_28_C93_U999 : BUFD1 port map( A => data_in(12), Z => mult_28_C93_n798);
   mult_28_C93_U998 : BUFD1 port map( A => data_in(13), Z => mult_28_C93_n797);
   mult_28_C93_U997 : BUFD1 port map( A => data_in(14), Z => mult_28_C93_n796);
   mult_28_C93_U996 : BUFD1 port map( A => data_in(11), Z => mult_28_C93_n799);
   mult_28_C93_U995 : BUFD1 port map( A => data_in(3), Z => mult_28_C93_n807);
   mult_28_C93_U994 : BUFD1 port map( A => data_in(7), Z => mult_28_C93_n803);
   mult_28_C93_U993 : BUFD1 port map( A => data_in(2), Z => mult_28_C93_n808);
   mult_28_C93_U992 : BUFD1 port map( A => data_in(8), Z => mult_28_C93_n802);
   mult_28_C93_U991 : BUFD1 port map( A => data_in(4), Z => mult_28_C93_n806);
   mult_28_C93_U990 : BUFD1 port map( A => data_in(1), Z => mult_28_C93_n809);
   mult_28_C93_U989 : OA22D1 port map( A1 => mult_28_C93_n46, A2 => 
                           mult_28_C93_n659, B1 => mult_28_C93_n48, B2 => 
                           mult_28_C93_n660, Z => mult_28_C93_n938);
   mult_28_C93_U988 : INVD1 port map( A => mult_28_C93_n1, Z => 
                           mult_28_C93_n842);
   mult_28_C93_U987 : BUFD1 port map( A => mult_28_C93_n834, Z => 
                           mult_28_C93_n3);
   mult_28_C93_U986 : BUFD1 port map( A => mult_28_C93_n834, Z => 
                           mult_28_C93_n4);
   mult_28_C93_U985 : BUFD1 port map( A => mult_28_C93_n832, Z => 
                           mult_28_C93_n16);
   mult_28_C93_U984 : BUFD1 port map( A => mult_28_C93_n827, Z => 
                           mult_28_C93_n46);
   mult_28_C93_U983 : BUFD1 port map( A => mult_28_C93_n828, Z => 
                           mult_28_C93_n40);
   mult_28_C93_U982 : BUFD1 port map( A => mult_28_C93_n826, Z => 
                           mult_28_C93_n5);
   mult_28_C93_U981 : BUFD1 port map( A => mult_28_C93_n827, Z => 
                           mult_28_C93_n45);
   mult_28_C93_U980 : BUFD1 port map( A => mult_28_C93_n826, Z => 
                           mult_28_C93_n6);
   mult_28_C93_U979 : BUFD1 port map( A => mult_28_C93_n828, Z => 
                           mult_28_C93_n39);
   mult_28_C93_U978 : BUFD1 port map( A => mult_28_C93_n829, Z => 
                           mult_28_C93_n34);
   mult_28_C93_U977 : BUFD1 port map( A => mult_28_C93_n830, Z => 
                           mult_28_C93_n28);
   mult_28_C93_U976 : BUFD1 port map( A => mult_28_C93_n833, Z => 
                           mult_28_C93_n9);
   mult_28_C93_U975 : BUFD1 port map( A => mult_28_C93_n819, Z => 
                           mult_28_C93_n47);
   mult_28_C93_U974 : BUFD1 port map( A => mult_28_C93_n833, Z => 
                           mult_28_C93_n10);
   mult_28_C93_U973 : BUFD1 port map( A => mult_28_C93_n831, Z => 
                           mult_28_C93_n22);
   mult_28_C93_U972 : BUFD1 port map( A => mult_28_C93_n830, Z => 
                           mult_28_C93_n27);
   mult_28_C93_U971 : BUFD1 port map( A => mult_28_C93_n832, Z => 
                           mult_28_C93_n15);
   mult_28_C93_U970 : BUFD1 port map( A => mult_28_C93_n829, Z => 
                           mult_28_C93_n33);
   mult_28_C93_U969 : BUFD1 port map( A => mult_28_C93_n831, Z => 
                           mult_28_C93_n21);
   mult_28_C93_U968 : BUFD1 port map( A => mult_28_C93_n824, Z => 
                           mult_28_C93_n18);
   mult_28_C93_U967 : BUFD1 port map( A => mult_28_C93_n820, Z => 
                           mult_28_C93_n42);
   mult_28_C93_U966 : BUFD1 port map( A => mult_28_C93_n819, Z => 
                           mult_28_C93_n48);
   mult_28_C93_U965 : BUFD1 port map( A => mult_28_C93_n820, Z => 
                           mult_28_C93_n41);
   mult_28_C93_U964 : BUFD1 port map( A => mult_28_C93_n821, Z => 
                           mult_28_C93_n36);
   mult_28_C93_U963 : BUFD1 port map( A => mult_28_C93_n825, Z => 
                           mult_28_C93_n11);
   mult_28_C93_U962 : BUFD1 port map( A => mult_28_C93_n822, Z => 
                           mult_28_C93_n30);
   mult_28_C93_U961 : BUFD1 port map( A => mult_28_C93_n823, Z => 
                           mult_28_C93_n24);
   mult_28_C93_U960 : BUFD1 port map( A => mult_28_C93_n822, Z => 
                           mult_28_C93_n29);
   mult_28_C93_U959 : BUFD1 port map( A => mult_28_C93_n825, Z => 
                           mult_28_C93_n12);
   mult_28_C93_U958 : BUFD1 port map( A => mult_28_C93_n824, Z => 
                           mult_28_C93_n17);
   mult_28_C93_U957 : BUFD1 port map( A => mult_28_C93_n821, Z => 
                           mult_28_C93_n35);
   mult_28_C93_U956 : BUFD1 port map( A => mult_28_C93_n823, Z => 
                           mult_28_C93_n23);
   mult_28_C93_U955 : AND2D1 port map( A1 => mult_28_C93_n658, A2 => 
                           mult_28_C93_n530, Z => mult_28_C93_n937);
   mult_28_C93_U954 : NOR2D1 port map( A1 => mult_28_C93_n522, A2 => 
                           mult_28_C93_n529, Z => mult_28_C93_n275);
   mult_28_C93_U953 : OAI22M10D1 port map( A1 => mult_28_C93_n37, A2 => 
                           mult_28_C93_n42, B1 => mult_28_C93_n40, B2 => 
                           mult_28_C93_n692, Z => mult_28_C93_n524);
   mult_28_C93_U952 : INVD1 port map( A => mult_28_C93_n13, Z => 
                           mult_28_C93_n840);
   mult_28_C93_U951 : ADHALFDL port map( A => mult_28_C93_n528, B => 
                           mult_28_C93_n654, CO => mult_28_C93_n517, S => 
                           mult_28_C93_n518);
   mult_28_C93_U950 : AND2DL port map( A1 => mult_28_C93_n520, A2 => 
                           mult_28_C93_n521, Z => mult_28_C93_n934);
   mult_28_C93_U949 : OAI22M10D1 port map( A1 => mult_28_C93_n43, A2 => 
                           mult_28_C93_n48, B1 => mult_28_C93_n46, B2 => 
                           mult_28_C93_n675, Z => mult_28_C93_n523);
   mult_28_C93_U948 : OR2D1 port map( A1 => mult_28_C93_n520, A2 => 
                           mult_28_C93_n521, Z => mult_28_C93_n933);
   mult_28_C93_U947 : NAN2DL port map( A1 => mult_28_C93_n516, A2 => 
                           mult_28_C93_n519, Z => mult_28_C93_n268);
   mult_28_C93_U946 : INVD1 port map( A => mult_28_C93_n31, Z => 
                           mult_28_C93_n837);
   mult_28_C93_U945 : ADHALFDL port map( A => mult_28_C93_n525, B => 
                           mult_28_C93_n648, CO => mult_28_C93_n481, S => 
                           mult_28_C93_n482);
   mult_28_C93_U944 : INVD1 port map( A => mult_28_C93_n25, Z => 
                           mult_28_C93_n838);
   mult_28_C93_U943 : ADHALFDL port map( A => mult_28_C93_n526, B => 
                           mult_28_C93_n650, CO => mult_28_C93_n497, S => 
                           mult_28_C93_n498);
   mult_28_C93_U942 : INVD1 port map( A => mult_28_C93_n19, Z => 
                           mult_28_C93_n839);
   mult_28_C93_U941 : ADHALFDL port map( A => mult_28_C93_n527, B => 
                           mult_28_C93_n652, CO => mult_28_C93_n509, S => 
                           mult_28_C93_n510);
   mult_28_C93_U940 : OR2D1 port map( A1 => mult_28_C93_n315, A2 => 
                           mult_28_C93_n938, Z => mult_28_C93_n930);
   mult_28_C93_U939 : AO21D1 port map( A1 => mult_28_C93_n42, A2 => 
                           mult_28_C93_n40, B => mult_28_C93_n676, Z => 
                           mult_28_C93_n547);
   mult_28_C93_U938 : INVD1 port map( A => mult_28_C93_n319, Z => 
                           mult_28_C93_n320);
   mult_28_C93_U937 : AO21D1 port map( A1 => mult_28_C93_n36, A2 => 
                           mult_28_C93_n34, B => mult_28_C93_n693, Z => 
                           mult_28_C93_n563);
   mult_28_C93_U936 : INVDL port map( A => mult_28_C93_n329, Z => 
                           mult_28_C93_n330);
   mult_28_C93_U935 : AO21D1 port map( A1 => mult_28_C93_n30, A2 => 
                           mult_28_C93_n28, B => mult_28_C93_n710, Z => 
                           mult_28_C93_n579);
   mult_28_C93_U934 : NAN2D1 port map( A1 => mult_28_C93_n315, A2 => 
                           mult_28_C93_n938, Z => mult_28_C93_n84);
   mult_28_C93_U933 : NAN2D1 port map( A1 => mult_28_C93_n930, A2 => 
                           mult_28_C93_n84, Z => mult_28_C93_n54);
   mult_28_C93_U932 : INVDL port map( A => mult_28_C93_n361, Z => 
                           mult_28_C93_n362);
   mult_28_C93_U931 : AO21D1 port map( A1 => mult_28_C93_n24, A2 => 
                           mult_28_C93_n22, B => mult_28_C93_n727, Z => 
                           mult_28_C93_n595);
   mult_28_C93_U930 : AO21D1 port map( A1 => mult_28_C93_n18, A2 => 
                           mult_28_C93_n16, B => mult_28_C93_n744, Z => 
                           mult_28_C93_n611);
   mult_28_C93_U929 : AO21D1 port map( A1 => mult_28_C93_n6, A2 => 
                           mult_28_C93_n4, B => mult_28_C93_n778, Z => 
                           mult_28_C93_n643);
   mult_28_C93_U928 : AO21D1 port map( A1 => mult_28_C93_n12, A2 => 
                           mult_28_C93_n10, B => mult_28_C93_n761, Z => 
                           mult_28_C93_n627);
   mult_28_C93_U927 : INVDL port map( A => mult_28_C93_n383, Z => 
                           mult_28_C93_n384);
   mult_28_C93_U926 : EXNOR2D1 port map( A1 => mult_28_C93_n600, A2 => 
                           mult_28_C93_n558, Z => mult_28_C93_n424);
   mult_28_C93_U925 : AND2DL port map( A1 => mult_28_C93_n492, A2 => 
                           mult_28_C93_n499, Z => mult_28_C93_n929);
   mult_28_C93_U924 : AND2D1 port map( A1 => mult_28_C93_n506, A2 => 
                           mult_28_C93_n511, Z => mult_28_C93_n927);
   mult_28_C93_U923 : OR2D1 port map( A1 => mult_28_C93_n492, A2 => 
                           mult_28_C93_n499, Z => mult_28_C93_n926);
   mult_28_C93_U922 : AND2DL port map( A1 => mult_28_C93_n500, A2 => 
                           mult_28_C93_n505, Z => mult_28_C93_n925);
   mult_28_C93_U921 : OR2D1 port map( A1 => mult_28_C93_n500, A2 => 
                           mult_28_C93_n505, Z => mult_28_C93_n924);
   mult_28_C93_U920 : NAN2D1 port map( A1 => mult_28_C93_n317, A2 => 
                           mult_28_C93_n316, Z => mult_28_C93_n93);
   mult_28_C93_U919 : NOR2D1 port map( A1 => mult_28_C93_n317, A2 => 
                           mult_28_C93_n316, Z => mult_28_C93_n92);
   mult_28_C93_U918 : NAN2DL port map( A1 => mult_28_C93_n318, A2 => 
                           mult_28_C93_n321, Z => mult_28_C93_n104);
   mult_28_C93_U917 : NOR2D1 port map( A1 => mult_28_C93_n318, A2 => 
                           mult_28_C93_n321, Z => mult_28_C93_n103);
   mult_28_C93_U916 : NOR2D1 port map( A1 => mult_28_C93_n325, A2 => 
                           mult_28_C93_n322, Z => mult_28_C93_n112);
   mult_28_C93_U915 : INVDL port map( A => mult_28_C93_n343, Z => 
                           mult_28_C93_n344);
   mult_28_C93_U914 : NAN2DL port map( A1 => mult_28_C93_n440, A2 => 
                           mult_28_C93_n451, Z => mult_28_C93_n214);
   mult_28_C93_U913 : NAN2D1 port map( A1 => mult_28_C93_n923, A2 => 
                           mult_28_C93_n915, Z => mult_28_C93_n216);
   mult_28_C93_U912 : OR2D1 port map( A1 => mult_28_C93_n452, A2 => 
                           mult_28_C93_n463, Z => mult_28_C93_n923);
   mult_28_C93_U911 : AND2DL port map( A1 => mult_28_C93_n474, A2 => 
                           mult_28_C93_n483, Z => mult_28_C93_n922);
   mult_28_C93_U910 : OR2D1 port map( A1 => mult_28_C93_n484, A2 => 
                           mult_28_C93_n491, Z => mult_28_C93_n920);
   mult_28_C93_U909 : OR2D1 port map( A1 => mult_28_C93_n474, A2 => 
                           mult_28_C93_n483, Z => mult_28_C93_n919);
   mult_28_C93_U908 : NOR2D1 port map( A1 => mult_28_C93_n112, A2 => 
                           mult_28_C93_n103, Z => mult_28_C93_n101);
   mult_28_C93_U907 : NAN2DL port map( A1 => mult_28_C93_n326, A2 => 
                           mult_28_C93_n331, Z => mult_28_C93_n126);
   mult_28_C93_U906 : NOR2D1 port map( A1 => mult_28_C93_n326, A2 => 
                           mult_28_C93_n331, Z => mult_28_C93_n125);
   mult_28_C93_U905 : NAN2DL port map( A1 => mult_28_C93_n332, A2 => 
                           mult_28_C93_n337, Z => mult_28_C93_n133);
   mult_28_C93_U904 : OA21DL port map( A1 => mult_28_C93_n100, A2 => 
                           mult_28_C93_n92, B => mult_28_C93_n93, Z => 
                           mult_28_C93_n917);
   mult_28_C93_U903 : INVDL port map( A => mult_28_C93_n208, Z => 
                           mult_28_C93_n206);
   mult_28_C93_U902 : INVDL port map( A => mult_28_C93_n207, Z => 
                           mult_28_C93_n205);
   mult_28_C93_U901 : NAN2D1 port map( A1 => mult_28_C93_n338, A2 => 
                           mult_28_C93_n345, Z => mult_28_C93_n146);
   mult_28_C93_U900 : NAN2D1 port map( A1 => mult_28_C93_n354, A2 => 
                           mult_28_C93_n363, Z => mult_28_C93_n166);
   mult_28_C93_U899 : INVDL port map( A => mult_28_C93_n230, Z => 
                           mult_28_C93_n229);
   mult_28_C93_U898 : NOR2DL port map( A1 => mult_28_C93_n911, A2 => 
                           mult_28_C93_n918, Z => mult_28_C93_n86);
   mult_28_C93_U897 : INVDL port map( A => mult_28_C93_n132, Z => 
                           mult_28_C93_n131);
   mult_28_C93_U896 : INVD1 port map( A => mult_28_C93_n131, Z => 
                           mult_28_C93_n130);
   mult_28_C93_U895 : INVDL port map( A => mult_28_C93_n193, Z => 
                           mult_28_C93_n192);
   mult_28_C93_U894 : INVDL port map( A => mult_28_C93_n165, Z => 
                           mult_28_C93_n163);
   mult_28_C93_U893 : INVD1 port map( A => mult_28_C93_n157, Z => 
                           mult_28_C93_n155);
   mult_28_C93_U892 : INVDL port map( A => mult_28_C93_n201, Z => 
                           mult_28_C93_n199);
   mult_28_C93_U891 : INVD1 port map( A => mult_28_C93_n145, Z => 
                           mult_28_C93_n143);
   mult_28_C93_U890 : NOR2D1 port map( A1 => mult_28_C93_n179, A2 => 
                           mult_28_C93_n174, Z => mult_28_C93_n172);
   mult_28_C93_U889 : NOR2D1 port map( A1 => mult_28_C93_n374, A2 => 
                           mult_28_C93_n385, Z => mult_28_C93_n179);
   mult_28_C93_U888 : NOR2D1 port map( A1 => mult_28_C93_n141, A2 => 
                           mult_28_C93_n165, Z => mult_28_C93_n139);
   mult_28_C93_U887 : INVDL port map( A => mult_28_C93_n186, Z => 
                           mult_28_C93_n296);
   mult_28_C93_U886 : INVDL port map( A => mult_28_C93_n202, Z => 
                           mult_28_C93_n298);
   mult_28_C93_U885 : INVDL port map( A => mult_28_C93_n193, Z => 
                           mult_28_C93_n297);
   mult_28_C93_U884 : INVD1 port map( A => mult_28_C93_n210, Z => 
                           mult_28_C93_n209);
   mult_28_C93_U883 : INVDL port map( A => mult_28_C93_n174, Z => 
                           mult_28_C93_n294);
   mult_28_C93_U882 : AND2D1 port map( A1 => mult_28_C93_n292, A2 => 
                           mult_28_C93_n157, Z => mult_28_C93_n916);
   mult_28_C93_U881 : EXNOR2D1 port map( A1 => mult_28_C93_n158, A2 => 
                           mult_28_C93_n916, Z => m2_8);
   mult_28_C93_U880 : NAN2DL port map( A1 => mult_28_C93_n200, A2 => 
                           mult_28_C93_n184, Z => mult_28_C93_n182);
   mult_28_C93_U879 : BUFD4 port map( A => mult_28_C93_n181, Z => 
                           mult_28_C93_n51);
   mult_28_C93_U878 : INVD1 port map( A => mult_28_C93_n99, Z => 
                           mult_28_C93_n98);
   mult_28_C93_U877 : INVD1 port map( A => mult_28_C93_n98, Z => 
                           mult_28_C93_n97);
   mult_28_C93_U876 : INVDL port map( A => mult_28_C93_n180, Z => 
                           mult_28_C93_n178);
   mult_28_C93_U875 : NOR2DL port map( A1 => mult_28_C93_n911, A2 => 
                           mult_28_C93_n108, Z => mult_28_C93_n106);
   mult_28_C93_U874 : INVD1 port map( A => mult_28_C93_n156, Z => 
                           mult_28_C93_n152);
   mult_28_C93_U873 : NAN2D1 port map( A1 => mult_28_C93_n163, A2 => 
                           mult_28_C93_n152, Z => mult_28_C93_n150);
   mult_28_C93_U872 : NOR2D1 port map( A1 => mult_28_C93_n198, A2 => 
                           mult_28_C93_n191, Z => mult_28_C93_n189);
   mult_28_C93_U871 : NOR2DL port map( A1 => mult_28_C93_n911, A2 => 
                           mult_28_C93_n130, Z => mult_28_C93_n128);
   mult_28_C93_U870 : INVDL port map( A => mult_28_C93_n173, Z => 
                           mult_28_C93_n171);
   mult_28_C93_U869 : NAN2D1 port map( A1 => mult_28_C93_n292, A2 => 
                           mult_28_C93_n143, Z => mult_28_C93_n141);
   mult_28_C93_U868 : INVD1 port map( A => mult_28_C93_n52, Z => 
                           mult_28_C93_n136);
   mult_28_C93_U867 : INVD1 port map( A => mult_28_C93_n123, Z => 
                           mult_28_C93_n117);
   mult_28_C93_U866 : INVD1 port map( A => mult_28_C93_n170, Z => 
                           mult_28_C93_n168);
   mult_28_C93_U865 : NOR2D1 port map( A1 => mult_28_C93_n170, A2 => 
                           mult_28_C93_n161, Z => mult_28_C93_n159);
   mult_28_C93_U864 : INVD1 port map( A => mult_28_C93_n911, Z => 
                           mult_28_C93_n135);
   mult_28_C93_U863 : NAN2DL port map( A1 => mult_28_C93_n522, A2 => 
                           mult_28_C93_n529, Z => mult_28_C93_n276);
   mult_28_C93_U862 : NOR2D1 port map( A1 => mult_28_C93_n516, A2 => 
                           mult_28_C93_n519, Z => mult_28_C93_n267);
   mult_28_C93_U861 : OAI22DL port map( A1 => mult_28_C93_n778, A2 => 
                           mult_28_C93_n4, B1 => mult_28_C93_n6, B2 => 
                           mult_28_C93_n779, Z => mult_28_C93_n644);
   mult_28_C93_U860 : OR2DL port map( A1 => mult_28_C93_n506, A2 => 
                           mult_28_C93_n511, Z => mult_28_C93_n928);
   mult_28_C93_U859 : NAN2DL port map( A1 => mult_28_C93_n325, A2 => 
                           mult_28_C93_n322, Z => mult_28_C93_n113);
   mult_28_C93_U858 : AND2D1 port map( A1 => mult_28_C93_n484, A2 => 
                           mult_28_C93_n491, Z => mult_28_C93_n921);
   mult_28_C93_U857 : NAN2DL port map( A1 => mult_28_C93_n919, A2 => 
                           mult_28_C93_n920, Z => mult_28_C93_n231);
   mult_28_C93_U856 : OR2D1 port map( A1 => mult_28_C93_n464, A2 => 
                           mult_28_C93_n473, Z => mult_28_C93_n915);
   mult_28_C93_U855 : OR2DL port map( A1 => mult_28_C93_n600, A2 => 
                           mult_28_C93_n558, Z => mult_28_C93_n423);
   mult_28_C93_U854 : AND2DL port map( A1 => mult_28_C93_n452, A2 => 
                           mult_28_C93_n463, Z => mult_28_C93_n914);
   mult_28_C93_U853 : OR2DL port map( A1 => mult_28_C93_n99, A2 => 
                           mult_28_C93_n92, Z => mult_28_C93_n918);
   mult_28_C93_U852 : NAN2M1D1 port map( A1 => mult_28_C93_n92, A2 => 
                           mult_28_C93_n93, Z => mult_28_C93_n55);
   mult_28_C93_U851 : OA21M20DL port map( A1 => mult_28_C93_n124, A2 => 
                           mult_28_C93_n110, B => mult_28_C93_n113, Z => 
                           mult_28_C93_n109);
   mult_28_C93_U850 : NAN2M1DL port map( A1 => mult_28_C93_n213, A2 => 
                           mult_28_C93_n214, Z => mult_28_C93_n69);
   mult_28_C93_U849 : NAN2M1D1 port map( A1 => mult_28_C93_n103, A2 => 
                           mult_28_C93_n104, Z => mult_28_C93_n56);
   mult_28_C93_U848 : NAN2M1DL port map( A1 => mult_28_C93_n112, A2 => 
                           mult_28_C93_n113, Z => mult_28_C93_n57);
   mult_28_C93_U847 : NAN2DL port map( A1 => mult_28_C93_n346, A2 => 
                           mult_28_C93_n353, Z => mult_28_C93_n157);
   mult_28_C93_U846 : NAN2M1DL port map( A1 => mult_28_C93_n207, A2 => 
                           mult_28_C93_n208, Z => mult_28_C93_n68);
   mult_28_C93_U845 : NAN2D1 port map( A1 => mult_28_C93_n364, A2 => 
                           mult_28_C93_n373, Z => mult_28_C93_n175);
   mult_28_C93_U844 : NAN2D1 port map( A1 => mult_28_C93_n386, A2 => 
                           mult_28_C93_n397, Z => mult_28_C93_n187);
   mult_28_C93_U843 : OAI21D1 port map( A1 => mult_28_C93_n217, A2 => 
                           mult_28_C93_n213, B => mult_28_C93_n214, Z => 
                           mult_28_C93_n913);
   mult_28_C93_U842 : NOR2DL port map( A1 => mult_28_C93_n216, A2 => 
                           mult_28_C93_n213, Z => mult_28_C93_n912);
   mult_28_C93_U841 : AOI21D1 port map( A1 => mult_28_C93_n912, A2 => 
                           mult_28_C93_n230, B => mult_28_C93_n913, Z => 
                           mult_28_C93_n210);
   mult_28_C93_U840 : NAN2D1 port map( A1 => mult_28_C93_n412, A2 => 
                           mult_28_C93_n425, Z => mult_28_C93_n203);
   mult_28_C93_U839 : NAN2DL port map( A1 => mult_28_C93_n123, A2 => 
                           mult_28_C93_n101, Z => mult_28_C93_n99);
   mult_28_C93_U838 : NOR2DL port map( A1 => mult_28_C93_n132, A2 => 
                           mult_28_C93_n125, Z => mult_28_C93_n123);
   mult_28_C93_U837 : INVDL port map( A => mult_28_C93_n166, Z => 
                           mult_28_C93_n164);
   mult_28_C93_U836 : INVDL port map( A => mult_28_C93_n146, Z => 
                           mult_28_C93_n144);
   mult_28_C93_U835 : INVD1 port map( A => mult_28_C93_n192, Z => 
                           mult_28_C93_n191);
   mult_28_C93_U834 : BUFD1 port map( A => mult_28_C93_n138, Z => 
                           mult_28_C93_n52);
   mult_28_C93_U833 : NAN2M1DL port map( A1 => mult_28_C93_n125, A2 => 
                           mult_28_C93_n126, Z => mult_28_C93_n58);
   mult_28_C93_U832 : NAN2M1DL port map( A1 => mult_28_C93_n132, A2 => 
                           mult_28_C93_n133, Z => mult_28_C93_n59);
   mult_28_C93_U831 : NAN2M1DL port map( A1 => mult_28_C93_n145, A2 => 
                           mult_28_C93_n146, Z => mult_28_C93_n60);
   mult_28_C93_U830 : INVDL port map( A => mult_28_C93_n165, Z => 
                           mult_28_C93_n293);
   mult_28_C93_U829 : INVDL port map( A => mult_28_C93_n163, Z => 
                           mult_28_C93_n161);
   mult_28_C93_U828 : AO21M20DL port map( A1 => mult_28_C93_n52, A2 => 
                           mult_28_C93_n117, B => mult_28_C93_n124, Z => 
                           mult_28_C93_n116);
   mult_28_C93_U827 : AO21M20DL port map( A1 => mult_28_C93_n171, A2 => 
                           mult_28_C93_n161, B => mult_28_C93_n164, Z => 
                           mult_28_C93_n160);
   mult_28_C93_U826 : INVDL port map( A => mult_28_C93_n179, Z => 
                           mult_28_C93_n177);
   mult_28_C93_U825 : INVDL port map( A => mult_28_C93_n199, Z => 
                           mult_28_C93_n197);
   mult_28_C93_U824 : NAN2M1DL port map( A1 => mult_28_C93_n179, A2 => 
                           mult_28_C93_n180, Z => mult_28_C93_n64);
   mult_28_C93_U823 : NOR2DL port map( A1 => mult_28_C93_n911, A2 => 
                           mult_28_C93_n97, Z => mult_28_C93_n95);
   mult_28_C93_U822 : NOR2DL port map( A1 => mult_28_C93_n911, A2 => 
                           mult_28_C93_n117, Z => mult_28_C93_n115);
   mult_28_C93_U821 : NOR2DL port map( A1 => mult_28_C93_n170, A2 => 
                           mult_28_C93_n150, Z => mult_28_C93_n148);
   mult_28_C93_U820 : INVDL port map( A => mult_28_C93_n171, Z => 
                           mult_28_C93_n169);
   mult_28_C93_U819 : AND2DL port map( A1 => mult_28_C93_n512, A2 => 
                           mult_28_C93_n515, Z => mult_28_C93_n932);
   mult_28_C93_U818 : OR2D1 port map( A1 => mult_28_C93_n512, A2 => 
                           mult_28_C93_n515, Z => mult_28_C93_n931);
   mult_28_C93_U817 : NAN2DL port map( A1 => mult_28_C93_n924, A2 => 
                           mult_28_C93_n928, Z => mult_28_C93_n249);
   mult_28_C93_U816 : AOI21D1 port map( A1 => mult_28_C93_n924, A2 => 
                           mult_28_C93_n927, B => mult_28_C93_n925, Z => 
                           mult_28_C93_n250);
   mult_28_C93_U815 : AOI21DL port map( A1 => mult_28_C93_n51, A2 => 
                           mult_28_C93_n95, B => mult_28_C93_n96, Z => 
                           mult_28_C93_n94);
   mult_28_C93_U814 : OAI21DL port map( A1 => mult_28_C93_n229, A2 => 
                           mult_28_C93_n216, B => mult_28_C93_n217, Z => 
                           mult_28_C93_n215);
   mult_28_C93_U813 : AOI21DL port map( A1 => mult_28_C93_n51, A2 => 
                           mult_28_C93_n106, B => mult_28_C93_n107, Z => 
                           mult_28_C93_n105);
   mult_28_C93_U812 : AOI21DL port map( A1 => mult_28_C93_n51, A2 => 
                           mult_28_C93_n115, B => mult_28_C93_n116, Z => 
                           mult_28_C93_n114);
   mult_28_C93_U811 : NAN2D1 port map( A1 => mult_28_C93_n398, A2 => 
                           mult_28_C93_n411, Z => mult_28_C93_n194);
   mult_28_C93_U810 : NAN2D1 port map( A1 => mult_28_C93_n123, A2 => 
                           mult_28_C93_n110, Z => mult_28_C93_n108);
   mult_28_C93_U809 : AOI21DL port map( A1 => mult_28_C93_n51, A2 => 
                           mult_28_C93_n135, B => mult_28_C93_n136, Z => 
                           mult_28_C93_n134);
   mult_28_C93_U808 : AOI21DL port map( A1 => mult_28_C93_n51, A2 => 
                           mult_28_C93_n148, B => mult_28_C93_n149, Z => 
                           mult_28_C93_n147);
   mult_28_C93_U807 : AOI21DL port map( A1 => mult_28_C93_n51, A2 => 
                           mult_28_C93_n128, B => mult_28_C93_n129, Z => 
                           mult_28_C93_n127);
   mult_28_C93_U806 : AOI21D1 port map( A1 => mult_28_C93_n51, A2 => 
                           mult_28_C93_n168, B => mult_28_C93_n169, Z => 
                           mult_28_C93_n167);
   mult_28_C93_U805 : NAN2DL port map( A1 => mult_28_C93_n172, A2 => 
                           mult_28_C93_n139, Z => mult_28_C93_n911);
   mult_28_C93_U804 : INVDL port map( A => mult_28_C93_n112, Z => 
                           mult_28_C93_n110);
   mult_28_C93_U803 : INVDL port map( A => mult_28_C93_n172, Z => 
                           mult_28_C93_n170);
   mult_28_C93_U802 : OR2DL port map( A1 => mult_28_C93_n657, A2 => 
                           mult_28_C93_n642, Z => mult_28_C93_n935);
   mult_28_C93_U801 : AND2D1 port map( A1 => mult_28_C93_n657, A2 => 
                           mult_28_C93_n642, Z => mult_28_C93_n936);
   mult_28_C93_U800 : BUFD20 port map( A => data_in(5), Z => mult_28_C93_n805);
   mult_28_C93_U799 : BUFD20 port map( A => data_in(9), Z => mult_28_C93_n801);
   mult_28_C93_U798 : BUFD20 port map( A => data_in(10), Z => mult_28_C93_n800)
                           ;
   mult_28_C93_U797 : NOR2D1 port map( A1 => mult_28_C93_n202, A2 => 
                           mult_28_C93_n207, Z => mult_28_C93_n200);
   mult_28_C93_U796 : INVD1 port map( A => mult_28_C93_n200, Z => 
                           mult_28_C93_n198);
   mult_28_C93_U795 : AND2D1 port map( A1 => mult_28_C93_n464, A2 => 
                           mult_28_C93_n473, Z => mult_28_C93_n910);
   mult_28_C93_U794 : INVDL port map( A => mult_28_C93_n156, Z => 
                           mult_28_C93_n292);
   mult_28_C93_U793 : NOR2D1 port map( A1 => mult_28_C93_n346, A2 => 
                           mult_28_C93_n353, Z => mult_28_C93_n156);
   mult_28_C93_U792 : NAN2DL port map( A1 => mult_28_C93_n296, A2 => 
                           mult_28_C93_n187, Z => mult_28_C93_n65);
   mult_28_C93_U791 : NOR2D1 port map( A1 => mult_28_C93_n193, A2 => 
                           mult_28_C93_n186, Z => mult_28_C93_n184);
   mult_28_C93_U790 : NAN2D1 port map( A1 => mult_28_C93_n426, A2 => 
                           mult_28_C93_n439, Z => mult_28_C93_n208);
   mult_28_C93_U789 : NAN2D1 port map( A1 => mult_28_C93_n811, A2 => 
                           mult_28_C93_n827, Z => mult_28_C93_n819);
   mult_28_C93_U788 : NAN2D1 port map( A1 => mult_28_C93_n812, A2 => 
                           mult_28_C93_n828, Z => mult_28_C93_n820);
   mult_28_C93_U787 : NOR2D1 port map( A1 => mult_28_C93_n338, A2 => 
                           mult_28_C93_n345, Z => mult_28_C93_n145);
   mult_28_C93_U786 : NAN2D1 port map( A1 => mult_28_C93_n814, A2 => 
                           mult_28_C93_n830, Z => mult_28_C93_n822);
   mult_28_C93_U785 : NAN2D1 port map( A1 => mult_28_C93_n816, A2 => 
                           mult_28_C93_n832, Z => mult_28_C93_n824);
   mult_28_C93_U784 : NAN2D1 port map( A1 => mult_28_C93_n815, A2 => 
                           mult_28_C93_n831, Z => mult_28_C93_n823);
   mult_28_C93_U783 : INVDL port map( A => mult_28_C93_n409, Z => 
                           mult_28_C93_n410);
   mult_28_C93_U782 : NAN2D1 port map( A1 => mult_28_C93_n817, A2 => 
                           mult_28_C93_n833, Z => mult_28_C93_n825);
   mult_28_C93_U781 : NAN2D1 port map( A1 => mult_28_C93_n813, A2 => 
                           mult_28_C93_n829, Z => mult_28_C93_n821);
   mult_28_C93_U780 : NAN2DL port map( A1 => mult_28_C93_n297, A2 => 
                           mult_28_C93_n194, Z => mult_28_C93_n66);
   mult_28_C93_U779 : NAN2DL port map( A1 => mult_28_C93_n298, A2 => 
                           mult_28_C93_n203, Z => mult_28_C93_n67);
   mult_28_C93_U778 : NAN2DL port map( A1 => mult_28_C93_n293, A2 => 
                           mult_28_C93_n166, Z => mult_28_C93_n62);
   mult_28_C93_U777 : NAN2DL port map( A1 => mult_28_C93_n294, A2 => 
                           mult_28_C93_n175, Z => mult_28_C93_n63);
   mult_28_C93_U773 : EXOR2D1 port map( A1 => coeff_memory_48_port, A2 => 
                           coeff_memory_49_port, Z => mult_28_C93_n818);
   mult_28_C93_U771 : EXNOR2D1 port map( A1 => coeff_memory_50_port, A2 => 
                           coeff_memory_49_port, Z => mult_28_C93_n833);
   mult_28_C93_U770 : EXOR2D1 port map( A1 => coeff_memory_50_port, A2 => 
                           coeff_memory_51_port, Z => mult_28_C93_n817);
   mult_28_C93_U768 : EXNOR2D1 port map( A1 => coeff_memory_52_port, A2 => 
                           coeff_memory_51_port, Z => mult_28_C93_n832);
   mult_28_C93_U767 : EXOR2D1 port map( A1 => coeff_memory_52_port, A2 => 
                           coeff_memory_53_port, Z => mult_28_C93_n816);
   mult_28_C93_U765 : EXNOR2D1 port map( A1 => coeff_memory_54_port, A2 => 
                           coeff_memory_53_port, Z => mult_28_C93_n831);
   mult_28_C93_U764 : EXOR2D1 port map( A1 => coeff_memory_54_port, A2 => 
                           coeff_memory_55_port, Z => mult_28_C93_n815);
   mult_28_C93_U762 : EXNOR2D1 port map( A1 => coeff_memory_56_port, A2 => 
                           coeff_memory_55_port, Z => mult_28_C93_n830);
   mult_28_C93_U761 : EXOR2D1 port map( A1 => coeff_memory_56_port, A2 => 
                           coeff_memory_57_port, Z => mult_28_C93_n814);
   mult_28_C93_U759 : EXNOR2D1 port map( A1 => coeff_memory_58_port, A2 => 
                           coeff_memory_57_port, Z => mult_28_C93_n829);
   mult_28_C93_U758 : EXOR2D1 port map( A1 => coeff_memory_58_port, A2 => 
                           coeff_memory_59_port, Z => mult_28_C93_n813);
   mult_28_C93_U756 : EXNOR2D1 port map( A1 => coeff_memory_60_port, A2 => 
                           coeff_memory_59_port, Z => mult_28_C93_n828);
   mult_28_C93_U755 : EXOR2D1 port map( A1 => coeff_memory_60_port, A2 => 
                           coeff_memory_61_port, Z => mult_28_C93_n812);
   mult_28_C93_U753 : EXNOR2D1 port map( A1 => coeff_memory_62_port, A2 => 
                           coeff_memory_61_port, Z => mult_28_C93_n827);
   mult_28_C93_U752 : EXOR2D1 port map( A1 => coeff_memory_62_port, A2 => 
                           coeff_memory_63_port, Z => mult_28_C93_n811);
   mult_28_C93_U727 : NAN2M1D1 port map( A1 => data_in(0), A2 => mult_28_C93_n1
                           , Z => mult_28_C93_n794);
   mult_28_C93_U726 : EXNOR2D1 port map( A1 => mult_28_C93_n1, A2 => data_in(0)
                           , Z => mult_28_C93_n793);
   mult_28_C93_U725 : EXNOR2D1 port map( A1 => mult_28_C93_n1, A2 => 
                           mult_28_C93_n809, Z => mult_28_C93_n792);
   mult_28_C93_U724 : EXNOR2D1 port map( A1 => mult_28_C93_n1, A2 => 
                           mult_28_C93_n808, Z => mult_28_C93_n791);
   mult_28_C93_U723 : EXNOR2D1 port map( A1 => mult_28_C93_n1, A2 => 
                           mult_28_C93_n807, Z => mult_28_C93_n790);
   mult_28_C93_U722 : EXNOR2D1 port map( A1 => mult_28_C93_n1, A2 => 
                           mult_28_C93_n806, Z => mult_28_C93_n789);
   mult_28_C93_U721 : EXNOR2D1 port map( A1 => mult_28_C93_n1, A2 => 
                           mult_28_C93_n805, Z => mult_28_C93_n788);
   mult_28_C93_U720 : EXNOR2D1 port map( A1 => mult_28_C93_n1, A2 => data_in(6)
                           , Z => mult_28_C93_n787);
   mult_28_C93_U719 : EXNOR2D1 port map( A1 => mult_28_C93_n1, A2 => 
                           mult_28_C93_n803, Z => mult_28_C93_n786);
   mult_28_C93_U718 : EXNOR2D1 port map( A1 => mult_28_C93_n1, A2 => 
                           mult_28_C93_n802, Z => mult_28_C93_n785);
   mult_28_C93_U717 : EXNOR2D1 port map( A1 => mult_28_C93_n1, A2 => 
                           mult_28_C93_n801, Z => mult_28_C93_n784);
   mult_28_C93_U716 : EXNOR2D1 port map( A1 => mult_28_C93_n1, A2 => 
                           mult_28_C93_n800, Z => mult_28_C93_n783);
   mult_28_C93_U715 : EXNOR2D1 port map( A1 => mult_28_C93_n1, A2 => 
                           mult_28_C93_n799, Z => mult_28_C93_n782);
   mult_28_C93_U714 : EXNOR2D1 port map( A1 => mult_28_C93_n1, A2 => 
                           mult_28_C93_n798, Z => mult_28_C93_n781);
   mult_28_C93_U713 : EXNOR2D1 port map( A1 => mult_28_C93_n1, A2 => 
                           mult_28_C93_n797, Z => mult_28_C93_n780);
   mult_28_C93_U712 : EXNOR2D1 port map( A1 => mult_28_C93_n1, A2 => 
                           mult_28_C93_n796, Z => mult_28_C93_n779);
   mult_28_C93_U711 : EXNOR2D1 port map( A1 => mult_28_C93_n1, A2 => 
                           mult_28_C93_n795, Z => mult_28_C93_n778);
   mult_28_C93_U709 : OAI22D1 port map( A1 => mult_28_C93_n792, A2 => 
                           mult_28_C93_n3, B1 => mult_28_C93_n5, B2 => 
                           mult_28_C93_n793, Z => mult_28_C93_n658);
   mult_28_C93_U708 : OAI22D1 port map( A1 => mult_28_C93_n791, A2 => 
                           mult_28_C93_n3, B1 => mult_28_C93_n5, B2 => 
                           mult_28_C93_n792, Z => mult_28_C93_n657);
   mult_28_C93_U707 : OAI22D1 port map( A1 => mult_28_C93_n790, A2 => 
                           mult_28_C93_n3, B1 => mult_28_C93_n5, B2 => 
                           mult_28_C93_n791, Z => mult_28_C93_n656);
   mult_28_C93_U706 : OAI22D1 port map( A1 => mult_28_C93_n789, A2 => 
                           mult_28_C93_n3, B1 => mult_28_C93_n5, B2 => 
                           mult_28_C93_n790, Z => mult_28_C93_n655);
   mult_28_C93_U705 : OAI22D1 port map( A1 => mult_28_C93_n788, A2 => 
                           mult_28_C93_n3, B1 => mult_28_C93_n5, B2 => 
                           mult_28_C93_n789, Z => mult_28_C93_n654);
   mult_28_C93_U704 : OAI22D1 port map( A1 => mult_28_C93_n787, A2 => 
                           mult_28_C93_n3, B1 => mult_28_C93_n5, B2 => 
                           mult_28_C93_n788, Z => mult_28_C93_n653);
   mult_28_C93_U703 : OAI22D1 port map( A1 => mult_28_C93_n786, A2 => 
                           mult_28_C93_n3, B1 => mult_28_C93_n5, B2 => 
                           mult_28_C93_n787, Z => mult_28_C93_n652);
   mult_28_C93_U702 : OAI22D1 port map( A1 => mult_28_C93_n785, A2 => 
                           mult_28_C93_n3, B1 => mult_28_C93_n5, B2 => 
                           mult_28_C93_n786, Z => mult_28_C93_n651);
   mult_28_C93_U701 : OAI22D1 port map( A1 => mult_28_C93_n784, A2 => 
                           mult_28_C93_n4, B1 => mult_28_C93_n6, B2 => 
                           mult_28_C93_n785, Z => mult_28_C93_n650);
   mult_28_C93_U700 : OAI22D1 port map( A1 => mult_28_C93_n783, A2 => 
                           mult_28_C93_n4, B1 => mult_28_C93_n6, B2 => 
                           mult_28_C93_n784, Z => mult_28_C93_n649);
   mult_28_C93_U699 : OAI22D1 port map( A1 => mult_28_C93_n782, A2 => 
                           mult_28_C93_n4, B1 => mult_28_C93_n6, B2 => 
                           mult_28_C93_n783, Z => mult_28_C93_n648);
   mult_28_C93_U698 : OAI22D1 port map( A1 => mult_28_C93_n781, A2 => 
                           mult_28_C93_n4, B1 => mult_28_C93_n6, B2 => 
                           mult_28_C93_n782, Z => mult_28_C93_n647);
   mult_28_C93_U697 : OAI22D1 port map( A1 => mult_28_C93_n780, A2 => 
                           mult_28_C93_n4, B1 => mult_28_C93_n6, B2 => 
                           mult_28_C93_n781, Z => mult_28_C93_n646);
   mult_28_C93_U696 : OAI22D1 port map( A1 => mult_28_C93_n779, A2 => 
                           mult_28_C93_n4, B1 => mult_28_C93_n6, B2 => 
                           mult_28_C93_n780, Z => mult_28_C93_n645);
   mult_28_C93_U693 : OAI22D1 port map( A1 => mult_28_C93_n794, A2 => 
                           mult_28_C93_n4, B1 => mult_28_C93_n6, B2 => 
                           mult_28_C93_n842, Z => mult_28_C93_n530);
   mult_28_C93_U692 : NAN2M1D1 port map( A1 => data_in(0), A2 => mult_28_C93_n7
                           , Z => mult_28_C93_n777);
   mult_28_C93_U691 : EXNOR2D1 port map( A1 => mult_28_C93_n7, A2 => data_in(0)
                           , Z => mult_28_C93_n776);
   mult_28_C93_U690 : EXNOR2D1 port map( A1 => mult_28_C93_n7, A2 => 
                           mult_28_C93_n809, Z => mult_28_C93_n775);
   mult_28_C93_U689 : EXNOR2D1 port map( A1 => mult_28_C93_n7, A2 => 
                           mult_28_C93_n808, Z => mult_28_C93_n774);
   mult_28_C93_U688 : EXNOR2D1 port map( A1 => mult_28_C93_n7, A2 => 
                           mult_28_C93_n807, Z => mult_28_C93_n773);
   mult_28_C93_U687 : EXNOR2D1 port map( A1 => mult_28_C93_n7, A2 => 
                           mult_28_C93_n806, Z => mult_28_C93_n772);
   mult_28_C93_U686 : EXNOR2D1 port map( A1 => mult_28_C93_n7, A2 => 
                           mult_28_C93_n805, Z => mult_28_C93_n771);
   mult_28_C93_U685 : EXNOR2D1 port map( A1 => mult_28_C93_n7, A2 => data_in(6)
                           , Z => mult_28_C93_n770);
   mult_28_C93_U684 : EXNOR2D1 port map( A1 => mult_28_C93_n7, A2 => 
                           mult_28_C93_n803, Z => mult_28_C93_n769);
   mult_28_C93_U683 : EXNOR2D1 port map( A1 => mult_28_C93_n7, A2 => 
                           mult_28_C93_n802, Z => mult_28_C93_n768);
   mult_28_C93_U682 : EXNOR2D1 port map( A1 => mult_28_C93_n7, A2 => 
                           mult_28_C93_n801, Z => mult_28_C93_n767);
   mult_28_C93_U681 : EXNOR2D1 port map( A1 => mult_28_C93_n7, A2 => 
                           mult_28_C93_n800, Z => mult_28_C93_n766);
   mult_28_C93_U680 : EXNOR2D1 port map( A1 => mult_28_C93_n7, A2 => 
                           mult_28_C93_n799, Z => mult_28_C93_n765);
   mult_28_C93_U679 : EXNOR2D1 port map( A1 => mult_28_C93_n7, A2 => 
                           mult_28_C93_n798, Z => mult_28_C93_n764);
   mult_28_C93_U678 : EXNOR2D1 port map( A1 => mult_28_C93_n7, A2 => 
                           mult_28_C93_n797, Z => mult_28_C93_n763);
   mult_28_C93_U677 : EXNOR2D1 port map( A1 => mult_28_C93_n7, A2 => 
                           mult_28_C93_n796, Z => mult_28_C93_n762);
   mult_28_C93_U676 : EXNOR2D1 port map( A1 => mult_28_C93_n7, A2 => 
                           mult_28_C93_n795, Z => mult_28_C93_n761);
   mult_28_C93_U675 : NOR2M1D1 port map( A1 => data_in(0), A2 => mult_28_C93_n9
                           , Z => mult_28_C93_n642);
   mult_28_C93_U674 : OAI22D1 port map( A1 => mult_28_C93_n9, A2 => 
                           mult_28_C93_n775, B1 => mult_28_C93_n11, B2 => 
                           mult_28_C93_n776, Z => mult_28_C93_n641);
   mult_28_C93_U673 : OAI22D1 port map( A1 => mult_28_C93_n9, A2 => 
                           mult_28_C93_n774, B1 => mult_28_C93_n11, B2 => 
                           mult_28_C93_n775, Z => mult_28_C93_n640);
   mult_28_C93_U672 : OAI22D1 port map( A1 => mult_28_C93_n9, A2 => 
                           mult_28_C93_n773, B1 => mult_28_C93_n11, B2 => 
                           mult_28_C93_n774, Z => mult_28_C93_n639);
   mult_28_C93_U671 : OAI22D1 port map( A1 => mult_28_C93_n9, A2 => 
                           mult_28_C93_n772, B1 => mult_28_C93_n11, B2 => 
                           mult_28_C93_n773, Z => mult_28_C93_n638);
   mult_28_C93_U670 : OAI22D1 port map( A1 => mult_28_C93_n9, A2 => 
                           mult_28_C93_n771, B1 => mult_28_C93_n11, B2 => 
                           mult_28_C93_n772, Z => mult_28_C93_n637);
   mult_28_C93_U669 : OAI22D1 port map( A1 => mult_28_C93_n9, A2 => 
                           mult_28_C93_n770, B1 => mult_28_C93_n11, B2 => 
                           mult_28_C93_n771, Z => mult_28_C93_n636);
   mult_28_C93_U668 : OAI22D1 port map( A1 => mult_28_C93_n9, A2 => 
                           mult_28_C93_n769, B1 => mult_28_C93_n11, B2 => 
                           mult_28_C93_n770, Z => mult_28_C93_n635);
   mult_28_C93_U667 : OAI22D1 port map( A1 => mult_28_C93_n9, A2 => 
                           mult_28_C93_n768, B1 => mult_28_C93_n11, B2 => 
                           mult_28_C93_n769, Z => mult_28_C93_n634);
   mult_28_C93_U666 : OAI22D1 port map( A1 => mult_28_C93_n10, A2 => 
                           mult_28_C93_n767, B1 => mult_28_C93_n12, B2 => 
                           mult_28_C93_n768, Z => mult_28_C93_n633);
   mult_28_C93_U665 : OAI22D1 port map( A1 => mult_28_C93_n10, A2 => 
                           mult_28_C93_n766, B1 => mult_28_C93_n12, B2 => 
                           mult_28_C93_n767, Z => mult_28_C93_n632);
   mult_28_C93_U664 : OAI22D1 port map( A1 => mult_28_C93_n10, A2 => 
                           mult_28_C93_n765, B1 => mult_28_C93_n12, B2 => 
                           mult_28_C93_n766, Z => mult_28_C93_n631);
   mult_28_C93_U663 : OAI22D1 port map( A1 => mult_28_C93_n10, A2 => 
                           mult_28_C93_n764, B1 => mult_28_C93_n12, B2 => 
                           mult_28_C93_n765, Z => mult_28_C93_n630);
   mult_28_C93_U662 : OAI22D1 port map( A1 => mult_28_C93_n10, A2 => 
                           mult_28_C93_n763, B1 => mult_28_C93_n12, B2 => 
                           mult_28_C93_n764, Z => mult_28_C93_n629);
   mult_28_C93_U661 : OAI22D1 port map( A1 => mult_28_C93_n10, A2 => 
                           mult_28_C93_n762, B1 => mult_28_C93_n12, B2 => 
                           mult_28_C93_n763, Z => mult_28_C93_n628);
   mult_28_C93_U660 : OAI22D1 port map( A1 => mult_28_C93_n10, A2 => 
                           mult_28_C93_n761, B1 => mult_28_C93_n12, B2 => 
                           mult_28_C93_n762, Z => mult_28_C93_n409);
   mult_28_C93_U657 : NAN2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C93_n13, Z => mult_28_C93_n760);
   mult_28_C93_U656 : EXNOR2D1 port map( A1 => mult_28_C93_n13, A2 => 
                           data_in(0), Z => mult_28_C93_n759);
   mult_28_C93_U655 : EXNOR2D1 port map( A1 => mult_28_C93_n13, A2 => 
                           mult_28_C93_n809, Z => mult_28_C93_n758);
   mult_28_C93_U654 : EXNOR2D1 port map( A1 => mult_28_C93_n13, A2 => 
                           mult_28_C93_n808, Z => mult_28_C93_n757);
   mult_28_C93_U653 : EXNOR2D1 port map( A1 => mult_28_C93_n13, A2 => 
                           mult_28_C93_n807, Z => mult_28_C93_n756);
   mult_28_C93_U652 : EXNOR2D1 port map( A1 => mult_28_C93_n13, A2 => 
                           mult_28_C93_n806, Z => mult_28_C93_n755);
   mult_28_C93_U651 : EXNOR2D1 port map( A1 => mult_28_C93_n13, A2 => 
                           mult_28_C93_n805, Z => mult_28_C93_n754);
   mult_28_C93_U650 : EXNOR2D1 port map( A1 => mult_28_C93_n13, A2 => 
                           data_in(6), Z => mult_28_C93_n753);
   mult_28_C93_U649 : EXNOR2D1 port map( A1 => mult_28_C93_n13, A2 => 
                           mult_28_C93_n803, Z => mult_28_C93_n752);
   mult_28_C93_U648 : EXNOR2D1 port map( A1 => mult_28_C93_n13, A2 => 
                           mult_28_C93_n802, Z => mult_28_C93_n751);
   mult_28_C93_U647 : EXNOR2D1 port map( A1 => mult_28_C93_n13, A2 => 
                           mult_28_C93_n801, Z => mult_28_C93_n750);
   mult_28_C93_U646 : EXNOR2D1 port map( A1 => mult_28_C93_n13, A2 => 
                           mult_28_C93_n800, Z => mult_28_C93_n749);
   mult_28_C93_U645 : EXNOR2D1 port map( A1 => mult_28_C93_n13, A2 => 
                           mult_28_C93_n799, Z => mult_28_C93_n748);
   mult_28_C93_U644 : EXNOR2D1 port map( A1 => mult_28_C93_n13, A2 => 
                           mult_28_C93_n798, Z => mult_28_C93_n747);
   mult_28_C93_U643 : EXNOR2D1 port map( A1 => mult_28_C93_n13, A2 => 
                           mult_28_C93_n797, Z => mult_28_C93_n746);
   mult_28_C93_U642 : EXNOR2D1 port map( A1 => mult_28_C93_n13, A2 => 
                           mult_28_C93_n796, Z => mult_28_C93_n745);
   mult_28_C93_U641 : EXNOR2D1 port map( A1 => mult_28_C93_n13, A2 => 
                           mult_28_C93_n795, Z => mult_28_C93_n744);
   mult_28_C93_U640 : NOR2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C93_n15, Z => mult_28_C93_n626);
   mult_28_C93_U639 : OAI22D1 port map( A1 => mult_28_C93_n15, A2 => 
                           mult_28_C93_n758, B1 => mult_28_C93_n17, B2 => 
                           mult_28_C93_n759, Z => mult_28_C93_n625);
   mult_28_C93_U638 : OAI22D1 port map( A1 => mult_28_C93_n15, A2 => 
                           mult_28_C93_n757, B1 => mult_28_C93_n17, B2 => 
                           mult_28_C93_n758, Z => mult_28_C93_n624);
   mult_28_C93_U637 : OAI22D1 port map( A1 => mult_28_C93_n15, A2 => 
                           mult_28_C93_n756, B1 => mult_28_C93_n17, B2 => 
                           mult_28_C93_n757, Z => mult_28_C93_n623);
   mult_28_C93_U636 : OAI22D1 port map( A1 => mult_28_C93_n15, A2 => 
                           mult_28_C93_n755, B1 => mult_28_C93_n17, B2 => 
                           mult_28_C93_n756, Z => mult_28_C93_n622);
   mult_28_C93_U635 : OAI22D1 port map( A1 => mult_28_C93_n15, A2 => 
                           mult_28_C93_n754, B1 => mult_28_C93_n17, B2 => 
                           mult_28_C93_n755, Z => mult_28_C93_n621);
   mult_28_C93_U634 : OAI22D1 port map( A1 => mult_28_C93_n15, A2 => 
                           mult_28_C93_n753, B1 => mult_28_C93_n17, B2 => 
                           mult_28_C93_n754, Z => mult_28_C93_n620);
   mult_28_C93_U633 : OAI22D1 port map( A1 => mult_28_C93_n15, A2 => 
                           mult_28_C93_n752, B1 => mult_28_C93_n17, B2 => 
                           mult_28_C93_n753, Z => mult_28_C93_n619);
   mult_28_C93_U632 : OAI22D1 port map( A1 => mult_28_C93_n15, A2 => 
                           mult_28_C93_n751, B1 => mult_28_C93_n17, B2 => 
                           mult_28_C93_n752, Z => mult_28_C93_n618);
   mult_28_C93_U631 : OAI22D1 port map( A1 => mult_28_C93_n16, A2 => 
                           mult_28_C93_n750, B1 => mult_28_C93_n18, B2 => 
                           mult_28_C93_n751, Z => mult_28_C93_n617);
   mult_28_C93_U630 : OAI22D1 port map( A1 => mult_28_C93_n16, A2 => 
                           mult_28_C93_n749, B1 => mult_28_C93_n18, B2 => 
                           mult_28_C93_n750, Z => mult_28_C93_n616);
   mult_28_C93_U629 : OAI22D1 port map( A1 => mult_28_C93_n16, A2 => 
                           mult_28_C93_n748, B1 => mult_28_C93_n18, B2 => 
                           mult_28_C93_n749, Z => mult_28_C93_n615);
   mult_28_C93_U628 : OAI22D1 port map( A1 => mult_28_C93_n16, A2 => 
                           mult_28_C93_n747, B1 => mult_28_C93_n18, B2 => 
                           mult_28_C93_n748, Z => mult_28_C93_n614);
   mult_28_C93_U627 : OAI22D1 port map( A1 => mult_28_C93_n16, A2 => 
                           mult_28_C93_n746, B1 => mult_28_C93_n18, B2 => 
                           mult_28_C93_n747, Z => mult_28_C93_n613);
   mult_28_C93_U626 : OAI22D1 port map( A1 => mult_28_C93_n16, A2 => 
                           mult_28_C93_n745, B1 => mult_28_C93_n18, B2 => 
                           mult_28_C93_n746, Z => mult_28_C93_n612);
   mult_28_C93_U625 : OAI22D1 port map( A1 => mult_28_C93_n16, A2 => 
                           mult_28_C93_n744, B1 => mult_28_C93_n18, B2 => 
                           mult_28_C93_n745, Z => mult_28_C93_n383);
   mult_28_C93_U623 : OAI22D1 port map( A1 => mult_28_C93_n16, A2 => 
                           mult_28_C93_n760, B1 => mult_28_C93_n18, B2 => 
                           mult_28_C93_n840, Z => mult_28_C93_n528);
   mult_28_C93_U622 : NAN2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C93_n19, Z => mult_28_C93_n743);
   mult_28_C93_U621 : EXNOR2D1 port map( A1 => mult_28_C93_n19, A2 => 
                           data_in(0), Z => mult_28_C93_n742);
   mult_28_C93_U620 : EXNOR2D1 port map( A1 => mult_28_C93_n19, A2 => 
                           mult_28_C93_n809, Z => mult_28_C93_n741);
   mult_28_C93_U619 : EXNOR2D1 port map( A1 => mult_28_C93_n19, A2 => 
                           mult_28_C93_n808, Z => mult_28_C93_n740);
   mult_28_C93_U618 : EXNOR2D1 port map( A1 => mult_28_C93_n19, A2 => 
                           mult_28_C93_n807, Z => mult_28_C93_n739);
   mult_28_C93_U617 : EXNOR2D1 port map( A1 => mult_28_C93_n19, A2 => 
                           mult_28_C93_n806, Z => mult_28_C93_n738);
   mult_28_C93_U616 : EXNOR2D1 port map( A1 => mult_28_C93_n19, A2 => 
                           mult_28_C93_n805, Z => mult_28_C93_n737);
   mult_28_C93_U615 : EXNOR2D1 port map( A1 => mult_28_C93_n19, A2 => 
                           data_in(6), Z => mult_28_C93_n736);
   mult_28_C93_U614 : EXNOR2D1 port map( A1 => mult_28_C93_n19, A2 => 
                           mult_28_C93_n803, Z => mult_28_C93_n735);
   mult_28_C93_U613 : EXNOR2D1 port map( A1 => mult_28_C93_n19, A2 => 
                           mult_28_C93_n802, Z => mult_28_C93_n734);
   mult_28_C93_U612 : EXNOR2D1 port map( A1 => mult_28_C93_n19, A2 => 
                           mult_28_C93_n801, Z => mult_28_C93_n733);
   mult_28_C93_U611 : EXNOR2D1 port map( A1 => mult_28_C93_n19, A2 => 
                           mult_28_C93_n800, Z => mult_28_C93_n732);
   mult_28_C93_U610 : EXNOR2D1 port map( A1 => mult_28_C93_n19, A2 => 
                           mult_28_C93_n799, Z => mult_28_C93_n731);
   mult_28_C93_U609 : EXNOR2D1 port map( A1 => mult_28_C93_n19, A2 => 
                           mult_28_C93_n798, Z => mult_28_C93_n730);
   mult_28_C93_U608 : EXNOR2D1 port map( A1 => mult_28_C93_n19, A2 => 
                           mult_28_C93_n797, Z => mult_28_C93_n729);
   mult_28_C93_U607 : EXNOR2D1 port map( A1 => mult_28_C93_n19, A2 => 
                           mult_28_C93_n796, Z => mult_28_C93_n728);
   mult_28_C93_U606 : EXNOR2D1 port map( A1 => mult_28_C93_n19, A2 => 
                           mult_28_C93_n795, Z => mult_28_C93_n727);
   mult_28_C93_U605 : NOR2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C93_n21, Z => mult_28_C93_n610);
   mult_28_C93_U604 : OAI22D1 port map( A1 => mult_28_C93_n21, A2 => 
                           mult_28_C93_n741, B1 => mult_28_C93_n23, B2 => 
                           mult_28_C93_n742, Z => mult_28_C93_n609);
   mult_28_C93_U603 : OAI22D1 port map( A1 => mult_28_C93_n21, A2 => 
                           mult_28_C93_n740, B1 => mult_28_C93_n23, B2 => 
                           mult_28_C93_n741, Z => mult_28_C93_n608);
   mult_28_C93_U602 : OAI22D1 port map( A1 => mult_28_C93_n21, A2 => 
                           mult_28_C93_n739, B1 => mult_28_C93_n23, B2 => 
                           mult_28_C93_n740, Z => mult_28_C93_n607);
   mult_28_C93_U601 : OAI22D1 port map( A1 => mult_28_C93_n21, A2 => 
                           mult_28_C93_n738, B1 => mult_28_C93_n23, B2 => 
                           mult_28_C93_n739, Z => mult_28_C93_n606);
   mult_28_C93_U600 : OAI22D1 port map( A1 => mult_28_C93_n21, A2 => 
                           mult_28_C93_n737, B1 => mult_28_C93_n23, B2 => 
                           mult_28_C93_n738, Z => mult_28_C93_n605);
   mult_28_C93_U599 : OAI22D1 port map( A1 => mult_28_C93_n21, A2 => 
                           mult_28_C93_n736, B1 => mult_28_C93_n23, B2 => 
                           mult_28_C93_n737, Z => mult_28_C93_n604);
   mult_28_C93_U598 : OAI22D1 port map( A1 => mult_28_C93_n21, A2 => 
                           mult_28_C93_n735, B1 => mult_28_C93_n23, B2 => 
                           mult_28_C93_n736, Z => mult_28_C93_n603);
   mult_28_C93_U597 : OAI22D1 port map( A1 => mult_28_C93_n21, A2 => 
                           mult_28_C93_n734, B1 => mult_28_C93_n23, B2 => 
                           mult_28_C93_n735, Z => mult_28_C93_n602);
   mult_28_C93_U596 : OAI22D1 port map( A1 => mult_28_C93_n22, A2 => 
                           mult_28_C93_n733, B1 => mult_28_C93_n24, B2 => 
                           mult_28_C93_n734, Z => mult_28_C93_n601);
   mult_28_C93_U595 : OAI22D1 port map( A1 => mult_28_C93_n22, A2 => 
                           mult_28_C93_n732, B1 => mult_28_C93_n24, B2 => 
                           mult_28_C93_n733, Z => mult_28_C93_n600);
   mult_28_C93_U594 : OAI22D1 port map( A1 => mult_28_C93_n22, A2 => 
                           mult_28_C93_n731, B1 => mult_28_C93_n24, B2 => 
                           mult_28_C93_n732, Z => mult_28_C93_n599);
   mult_28_C93_U593 : OAI22D1 port map( A1 => mult_28_C93_n22, A2 => 
                           mult_28_C93_n730, B1 => mult_28_C93_n24, B2 => 
                           mult_28_C93_n731, Z => mult_28_C93_n598);
   mult_28_C93_U592 : OAI22D1 port map( A1 => mult_28_C93_n22, A2 => 
                           mult_28_C93_n729, B1 => mult_28_C93_n24, B2 => 
                           mult_28_C93_n730, Z => mult_28_C93_n597);
   mult_28_C93_U591 : OAI22D1 port map( A1 => mult_28_C93_n22, A2 => 
                           mult_28_C93_n728, B1 => mult_28_C93_n24, B2 => 
                           mult_28_C93_n729, Z => mult_28_C93_n596);
   mult_28_C93_U590 : OAI22D1 port map( A1 => mult_28_C93_n22, A2 => 
                           mult_28_C93_n727, B1 => mult_28_C93_n24, B2 => 
                           mult_28_C93_n728, Z => mult_28_C93_n361);
   mult_28_C93_U588 : OAI22D1 port map( A1 => mult_28_C93_n22, A2 => 
                           mult_28_C93_n743, B1 => mult_28_C93_n24, B2 => 
                           mult_28_C93_n839, Z => mult_28_C93_n527);
   mult_28_C93_U587 : NAN2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C93_n25, Z => mult_28_C93_n726);
   mult_28_C93_U586 : EXNOR2D1 port map( A1 => mult_28_C93_n25, A2 => 
                           data_in(0), Z => mult_28_C93_n725);
   mult_28_C93_U585 : EXNOR2D1 port map( A1 => mult_28_C93_n25, A2 => 
                           mult_28_C93_n809, Z => mult_28_C93_n724);
   mult_28_C93_U584 : EXNOR2D1 port map( A1 => mult_28_C93_n25, A2 => 
                           mult_28_C93_n808, Z => mult_28_C93_n723);
   mult_28_C93_U583 : EXNOR2D1 port map( A1 => mult_28_C93_n25, A2 => 
                           mult_28_C93_n807, Z => mult_28_C93_n722);
   mult_28_C93_U582 : EXNOR2D1 port map( A1 => mult_28_C93_n25, A2 => 
                           mult_28_C93_n806, Z => mult_28_C93_n721);
   mult_28_C93_U581 : EXNOR2D1 port map( A1 => mult_28_C93_n25, A2 => 
                           mult_28_C93_n805, Z => mult_28_C93_n720);
   mult_28_C93_U580 : EXNOR2D1 port map( A1 => mult_28_C93_n25, A2 => 
                           data_in(6), Z => mult_28_C93_n719);
   mult_28_C93_U579 : EXNOR2D1 port map( A1 => mult_28_C93_n25, A2 => 
                           mult_28_C93_n803, Z => mult_28_C93_n718);
   mult_28_C93_U578 : EXNOR2D1 port map( A1 => mult_28_C93_n25, A2 => 
                           mult_28_C93_n802, Z => mult_28_C93_n717);
   mult_28_C93_U577 : EXNOR2D1 port map( A1 => mult_28_C93_n25, A2 => 
                           mult_28_C93_n801, Z => mult_28_C93_n716);
   mult_28_C93_U576 : EXNOR2D1 port map( A1 => mult_28_C93_n25, A2 => 
                           mult_28_C93_n800, Z => mult_28_C93_n715);
   mult_28_C93_U575 : EXNOR2D1 port map( A1 => mult_28_C93_n25, A2 => 
                           mult_28_C93_n799, Z => mult_28_C93_n714);
   mult_28_C93_U574 : EXNOR2D1 port map( A1 => mult_28_C93_n25, A2 => 
                           mult_28_C93_n798, Z => mult_28_C93_n713);
   mult_28_C93_U573 : EXNOR2D1 port map( A1 => mult_28_C93_n25, A2 => 
                           mult_28_C93_n797, Z => mult_28_C93_n712);
   mult_28_C93_U572 : EXNOR2D1 port map( A1 => mult_28_C93_n25, A2 => 
                           mult_28_C93_n796, Z => mult_28_C93_n711);
   mult_28_C93_U571 : EXNOR2D1 port map( A1 => mult_28_C93_n25, A2 => 
                           mult_28_C93_n795, Z => mult_28_C93_n710);
   mult_28_C93_U570 : NOR2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C93_n27, Z => mult_28_C93_n594);
   mult_28_C93_U569 : OAI22D1 port map( A1 => mult_28_C93_n27, A2 => 
                           mult_28_C93_n724, B1 => mult_28_C93_n29, B2 => 
                           mult_28_C93_n725, Z => mult_28_C93_n593);
   mult_28_C93_U568 : OAI22D1 port map( A1 => mult_28_C93_n27, A2 => 
                           mult_28_C93_n723, B1 => mult_28_C93_n29, B2 => 
                           mult_28_C93_n724, Z => mult_28_C93_n592);
   mult_28_C93_U567 : OAI22D1 port map( A1 => mult_28_C93_n27, A2 => 
                           mult_28_C93_n722, B1 => mult_28_C93_n29, B2 => 
                           mult_28_C93_n723, Z => mult_28_C93_n591);
   mult_28_C93_U566 : OAI22D1 port map( A1 => mult_28_C93_n27, A2 => 
                           mult_28_C93_n721, B1 => mult_28_C93_n29, B2 => 
                           mult_28_C93_n722, Z => mult_28_C93_n590);
   mult_28_C93_U565 : OAI22D1 port map( A1 => mult_28_C93_n27, A2 => 
                           mult_28_C93_n720, B1 => mult_28_C93_n29, B2 => 
                           mult_28_C93_n721, Z => mult_28_C93_n589);
   mult_28_C93_U564 : OAI22D1 port map( A1 => mult_28_C93_n27, A2 => 
                           mult_28_C93_n719, B1 => mult_28_C93_n29, B2 => 
                           mult_28_C93_n720, Z => mult_28_C93_n588);
   mult_28_C93_U563 : OAI22D1 port map( A1 => mult_28_C93_n27, A2 => 
                           mult_28_C93_n718, B1 => mult_28_C93_n29, B2 => 
                           mult_28_C93_n719, Z => mult_28_C93_n587);
   mult_28_C93_U562 : OAI22D1 port map( A1 => mult_28_C93_n27, A2 => 
                           mult_28_C93_n717, B1 => mult_28_C93_n29, B2 => 
                           mult_28_C93_n718, Z => mult_28_C93_n586);
   mult_28_C93_U561 : OAI22D1 port map( A1 => mult_28_C93_n28, A2 => 
                           mult_28_C93_n716, B1 => mult_28_C93_n30, B2 => 
                           mult_28_C93_n717, Z => mult_28_C93_n585);
   mult_28_C93_U560 : OAI22D1 port map( A1 => mult_28_C93_n28, A2 => 
                           mult_28_C93_n715, B1 => mult_28_C93_n30, B2 => 
                           mult_28_C93_n716, Z => mult_28_C93_n584);
   mult_28_C93_U559 : OAI22D1 port map( A1 => mult_28_C93_n28, A2 => 
                           mult_28_C93_n714, B1 => mult_28_C93_n30, B2 => 
                           mult_28_C93_n715, Z => mult_28_C93_n583);
   mult_28_C93_U558 : OAI22D1 port map( A1 => mult_28_C93_n28, A2 => 
                           mult_28_C93_n713, B1 => mult_28_C93_n30, B2 => 
                           mult_28_C93_n714, Z => mult_28_C93_n582);
   mult_28_C93_U557 : OAI22D1 port map( A1 => mult_28_C93_n28, A2 => 
                           mult_28_C93_n712, B1 => mult_28_C93_n30, B2 => 
                           mult_28_C93_n713, Z => mult_28_C93_n581);
   mult_28_C93_U556 : OAI22D1 port map( A1 => mult_28_C93_n28, A2 => 
                           mult_28_C93_n711, B1 => mult_28_C93_n30, B2 => 
                           mult_28_C93_n712, Z => mult_28_C93_n580);
   mult_28_C93_U555 : OAI22D1 port map( A1 => mult_28_C93_n28, A2 => 
                           mult_28_C93_n710, B1 => mult_28_C93_n30, B2 => 
                           mult_28_C93_n711, Z => mult_28_C93_n343);
   mult_28_C93_U553 : OAI22D1 port map( A1 => mult_28_C93_n28, A2 => 
                           mult_28_C93_n726, B1 => mult_28_C93_n30, B2 => 
                           mult_28_C93_n838, Z => mult_28_C93_n526);
   mult_28_C93_U552 : NAN2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C93_n31, Z => mult_28_C93_n709);
   mult_28_C93_U551 : EXNOR2D1 port map( A1 => mult_28_C93_n31, A2 => 
                           data_in(0), Z => mult_28_C93_n708);
   mult_28_C93_U550 : EXNOR2D1 port map( A1 => mult_28_C93_n31, A2 => 
                           mult_28_C93_n809, Z => mult_28_C93_n707);
   mult_28_C93_U549 : EXNOR2D1 port map( A1 => mult_28_C93_n31, A2 => 
                           mult_28_C93_n808, Z => mult_28_C93_n706);
   mult_28_C93_U548 : EXNOR2D1 port map( A1 => mult_28_C93_n31, A2 => 
                           mult_28_C93_n807, Z => mult_28_C93_n705);
   mult_28_C93_U547 : EXNOR2D1 port map( A1 => mult_28_C93_n31, A2 => 
                           mult_28_C93_n806, Z => mult_28_C93_n704);
   mult_28_C93_U546 : EXNOR2D1 port map( A1 => mult_28_C93_n31, A2 => 
                           mult_28_C93_n805, Z => mult_28_C93_n703);
   mult_28_C93_U545 : EXNOR2D1 port map( A1 => mult_28_C93_n31, A2 => 
                           data_in(6), Z => mult_28_C93_n702);
   mult_28_C93_U544 : EXNOR2D1 port map( A1 => mult_28_C93_n31, A2 => 
                           mult_28_C93_n803, Z => mult_28_C93_n701);
   mult_28_C93_U543 : EXNOR2D1 port map( A1 => mult_28_C93_n31, A2 => 
                           mult_28_C93_n802, Z => mult_28_C93_n700);
   mult_28_C93_U542 : EXNOR2D1 port map( A1 => mult_28_C93_n31, A2 => 
                           mult_28_C93_n801, Z => mult_28_C93_n699);
   mult_28_C93_U541 : EXNOR2D1 port map( A1 => mult_28_C93_n31, A2 => 
                           mult_28_C93_n800, Z => mult_28_C93_n698);
   mult_28_C93_U540 : EXNOR2D1 port map( A1 => mult_28_C93_n31, A2 => 
                           mult_28_C93_n799, Z => mult_28_C93_n697);
   mult_28_C93_U539 : EXNOR2D1 port map( A1 => mult_28_C93_n31, A2 => 
                           mult_28_C93_n798, Z => mult_28_C93_n696);
   mult_28_C93_U538 : EXNOR2D1 port map( A1 => mult_28_C93_n31, A2 => 
                           mult_28_C93_n797, Z => mult_28_C93_n695);
   mult_28_C93_U537 : EXNOR2D1 port map( A1 => mult_28_C93_n31, A2 => 
                           mult_28_C93_n796, Z => mult_28_C93_n694);
   mult_28_C93_U536 : EXNOR2D1 port map( A1 => mult_28_C93_n31, A2 => 
                           mult_28_C93_n795, Z => mult_28_C93_n693);
   mult_28_C93_U535 : NOR2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C93_n33, Z => mult_28_C93_n578);
   mult_28_C93_U534 : OAI22D1 port map( A1 => mult_28_C93_n33, A2 => 
                           mult_28_C93_n707, B1 => mult_28_C93_n35, B2 => 
                           mult_28_C93_n708, Z => mult_28_C93_n577);
   mult_28_C93_U533 : OAI22D1 port map( A1 => mult_28_C93_n33, A2 => 
                           mult_28_C93_n706, B1 => mult_28_C93_n35, B2 => 
                           mult_28_C93_n707, Z => mult_28_C93_n576);
   mult_28_C93_U532 : OAI22D1 port map( A1 => mult_28_C93_n33, A2 => 
                           mult_28_C93_n705, B1 => mult_28_C93_n35, B2 => 
                           mult_28_C93_n706, Z => mult_28_C93_n575);
   mult_28_C93_U531 : OAI22D1 port map( A1 => mult_28_C93_n33, A2 => 
                           mult_28_C93_n704, B1 => mult_28_C93_n35, B2 => 
                           mult_28_C93_n705, Z => mult_28_C93_n574);
   mult_28_C93_U530 : OAI22D1 port map( A1 => mult_28_C93_n33, A2 => 
                           mult_28_C93_n703, B1 => mult_28_C93_n35, B2 => 
                           mult_28_C93_n704, Z => mult_28_C93_n573);
   mult_28_C93_U529 : OAI22D1 port map( A1 => mult_28_C93_n33, A2 => 
                           mult_28_C93_n702, B1 => mult_28_C93_n35, B2 => 
                           mult_28_C93_n703, Z => mult_28_C93_n572);
   mult_28_C93_U528 : OAI22D1 port map( A1 => mult_28_C93_n33, A2 => 
                           mult_28_C93_n701, B1 => mult_28_C93_n35, B2 => 
                           mult_28_C93_n702, Z => mult_28_C93_n571);
   mult_28_C93_U527 : OAI22D1 port map( A1 => mult_28_C93_n33, A2 => 
                           mult_28_C93_n700, B1 => mult_28_C93_n35, B2 => 
                           mult_28_C93_n701, Z => mult_28_C93_n570);
   mult_28_C93_U526 : OAI22D1 port map( A1 => mult_28_C93_n34, A2 => 
                           mult_28_C93_n699, B1 => mult_28_C93_n36, B2 => 
                           mult_28_C93_n700, Z => mult_28_C93_n569);
   mult_28_C93_U525 : OAI22D1 port map( A1 => mult_28_C93_n34, A2 => 
                           mult_28_C93_n698, B1 => mult_28_C93_n36, B2 => 
                           mult_28_C93_n699, Z => mult_28_C93_n568);
   mult_28_C93_U524 : OAI22D1 port map( A1 => mult_28_C93_n34, A2 => 
                           mult_28_C93_n697, B1 => mult_28_C93_n36, B2 => 
                           mult_28_C93_n698, Z => mult_28_C93_n567);
   mult_28_C93_U523 : OAI22D1 port map( A1 => mult_28_C93_n34, A2 => 
                           mult_28_C93_n696, B1 => mult_28_C93_n36, B2 => 
                           mult_28_C93_n697, Z => mult_28_C93_n566);
   mult_28_C93_U522 : OAI22D1 port map( A1 => mult_28_C93_n34, A2 => 
                           mult_28_C93_n695, B1 => mult_28_C93_n36, B2 => 
                           mult_28_C93_n696, Z => mult_28_C93_n565);
   mult_28_C93_U521 : OAI22D1 port map( A1 => mult_28_C93_n34, A2 => 
                           mult_28_C93_n694, B1 => mult_28_C93_n36, B2 => 
                           mult_28_C93_n695, Z => mult_28_C93_n564);
   mult_28_C93_U520 : OAI22D1 port map( A1 => mult_28_C93_n34, A2 => 
                           mult_28_C93_n693, B1 => mult_28_C93_n36, B2 => 
                           mult_28_C93_n694, Z => mult_28_C93_n329);
   mult_28_C93_U518 : OAI22D1 port map( A1 => mult_28_C93_n34, A2 => 
                           mult_28_C93_n709, B1 => mult_28_C93_n36, B2 => 
                           mult_28_C93_n837, Z => mult_28_C93_n525);
   mult_28_C93_U517 : NAN2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C93_n37, Z => mult_28_C93_n692);
   mult_28_C93_U516 : EXNOR2D1 port map( A1 => mult_28_C93_n37, A2 => 
                           data_in(0), Z => mult_28_C93_n691);
   mult_28_C93_U515 : EXNOR2D1 port map( A1 => mult_28_C93_n37, A2 => 
                           mult_28_C93_n809, Z => mult_28_C93_n690);
   mult_28_C93_U514 : EXNOR2D1 port map( A1 => mult_28_C93_n37, A2 => 
                           mult_28_C93_n808, Z => mult_28_C93_n689);
   mult_28_C93_U513 : EXNOR2D1 port map( A1 => mult_28_C93_n37, A2 => 
                           mult_28_C93_n807, Z => mult_28_C93_n688);
   mult_28_C93_U512 : EXNOR2D1 port map( A1 => mult_28_C93_n37, A2 => 
                           mult_28_C93_n806, Z => mult_28_C93_n687);
   mult_28_C93_U511 : EXNOR2D1 port map( A1 => mult_28_C93_n37, A2 => 
                           mult_28_C93_n805, Z => mult_28_C93_n686);
   mult_28_C93_U510 : EXNOR2D1 port map( A1 => mult_28_C93_n37, A2 => 
                           data_in(6), Z => mult_28_C93_n685);
   mult_28_C93_U509 : EXNOR2D1 port map( A1 => mult_28_C93_n37, A2 => 
                           mult_28_C93_n803, Z => mult_28_C93_n684);
   mult_28_C93_U508 : EXNOR2D1 port map( A1 => mult_28_C93_n37, A2 => 
                           mult_28_C93_n802, Z => mult_28_C93_n683);
   mult_28_C93_U507 : EXNOR2D1 port map( A1 => mult_28_C93_n37, A2 => 
                           mult_28_C93_n801, Z => mult_28_C93_n682);
   mult_28_C93_U506 : EXNOR2D1 port map( A1 => mult_28_C93_n37, A2 => 
                           mult_28_C93_n800, Z => mult_28_C93_n681);
   mult_28_C93_U505 : EXNOR2D1 port map( A1 => mult_28_C93_n37, A2 => 
                           mult_28_C93_n799, Z => mult_28_C93_n680);
   mult_28_C93_U504 : EXNOR2D1 port map( A1 => mult_28_C93_n37, A2 => 
                           mult_28_C93_n798, Z => mult_28_C93_n679);
   mult_28_C93_U503 : EXNOR2D1 port map( A1 => mult_28_C93_n37, A2 => 
                           mult_28_C93_n797, Z => mult_28_C93_n678);
   mult_28_C93_U502 : EXNOR2D1 port map( A1 => mult_28_C93_n37, A2 => 
                           mult_28_C93_n796, Z => mult_28_C93_n677);
   mult_28_C93_U501 : EXNOR2D1 port map( A1 => mult_28_C93_n37, A2 => 
                           mult_28_C93_n795, Z => mult_28_C93_n676);
   mult_28_C93_U500 : NOR2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C93_n39, Z => mult_28_C93_n562);
   mult_28_C93_U499 : OAI22D1 port map( A1 => mult_28_C93_n39, A2 => 
                           mult_28_C93_n690, B1 => mult_28_C93_n41, B2 => 
                           mult_28_C93_n691, Z => mult_28_C93_n561);
   mult_28_C93_U498 : OAI22D1 port map( A1 => mult_28_C93_n39, A2 => 
                           mult_28_C93_n689, B1 => mult_28_C93_n41, B2 => 
                           mult_28_C93_n690, Z => mult_28_C93_n560);
   mult_28_C93_U497 : OAI22D1 port map( A1 => mult_28_C93_n39, A2 => 
                           mult_28_C93_n688, B1 => mult_28_C93_n41, B2 => 
                           mult_28_C93_n689, Z => mult_28_C93_n559);
   mult_28_C93_U496 : OAI22D1 port map( A1 => mult_28_C93_n39, A2 => 
                           mult_28_C93_n687, B1 => mult_28_C93_n41, B2 => 
                           mult_28_C93_n688, Z => mult_28_C93_n558);
   mult_28_C93_U495 : OAI22D1 port map( A1 => mult_28_C93_n39, A2 => 
                           mult_28_C93_n686, B1 => mult_28_C93_n41, B2 => 
                           mult_28_C93_n687, Z => mult_28_C93_n557);
   mult_28_C93_U494 : OAI22D1 port map( A1 => mult_28_C93_n39, A2 => 
                           mult_28_C93_n685, B1 => mult_28_C93_n41, B2 => 
                           mult_28_C93_n686, Z => mult_28_C93_n556);
   mult_28_C93_U493 : OAI22D1 port map( A1 => mult_28_C93_n39, A2 => 
                           mult_28_C93_n684, B1 => mult_28_C93_n41, B2 => 
                           mult_28_C93_n685, Z => mult_28_C93_n555);
   mult_28_C93_U492 : OAI22D1 port map( A1 => mult_28_C93_n39, A2 => 
                           mult_28_C93_n683, B1 => mult_28_C93_n41, B2 => 
                           mult_28_C93_n684, Z => mult_28_C93_n554);
   mult_28_C93_U491 : OAI22D1 port map( A1 => mult_28_C93_n40, A2 => 
                           mult_28_C93_n682, B1 => mult_28_C93_n42, B2 => 
                           mult_28_C93_n683, Z => mult_28_C93_n553);
   mult_28_C93_U490 : OAI22D1 port map( A1 => mult_28_C93_n40, A2 => 
                           mult_28_C93_n681, B1 => mult_28_C93_n42, B2 => 
                           mult_28_C93_n682, Z => mult_28_C93_n552);
   mult_28_C93_U489 : OAI22D1 port map( A1 => mult_28_C93_n40, A2 => 
                           mult_28_C93_n680, B1 => mult_28_C93_n42, B2 => 
                           mult_28_C93_n681, Z => mult_28_C93_n551);
   mult_28_C93_U488 : OAI22D1 port map( A1 => mult_28_C93_n40, A2 => 
                           mult_28_C93_n679, B1 => mult_28_C93_n42, B2 => 
                           mult_28_C93_n680, Z => mult_28_C93_n550);
   mult_28_C93_U487 : OAI22D1 port map( A1 => mult_28_C93_n40, A2 => 
                           mult_28_C93_n678, B1 => mult_28_C93_n42, B2 => 
                           mult_28_C93_n679, Z => mult_28_C93_n549);
   mult_28_C93_U486 : OAI22D1 port map( A1 => mult_28_C93_n40, A2 => 
                           mult_28_C93_n677, B1 => mult_28_C93_n42, B2 => 
                           mult_28_C93_n678, Z => mult_28_C93_n548);
   mult_28_C93_U485 : OAI22D1 port map( A1 => mult_28_C93_n40, A2 => 
                           mult_28_C93_n676, B1 => mult_28_C93_n42, B2 => 
                           mult_28_C93_n677, Z => mult_28_C93_n319);
   mult_28_C93_U482 : NAN2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C93_n43, Z => mult_28_C93_n675);
   mult_28_C93_U481 : EXNOR2D1 port map( A1 => mult_28_C93_n43, A2 => 
                           data_in(0), Z => mult_28_C93_n674);
   mult_28_C93_U480 : EXNOR2D1 port map( A1 => mult_28_C93_n43, A2 => 
                           mult_28_C93_n809, Z => mult_28_C93_n673);
   mult_28_C93_U479 : EXNOR2D1 port map( A1 => mult_28_C93_n43, A2 => 
                           mult_28_C93_n808, Z => mult_28_C93_n672);
   mult_28_C93_U478 : EXNOR2D1 port map( A1 => mult_28_C93_n43, A2 => 
                           mult_28_C93_n807, Z => mult_28_C93_n671);
   mult_28_C93_U477 : EXNOR2D1 port map( A1 => mult_28_C93_n43, A2 => 
                           mult_28_C93_n806, Z => mult_28_C93_n670);
   mult_28_C93_U476 : EXNOR2D1 port map( A1 => mult_28_C93_n43, A2 => 
                           mult_28_C93_n805, Z => mult_28_C93_n669);
   mult_28_C93_U475 : EXNOR2D1 port map( A1 => mult_28_C93_n43, A2 => 
                           data_in(6), Z => mult_28_C93_n668);
   mult_28_C93_U474 : EXNOR2D1 port map( A1 => mult_28_C93_n43, A2 => 
                           mult_28_C93_n803, Z => mult_28_C93_n667);
   mult_28_C93_U473 : EXNOR2D1 port map( A1 => mult_28_C93_n43, A2 => 
                           mult_28_C93_n802, Z => mult_28_C93_n666);
   mult_28_C93_U472 : EXNOR2D1 port map( A1 => mult_28_C93_n43, A2 => 
                           mult_28_C93_n801, Z => mult_28_C93_n665);
   mult_28_C93_U471 : EXNOR2D1 port map( A1 => mult_28_C93_n43, A2 => 
                           mult_28_C93_n800, Z => mult_28_C93_n664);
   mult_28_C93_U470 : EXNOR2D1 port map( A1 => mult_28_C93_n43, A2 => 
                           mult_28_C93_n799, Z => mult_28_C93_n663);
   mult_28_C93_U469 : EXNOR2D1 port map( A1 => mult_28_C93_n43, A2 => 
                           mult_28_C93_n798, Z => mult_28_C93_n662);
   mult_28_C93_U468 : EXNOR2D1 port map( A1 => mult_28_C93_n43, A2 => 
                           mult_28_C93_n797, Z => mult_28_C93_n661);
   mult_28_C93_U467 : EXNOR2D1 port map( A1 => mult_28_C93_n43, A2 => 
                           mult_28_C93_n796, Z => mult_28_C93_n660);
   mult_28_C93_U466 : EXNOR2D1 port map( A1 => mult_28_C93_n43, A2 => 
                           mult_28_C93_n795, Z => mult_28_C93_n659);
   mult_28_C93_U465 : NOR2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C93_n45, Z => mult_28_C93_n546);
   mult_28_C93_U464 : OAI22D1 port map( A1 => mult_28_C93_n45, A2 => 
                           mult_28_C93_n673, B1 => mult_28_C93_n47, B2 => 
                           mult_28_C93_n674, Z => mult_28_C93_n545);
   mult_28_C93_U463 : OAI22D1 port map( A1 => mult_28_C93_n45, A2 => 
                           mult_28_C93_n672, B1 => mult_28_C93_n47, B2 => 
                           mult_28_C93_n673, Z => mult_28_C93_n544);
   mult_28_C93_U462 : OAI22D1 port map( A1 => mult_28_C93_n45, A2 => 
                           mult_28_C93_n671, B1 => mult_28_C93_n47, B2 => 
                           mult_28_C93_n672, Z => mult_28_C93_n543);
   mult_28_C93_U461 : OAI22D1 port map( A1 => mult_28_C93_n45, A2 => 
                           mult_28_C93_n670, B1 => mult_28_C93_n47, B2 => 
                           mult_28_C93_n671, Z => mult_28_C93_n542);
   mult_28_C93_U460 : OAI22D1 port map( A1 => mult_28_C93_n45, A2 => 
                           mult_28_C93_n669, B1 => mult_28_C93_n47, B2 => 
                           mult_28_C93_n670, Z => mult_28_C93_n541);
   mult_28_C93_U459 : OAI22D1 port map( A1 => mult_28_C93_n45, A2 => 
                           mult_28_C93_n668, B1 => mult_28_C93_n47, B2 => 
                           mult_28_C93_n669, Z => mult_28_C93_n540);
   mult_28_C93_U458 : OAI22D1 port map( A1 => mult_28_C93_n45, A2 => 
                           mult_28_C93_n667, B1 => mult_28_C93_n47, B2 => 
                           mult_28_C93_n668, Z => mult_28_C93_n539);
   mult_28_C93_U457 : OAI22D1 port map( A1 => mult_28_C93_n45, A2 => 
                           mult_28_C93_n666, B1 => mult_28_C93_n47, B2 => 
                           mult_28_C93_n667, Z => mult_28_C93_n538);
   mult_28_C93_U456 : OAI22D1 port map( A1 => mult_28_C93_n46, A2 => 
                           mult_28_C93_n665, B1 => mult_28_C93_n48, B2 => 
                           mult_28_C93_n666, Z => mult_28_C93_n537);
   mult_28_C93_U455 : OAI22D1 port map( A1 => mult_28_C93_n46, A2 => 
                           mult_28_C93_n664, B1 => mult_28_C93_n48, B2 => 
                           mult_28_C93_n665, Z => mult_28_C93_n536);
   mult_28_C93_U454 : OAI22D1 port map( A1 => mult_28_C93_n46, A2 => 
                           mult_28_C93_n663, B1 => mult_28_C93_n48, B2 => 
                           mult_28_C93_n664, Z => mult_28_C93_n535);
   mult_28_C93_U453 : OAI22D1 port map( A1 => mult_28_C93_n46, A2 => 
                           mult_28_C93_n662, B1 => mult_28_C93_n48, B2 => 
                           mult_28_C93_n663, Z => mult_28_C93_n534);
   mult_28_C93_U452 : OAI22D1 port map( A1 => mult_28_C93_n46, A2 => 
                           mult_28_C93_n661, B1 => mult_28_C93_n48, B2 => 
                           mult_28_C93_n662, Z => mult_28_C93_n533);
   mult_28_C93_U451 : OAI22D1 port map( A1 => mult_28_C93_n46, A2 => 
                           mult_28_C93_n660, B1 => mult_28_C93_n48, B2 => 
                           mult_28_C93_n661, Z => mult_28_C93_n532);
   mult_28_C93_U447 : ADFULD1 port map( A => mult_28_C93_n655, B => 
                           mult_28_C93_n626, CI => mult_28_C93_n640, CO => 
                           mult_28_C93_n519, S => mult_28_C93_n520);
   mult_28_C93_U445 : ADFULD1 port map( A => mult_28_C93_n625, B => 
                           mult_28_C93_n639, CI => mult_28_C93_n518, CO => 
                           mult_28_C93_n515, S => mult_28_C93_n516);
   mult_28_C93_U444 : ADFULD1 port map( A => mult_28_C93_n653, B => 
                           mult_28_C93_n610, CI => mult_28_C93_n638, CO => 
                           mult_28_C93_n513, S => mult_28_C93_n514);
   mult_28_C93_U443 : ADFULD1 port map( A => mult_28_C93_n517, B => 
                           mult_28_C93_n624, CI => mult_28_C93_n514, CO => 
                           mult_28_C93_n511, S => mult_28_C93_n512);
   mult_28_C93_U441 : ADFULD1 port map( A => mult_28_C93_n609, B => 
                           mult_28_C93_n637, CI => mult_28_C93_n623, CO => 
                           mult_28_C93_n507, S => mult_28_C93_n508);
   mult_28_C93_U440 : ADFULD1 port map( A => mult_28_C93_n513, B => 
                           mult_28_C93_n510, CI => mult_28_C93_n508, CO => 
                           mult_28_C93_n505, S => mult_28_C93_n506);
   mult_28_C93_U439 : ADFULD1 port map( A => mult_28_C93_n651, B => 
                           mult_28_C93_n594, CI => mult_28_C93_n636, CO => 
                           mult_28_C93_n503, S => mult_28_C93_n504);
   mult_28_C93_U438 : ADFULD1 port map( A => mult_28_C93_n608, B => 
                           mult_28_C93_n622, CI => mult_28_C93_n509, CO => 
                           mult_28_C93_n501, S => mult_28_C93_n502);
   mult_28_C93_U437 : ADFULD1 port map( A => mult_28_C93_n504, B => 
                           mult_28_C93_n507, CI => mult_28_C93_n502, CO => 
                           mult_28_C93_n499, S => mult_28_C93_n500);
   mult_28_C93_U435 : ADFULD1 port map( A => mult_28_C93_n593, B => 
                           mult_28_C93_n607, CI => mult_28_C93_n621, CO => 
                           mult_28_C93_n495, S => mult_28_C93_n496);
   mult_28_C93_U434 : ADFULD1 port map( A => mult_28_C93_n498, B => 
                           mult_28_C93_n635, CI => mult_28_C93_n503, CO => 
                           mult_28_C93_n493, S => mult_28_C93_n494);
   mult_28_C93_U433 : ADFULD1 port map( A => mult_28_C93_n496, B => 
                           mult_28_C93_n501, CI => mult_28_C93_n494, CO => 
                           mult_28_C93_n491, S => mult_28_C93_n492);
   mult_28_C93_U432 : ADFULD1 port map( A => mult_28_C93_n649, B => 
                           mult_28_C93_n578, CI => mult_28_C93_n634, CO => 
                           mult_28_C93_n489, S => mult_28_C93_n490);
   mult_28_C93_U431 : ADFULD1 port map( A => mult_28_C93_n592, B => 
                           mult_28_C93_n620, CI => mult_28_C93_n606, CO => 
                           mult_28_C93_n487, S => mult_28_C93_n488);
   mult_28_C93_U430 : ADFULD1 port map( A => mult_28_C93_n495, B => 
                           mult_28_C93_n497, CI => mult_28_C93_n490, CO => 
                           mult_28_C93_n485, S => mult_28_C93_n486);
   mult_28_C93_U429 : ADFULD1 port map( A => mult_28_C93_n493, B => 
                           mult_28_C93_n488, CI => mult_28_C93_n486, CO => 
                           mult_28_C93_n483, S => mult_28_C93_n484);
   mult_28_C93_U427 : ADFULD1 port map( A => mult_28_C93_n577, B => 
                           mult_28_C93_n605, CI => mult_28_C93_n633, CO => 
                           mult_28_C93_n479, S => mult_28_C93_n480);
   mult_28_C93_U426 : ADFULD1 port map( A => mult_28_C93_n591, B => 
                           mult_28_C93_n619, CI => mult_28_C93_n482, CO => 
                           mult_28_C93_n477, S => mult_28_C93_n478);
   mult_28_C93_U425 : ADFULD1 port map( A => mult_28_C93_n487, B => 
                           mult_28_C93_n489, CI => mult_28_C93_n480, CO => 
                           mult_28_C93_n475, S => mult_28_C93_n476);
   mult_28_C93_U424 : ADFULD1 port map( A => mult_28_C93_n485, B => 
                           mult_28_C93_n478, CI => mult_28_C93_n476, CO => 
                           mult_28_C93_n473, S => mult_28_C93_n474);
   mult_28_C93_U423 : ADFULD1 port map( A => mult_28_C93_n647, B => 
                           mult_28_C93_n562, CI => mult_28_C93_n632, CO => 
                           mult_28_C93_n471, S => mult_28_C93_n472);
   mult_28_C93_U422 : ADFULD1 port map( A => mult_28_C93_n576, B => 
                           mult_28_C93_n618, CI => mult_28_C93_n590, CO => 
                           mult_28_C93_n469, S => mult_28_C93_n470);
   mult_28_C93_U421 : ADFULD1 port map( A => mult_28_C93_n481, B => 
                           mult_28_C93_n604, CI => mult_28_C93_n479, CO => 
                           mult_28_C93_n467, S => mult_28_C93_n468);
   mult_28_C93_U420 : ADFULD1 port map( A => mult_28_C93_n470, B => 
                           mult_28_C93_n472, CI => mult_28_C93_n477, CO => 
                           mult_28_C93_n465, S => mult_28_C93_n466);
   mult_28_C93_U419 : ADFULD1 port map( A => mult_28_C93_n468, B => 
                           mult_28_C93_n475, CI => mult_28_C93_n466, CO => 
                           mult_28_C93_n463, S => mult_28_C93_n464);
   mult_28_C93_U418 : ADHALFD1 port map( A => mult_28_C93_n524, B => 
                           mult_28_C93_n646, CO => mult_28_C93_n461, S => 
                           mult_28_C93_n462);
   mult_28_C93_U417 : ADFULD1 port map( A => mult_28_C93_n631, B => 
                           mult_28_C93_n589, CI => mult_28_C93_n617, CO => 
                           mult_28_C93_n459, S => mult_28_C93_n460);
   mult_28_C93_U416 : ADFULD1 port map( A => mult_28_C93_n561, B => 
                           mult_28_C93_n603, CI => mult_28_C93_n575, CO => 
                           mult_28_C93_n457, S => mult_28_C93_n458);
   mult_28_C93_U415 : ADFULD1 port map( A => mult_28_C93_n471, B => 
                           mult_28_C93_n462, CI => mult_28_C93_n469, CO => 
                           mult_28_C93_n455, S => mult_28_C93_n456);
   mult_28_C93_U414 : ADFULD1 port map( A => mult_28_C93_n460, B => 
                           mult_28_C93_n458, CI => mult_28_C93_n467, CO => 
                           mult_28_C93_n453, S => mult_28_C93_n454);
   mult_28_C93_U413 : ADFULD1 port map( A => mult_28_C93_n465, B => 
                           mult_28_C93_n456, CI => mult_28_C93_n454, CO => 
                           mult_28_C93_n451, S => mult_28_C93_n452);
   mult_28_C93_U412 : ADFULD1 port map( A => mult_28_C93_n645, B => 
                           mult_28_C93_n546, CI => mult_28_C93_n630, CO => 
                           mult_28_C93_n449, S => mult_28_C93_n450);
   mult_28_C93_U411 : ADFULD1 port map( A => mult_28_C93_n560, B => 
                           mult_28_C93_n616, CI => mult_28_C93_n574, CO => 
                           mult_28_C93_n447, S => mult_28_C93_n448);
   mult_28_C93_U410 : ADFULD1 port map( A => mult_28_C93_n588, B => 
                           mult_28_C93_n602, CI => mult_28_C93_n461, CO => 
                           mult_28_C93_n445, S => mult_28_C93_n446);
   mult_28_C93_U409 : ADFULD1 port map( A => mult_28_C93_n457, B => 
                           mult_28_C93_n459, CI => mult_28_C93_n450, CO => 
                           mult_28_C93_n443, S => mult_28_C93_n444);
   mult_28_C93_U408 : ADFULD1 port map( A => mult_28_C93_n446, B => 
                           mult_28_C93_n448, CI => mult_28_C93_n455, CO => 
                           mult_28_C93_n441, S => mult_28_C93_n442);
   mult_28_C93_U407 : ADFULD1 port map( A => mult_28_C93_n453, B => 
                           mult_28_C93_n444, CI => mult_28_C93_n442, CO => 
                           mult_28_C93_n439, S => mult_28_C93_n440);
   mult_28_C93_U406 : ADHALFD1 port map( A => mult_28_C93_n523, B => 
                           mult_28_C93_n644, CO => mult_28_C93_n437, S => 
                           mult_28_C93_n438);
   mult_28_C93_U405 : ADFULD1 port map( A => mult_28_C93_n545, B => 
                           mult_28_C93_n587, CI => mult_28_C93_n559, CO => 
                           mult_28_C93_n435, S => mult_28_C93_n436);
   mult_28_C93_U404 : ADFULD1 port map( A => mult_28_C93_n629, B => 
                           mult_28_C93_n573, CI => mult_28_C93_n601, CO => 
                           mult_28_C93_n433, S => mult_28_C93_n434);
   mult_28_C93_U403 : ADFULD1 port map( A => mult_28_C93_n438, B => 
                           mult_28_C93_n615, CI => mult_28_C93_n449, CO => 
                           mult_28_C93_n431, S => mult_28_C93_n432);
   mult_28_C93_U402 : ADFULD1 port map( A => mult_28_C93_n445, B => 
                           mult_28_C93_n447, CI => mult_28_C93_n434, CO => 
                           mult_28_C93_n429, S => mult_28_C93_n430);
   mult_28_C93_U401 : ADFULD1 port map( A => mult_28_C93_n443, B => 
                           mult_28_C93_n436, CI => mult_28_C93_n432, CO => 
                           mult_28_C93_n427, S => mult_28_C93_n428);
   mult_28_C93_U400 : ADFULD1 port map( A => mult_28_C93_n441, B => 
                           mult_28_C93_n430, CI => mult_28_C93_n428, CO => 
                           mult_28_C93_n425, S => mult_28_C93_n426);
   mult_28_C93_U397 : ADFULD1 port map( A => mult_28_C93_n544, B => 
                           mult_28_C93_n586, CI => mult_28_C93_n572, CO => 
                           mult_28_C93_n421, S => mult_28_C93_n422);
   mult_28_C93_U396 : ADFULD1 port map( A => mult_28_C93_n614, B => 
                           mult_28_C93_n628, CI => mult_28_C93_n643, CO => 
                           mult_28_C93_n419, S => mult_28_C93_n420);
   mult_28_C93_U395 : ADFULD1 port map( A => mult_28_C93_n424, B => 
                           mult_28_C93_n437, CI => mult_28_C93_n435, CO => 
                           mult_28_C93_n417, S => mult_28_C93_n418);
   mult_28_C93_U394 : ADFULD1 port map( A => mult_28_C93_n422, B => 
                           mult_28_C93_n433, CI => mult_28_C93_n420, CO => 
                           mult_28_C93_n415, S => mult_28_C93_n416);
   mult_28_C93_U393 : ADFULD1 port map( A => mult_28_C93_n429, B => 
                           mult_28_C93_n431, CI => mult_28_C93_n418, CO => 
                           mult_28_C93_n413, S => mult_28_C93_n414);
   mult_28_C93_U392 : ADFULD1 port map( A => mult_28_C93_n427, B => 
                           mult_28_C93_n416, CI => mult_28_C93_n414, CO => 
                           mult_28_C93_n411, S => mult_28_C93_n412);
   mult_28_C93_U390 : ADFULD1 port map( A => mult_28_C93_n543, B => 
                           mult_28_C93_n571, CI => mult_28_C93_n613, CO => 
                           mult_28_C93_n407, S => mult_28_C93_n408);
   mult_28_C93_U389 : ADFULD1 port map( A => mult_28_C93_n557, B => 
                           mult_28_C93_n599, CI => mult_28_C93_n585, CO => 
                           mult_28_C93_n405, S => mult_28_C93_n406);
   mult_28_C93_U388 : ADFULD1 port map( A => mult_28_C93_n423, B => 
                           mult_28_C93_n410, CI => mult_28_C93_n421, CO => 
                           mult_28_C93_n403, S => mult_28_C93_n404);
   mult_28_C93_U387 : ADFULD1 port map( A => mult_28_C93_n406, B => 
                           mult_28_C93_n419, CI => mult_28_C93_n408, CO => 
                           mult_28_C93_n401, S => mult_28_C93_n402);
   mult_28_C93_U386 : ADFULD1 port map( A => mult_28_C93_n404, B => 
                           mult_28_C93_n417, CI => mult_28_C93_n415, CO => 
                           mult_28_C93_n399, S => mult_28_C93_n400);
   mult_28_C93_U385 : ADFULD1 port map( A => mult_28_C93_n413, B => 
                           mult_28_C93_n402, CI => mult_28_C93_n400, CO => 
                           mult_28_C93_n397, S => mult_28_C93_n398);
   mult_28_C93_U384 : ADFULD1 port map( A => mult_28_C93_n409, B => 
                           mult_28_C93_n542, CI => mult_28_C93_n556, CO => 
                           mult_28_C93_n395, S => mult_28_C93_n396);
   mult_28_C93_U383 : ADFULD1 port map( A => mult_28_C93_n570, B => 
                           mult_28_C93_n598, CI => mult_28_C93_n612, CO => 
                           mult_28_C93_n393, S => mult_28_C93_n394);
   mult_28_C93_U382 : ADFULD1 port map( A => mult_28_C93_n627, B => 
                           mult_28_C93_n584, CI => mult_28_C93_n407, CO => 
                           mult_28_C93_n391, S => mult_28_C93_n392);
   mult_28_C93_U381 : ADFULD1 port map( A => mult_28_C93_n394, B => 
                           mult_28_C93_n405, CI => mult_28_C93_n396, CO => 
                           mult_28_C93_n389, S => mult_28_C93_n390);
   mult_28_C93_U380 : ADFULD1 port map( A => mult_28_C93_n392, B => 
                           mult_28_C93_n403, CI => mult_28_C93_n401, CO => 
                           mult_28_C93_n387, S => mult_28_C93_n388);
   mult_28_C93_U379 : ADFULD1 port map( A => mult_28_C93_n399, B => 
                           mult_28_C93_n390, CI => mult_28_C93_n388, CO => 
                           mult_28_C93_n385, S => mult_28_C93_n386);
   mult_28_C93_U377 : ADFULD1 port map( A => mult_28_C93_n597, B => 
                           mult_28_C93_n569, CI => mult_28_C93_n583, CO => 
                           mult_28_C93_n381, S => mult_28_C93_n382);
   mult_28_C93_U376 : ADFULD1 port map( A => mult_28_C93_n541, B => 
                           mult_28_C93_n555, CI => mult_28_C93_n384, CO => 
                           mult_28_C93_n379, S => mult_28_C93_n380);
   mult_28_C93_U375 : ADFULD1 port map( A => mult_28_C93_n393, B => 
                           mult_28_C93_n395, CI => mult_28_C93_n382, CO => 
                           mult_28_C93_n377, S => mult_28_C93_n378);
   mult_28_C93_U374 : ADFULD1 port map( A => mult_28_C93_n391, B => 
                           mult_28_C93_n380, CI => mult_28_C93_n389, CO => 
                           mult_28_C93_n375, S => mult_28_C93_n376);
   mult_28_C93_U373 : ADFULD1 port map( A => mult_28_C93_n387, B => 
                           mult_28_C93_n378, CI => mult_28_C93_n376, CO => 
                           mult_28_C93_n373, S => mult_28_C93_n374);
   mult_28_C93_U372 : ADFULD1 port map( A => mult_28_C93_n383, B => 
                           mult_28_C93_n540, CI => mult_28_C93_n568, CO => 
                           mult_28_C93_n371, S => mult_28_C93_n372);
   mult_28_C93_U371 : ADFULD1 port map( A => mult_28_C93_n554, B => 
                           mult_28_C93_n582, CI => mult_28_C93_n596, CO => 
                           mult_28_C93_n369, S => mult_28_C93_n370);
   mult_28_C93_U370 : ADFULD1 port map( A => mult_28_C93_n381, B => 
                           mult_28_C93_n611, CI => mult_28_C93_n379, CO => 
                           mult_28_C93_n367, S => mult_28_C93_n368);
   mult_28_C93_U369 : ADFULD1 port map( A => mult_28_C93_n372, B => 
                           mult_28_C93_n370, CI => mult_28_C93_n377, CO => 
                           mult_28_C93_n365, S => mult_28_C93_n366);
   mult_28_C93_U368 : ADFULD1 port map( A => mult_28_C93_n375, B => 
                           mult_28_C93_n368, CI => mult_28_C93_n366, CO => 
                           mult_28_C93_n363, S => mult_28_C93_n364);
   mult_28_C93_U366 : ADFULD1 port map( A => mult_28_C93_n581, B => 
                           mult_28_C93_n553, CI => mult_28_C93_n539, CO => 
                           mult_28_C93_n359, S => mult_28_C93_n360);
   mult_28_C93_U365 : ADFULD1 port map( A => mult_28_C93_n362, B => 
                           mult_28_C93_n567, CI => mult_28_C93_n371, CO => 
                           mult_28_C93_n357, S => mult_28_C93_n358);
   mult_28_C93_U364 : ADFULD1 port map( A => mult_28_C93_n360, B => 
                           mult_28_C93_n369, CI => mult_28_C93_n367, CO => 
                           mult_28_C93_n355, S => mult_28_C93_n356);
   mult_28_C93_U363 : ADFULD1 port map( A => mult_28_C93_n365, B => 
                           mult_28_C93_n358, CI => mult_28_C93_n356, CO => 
                           mult_28_C93_n353, S => mult_28_C93_n354);
   mult_28_C93_U362 : ADFULD1 port map( A => mult_28_C93_n580, B => 
                           mult_28_C93_n538, CI => mult_28_C93_n361, CO => 
                           mult_28_C93_n351, S => mult_28_C93_n352);
   mult_28_C93_U361 : ADFULD1 port map( A => mult_28_C93_n566, B => 
                           mult_28_C93_n552, CI => mult_28_C93_n595, CO => 
                           mult_28_C93_n349, S => mult_28_C93_n350);
   mult_28_C93_U360 : ADFULD1 port map( A => mult_28_C93_n352, B => 
                           mult_28_C93_n359, CI => mult_28_C93_n350, CO => 
                           mult_28_C93_n347, S => mult_28_C93_n348);
   mult_28_C93_U359 : ADFULD1 port map( A => mult_28_C93_n348, B => 
                           mult_28_C93_n357, CI => mult_28_C93_n355, CO => 
                           mult_28_C93_n345, S => mult_28_C93_n346);
   mult_28_C93_U357 : ADFULD1 port map( A => mult_28_C93_n551, B => 
                           mult_28_C93_n537, CI => mult_28_C93_n565, CO => 
                           mult_28_C93_n341, S => mult_28_C93_n342);
   mult_28_C93_U356 : ADFULD1 port map( A => mult_28_C93_n351, B => 
                           mult_28_C93_n344, CI => mult_28_C93_n349, CO => 
                           mult_28_C93_n339, S => mult_28_C93_n340);
   mult_28_C93_U355 : ADFULD1 port map( A => mult_28_C93_n347, B => 
                           mult_28_C93_n342, CI => mult_28_C93_n340, CO => 
                           mult_28_C93_n337, S => mult_28_C93_n338);
   mult_28_C93_U354 : ADFULD1 port map( A => mult_28_C93_n550, B => 
                           mult_28_C93_n536, CI => mult_28_C93_n343, CO => 
                           mult_28_C93_n335, S => mult_28_C93_n336);
   mult_28_C93_U353 : ADFULD1 port map( A => mult_28_C93_n579, B => 
                           mult_28_C93_n564, CI => mult_28_C93_n341, CO => 
                           mult_28_C93_n333, S => mult_28_C93_n334);
   mult_28_C93_U352 : ADFULD1 port map( A => mult_28_C93_n339, B => 
                           mult_28_C93_n336, CI => mult_28_C93_n334, CO => 
                           mult_28_C93_n331, S => mult_28_C93_n332);
   mult_28_C93_U350 : ADFULD1 port map( A => mult_28_C93_n535, B => 
                           mult_28_C93_n549, CI => mult_28_C93_n330, CO => 
                           mult_28_C93_n327, S => mult_28_C93_n328);
   mult_28_C93_U349 : ADFULD1 port map( A => mult_28_C93_n328, B => 
                           mult_28_C93_n335, CI => mult_28_C93_n333, CO => 
                           mult_28_C93_n325, S => mult_28_C93_n326);
   mult_28_C93_U348 : ADFULD1 port map( A => mult_28_C93_n548, B => 
                           mult_28_C93_n329, CI => mult_28_C93_n534, CO => 
                           mult_28_C93_n323, S => mult_28_C93_n324);
   mult_28_C93_U347 : ADFULD1 port map( A => mult_28_C93_n327, B => 
                           mult_28_C93_n563, CI => mult_28_C93_n324, CO => 
                           mult_28_C93_n321, S => mult_28_C93_n322);
   mult_28_C93_U345 : ADFULD1 port map( A => mult_28_C93_n320, B => 
                           mult_28_C93_n533, CI => mult_28_C93_n323, CO => 
                           mult_28_C93_n317, S => mult_28_C93_n318);
   mult_28_C93_U344 : ADFULD1 port map( A => mult_28_C93_n532, B => 
                           mult_28_C93_n319, CI => mult_28_C93_n547, CO => 
                           mult_28_C93_n315, S => mult_28_C93_n316);
   mult_28_C93_U330 : AOI21D1 port map( A1 => mult_28_C93_n935, A2 => 
                           mult_28_C93_n937, B => mult_28_C93_n936, Z => 
                           mult_28_C93_n277);
   mult_28_C93_U324 : OAI21D1 port map( A1 => mult_28_C93_n275, A2 => 
                           mult_28_C93_n277, B => mult_28_C93_n276, Z => 
                           mult_28_C93_n274);
   mult_28_C93_U316 : AOI21D1 port map( A1 => mult_28_C93_n274, A2 => 
                           mult_28_C93_n933, B => mult_28_C93_n934, Z => 
                           mult_28_C93_n269);
   mult_28_C93_U310 : OAI21D1 port map( A1 => mult_28_C93_n267, A2 => 
                           mult_28_C93_n269, B => mult_28_C93_n268, Z => 
                           mult_28_C93_n266);
   mult_28_C93_U302 : AOI21D1 port map( A1 => mult_28_C93_n266, A2 => 
                           mult_28_C93_n931, B => mult_28_C93_n932, Z => 
                           mult_28_C93_n261);
   mult_28_C93_U283 : OAI21D1 port map( A1 => mult_28_C93_n249, A2 => 
                           mult_28_C93_n261, B => mult_28_C93_n250, Z => 
                           mult_28_C93_n248);
   mult_28_C93_U275 : AOI21D1 port map( A1 => mult_28_C93_n248, A2 => 
                           mult_28_C93_n926, B => mult_28_C93_n929, Z => 
                           mult_28_C93_n243);
   mult_28_C93_U258 : AOI21D1 port map( A1 => mult_28_C93_n919, A2 => 
                           mult_28_C93_n921, B => mult_28_C93_n922, Z => 
                           mult_28_C93_n232);
   mult_28_C93_U256 : OAI21D1 port map( A1 => mult_28_C93_n243, A2 => 
                           mult_28_C93_n231, B => mult_28_C93_n232, Z => 
                           mult_28_C93_n230);
   mult_28_C93_U237 : AOI21D1 port map( A1 => mult_28_C93_n923, A2 => 
                           mult_28_C93_n910, B => mult_28_C93_n914, Z => 
                           mult_28_C93_n217);
   mult_28_C93_U232 : NOR2D2 port map( A1 => mult_28_C93_n440, A2 => 
                           mult_28_C93_n451, Z => mult_28_C93_n213);
   mult_28_C93_U225 : EXNOR2D1 port map( A1 => mult_28_C93_n215, A2 => 
                           mult_28_C93_n69, Z => m2_0);
   mult_28_C93_U223 : NOR2D2 port map( A1 => mult_28_C93_n426, A2 => 
                           mult_28_C93_n439, Z => mult_28_C93_n207);
   mult_28_C93_U218 : AOI21D1 port map( A1 => mult_28_C93_n209, A2 => 
                           mult_28_C93_n205, B => mult_28_C93_n206, Z => 
                           mult_28_C93_n204);
   mult_28_C93_U217 : EXNOR2D1 port map( A1 => mult_28_C93_n209, A2 => 
                           mult_28_C93_n68, Z => m2_1);
   mult_28_C93_U215 : NOR2D2 port map( A1 => mult_28_C93_n412, A2 => 
                           mult_28_C93_n425, Z => mult_28_C93_n202);
   mult_28_C93_U212 : OAI21D1 port map( A1 => mult_28_C93_n202, A2 => 
                           mult_28_C93_n208, B => mult_28_C93_n203, Z => 
                           mult_28_C93_n201);
   mult_28_C93_U206 : AOI21D1 port map( A1 => mult_28_C93_n209, A2 => 
                           mult_28_C93_n200, B => mult_28_C93_n197, Z => 
                           mult_28_C93_n195);
   mult_28_C93_U205 : EXOR2D1 port map( A1 => mult_28_C93_n204, A2 => 
                           mult_28_C93_n67, Z => m2_2);
   mult_28_C93_U203 : NOR2D2 port map( A1 => mult_28_C93_n398, A2 => 
                           mult_28_C93_n411, Z => mult_28_C93_n193);
   mult_28_C93_U198 : OAI21D1 port map( A1 => mult_28_C93_n199, A2 => 
                           mult_28_C93_n191, B => mult_28_C93_n194, Z => 
                           mult_28_C93_n190);
   mult_28_C93_U196 : AOI21D1 port map( A1 => mult_28_C93_n189, A2 => 
                           mult_28_C93_n209, B => mult_28_C93_n190, Z => 
                           mult_28_C93_n188);
   mult_28_C93_U195 : EXOR2D1 port map( A1 => mult_28_C93_n195, A2 => 
                           mult_28_C93_n66, Z => m2_3);
   mult_28_C93_U193 : NOR2D2 port map( A1 => mult_28_C93_n386, A2 => 
                           mult_28_C93_n397, Z => mult_28_C93_n186);
   mult_28_C93_U190 : OAI21D1 port map( A1 => mult_28_C93_n186, A2 => 
                           mult_28_C93_n194, B => mult_28_C93_n187, Z => 
                           mult_28_C93_n185);
   mult_28_C93_U188 : AOI21D1 port map( A1 => mult_28_C93_n201, A2 => 
                           mult_28_C93_n184, B => mult_28_C93_n185, Z => 
                           mult_28_C93_n183);
   mult_28_C93_U186 : OAI21D1 port map( A1 => mult_28_C93_n182, A2 => 
                           mult_28_C93_n210, B => mult_28_C93_n183, Z => 
                           mult_28_C93_n181);
   mult_28_C93_U185 : EXOR2D1 port map( A1 => mult_28_C93_n188, A2 => 
                           mult_28_C93_n65, Z => m2_4);
   mult_28_C93_U184 : NAN2D2 port map( A1 => mult_28_C93_n374, A2 => 
                           mult_28_C93_n385, Z => mult_28_C93_n180);
   mult_28_C93_U178 : AOI21D1 port map( A1 => mult_28_C93_n51, A2 => 
                           mult_28_C93_n177, B => mult_28_C93_n178, Z => 
                           mult_28_C93_n176);
   mult_28_C93_U177 : EXNOR2D1 port map( A1 => mult_28_C93_n51, A2 => 
                           mult_28_C93_n64, Z => m2_5);
   mult_28_C93_U175 : NOR2D2 port map( A1 => mult_28_C93_n364, A2 => 
                           mult_28_C93_n373, Z => mult_28_C93_n174);
   mult_28_C93_U172 : OAI21D1 port map( A1 => mult_28_C93_n174, A2 => 
                           mult_28_C93_n180, B => mult_28_C93_n175, Z => 
                           mult_28_C93_n173);
   mult_28_C93_U165 : EXOR2D1 port map( A1 => mult_28_C93_n176, A2 => 
                           mult_28_C93_n63, Z => m2_6);
   mult_28_C93_U163 : NOR2D2 port map( A1 => mult_28_C93_n354, A2 => 
                           mult_28_C93_n363, Z => mult_28_C93_n165);
   mult_28_C93_U154 : AOI21D1 port map( A1 => mult_28_C93_n51, A2 => 
                           mult_28_C93_n159, B => mult_28_C93_n160, Z => 
                           mult_28_C93_n158);
   mult_28_C93_U153 : EXOR2D1 port map( A1 => mult_28_C93_n167, A2 => 
                           mult_28_C93_n62, Z => m2_7);
   mult_28_C93_U144 : AOI21D1 port map( A1 => mult_28_C93_n164, A2 => 
                           mult_28_C93_n152, B => mult_28_C93_n155, Z => 
                           mult_28_C93_n151);
   mult_28_C93_U142 : OAI21D1 port map( A1 => mult_28_C93_n171, A2 => 
                           mult_28_C93_n150, B => mult_28_C93_n151, Z => 
                           mult_28_C93_n149);
   mult_28_C93_U132 : AOI21D1 port map( A1 => mult_28_C93_n155, A2 => 
                           mult_28_C93_n143, B => mult_28_C93_n144, Z => 
                           mult_28_C93_n142);
   mult_28_C93_U130 : OAI21D1 port map( A1 => mult_28_C93_n141, A2 => 
                           mult_28_C93_n166, B => mult_28_C93_n142, Z => 
                           mult_28_C93_n140);
   mult_28_C93_U128 : AOI21D1 port map( A1 => mult_28_C93_n173, A2 => 
                           mult_28_C93_n139, B => mult_28_C93_n140, Z => 
                           mult_28_C93_n138);
   mult_28_C93_U123 : EXOR2D1 port map( A1 => mult_28_C93_n147, A2 => 
                           mult_28_C93_n60, Z => m2_9);
   mult_28_C93_U121 : NOR2D2 port map( A1 => mult_28_C93_n332, A2 => 
                           mult_28_C93_n337, Z => mult_28_C93_n132);
   mult_28_C93_U116 : OAI21D1 port map( A1 => mult_28_C93_n52, A2 => 
                           mult_28_C93_n130, B => mult_28_C93_n133, Z => 
                           mult_28_C93_n129);
   mult_28_C93_U113 : EXOR2D1 port map( A1 => mult_28_C93_n134, A2 => 
                           mult_28_C93_n59, Z => m2_10);
   mult_28_C93_U108 : OAI21D1 port map( A1 => mult_28_C93_n133, A2 => 
                           mult_28_C93_n125, B => mult_28_C93_n126, Z => 
                           mult_28_C93_n124);
   mult_28_C93_U97 : EXOR2D1 port map( A1 => mult_28_C93_n127, A2 => 
                           mult_28_C93_n58, Z => m2_11);
   mult_28_C93_U88 : OAI21D1 port map( A1 => mult_28_C93_n52, A2 => 
                           mult_28_C93_n108, B => mult_28_C93_n109, Z => 
                           mult_28_C93_n107);
   mult_28_C93_U85 : EXOR2D1 port map( A1 => mult_28_C93_n114, A2 => 
                           mult_28_C93_n57, Z => m2_12);
   mult_28_C93_U80 : OAI21D1 port map( A1 => mult_28_C93_n113, A2 => 
                           mult_28_C93_n103, B => mult_28_C93_n104, Z => 
                           mult_28_C93_n102);
   mult_28_C93_U78 : AOI21D1 port map( A1 => mult_28_C93_n124, A2 => 
                           mult_28_C93_n101, B => mult_28_C93_n102, Z => 
                           mult_28_C93_n100);
   mult_28_C93_U74 : OAI21D1 port map( A1 => mult_28_C93_n52, A2 => 
                           mult_28_C93_n97, B => mult_28_C93_n100, Z => 
                           mult_28_C93_n96);
   mult_28_C93_U71 : EXOR2D1 port map( A1 => mult_28_C93_n105, A2 => 
                           mult_28_C93_n56, Z => m2_13);
   mult_28_C93_U62 : OAI21D1 port map( A1 => mult_28_C93_n52, A2 => 
                           mult_28_C93_n918, B => mult_28_C93_n917, Z => 
                           mult_28_C93_n87);
   mult_28_C93_U60 : AOI21D1 port map( A1 => mult_28_C93_n51, A2 => 
                           mult_28_C93_n86, B => mult_28_C93_n87, Z => 
                           mult_28_C93_n85);
   mult_28_C93_U59 : EXOR2D1 port map( A1 => mult_28_C93_n94, A2 => 
                           mult_28_C93_n55, Z => m2_14);
   mult_28_C93_U54 : EXOR2D1 port map( A1 => mult_28_C93_n85, A2 => 
                           mult_28_C93_n54, Z => m2_15);
   add_1_root_add_0_root_add_101_U241 : NOR2D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n59, A2 => 
                           add_1_root_add_0_root_add_101_n52, Z => 
                           add_1_root_add_0_root_add_101_n50);
   add_1_root_add_0_root_add_101_U240 : NAN2D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n122, A2 => 
                           add_1_root_add_0_root_add_101_n53, Z => 
                           add_1_root_add_0_root_add_101_n8);
   add_1_root_add_0_root_add_101_U239 : NAN2DL port map( A1 => z1_11_port, A2 
                           => m2_11, Z => add_1_root_add_0_root_add_101_n53);
   add_1_root_add_0_root_add_101_U238 : OR2D1 port map( A1 => z1_15_port, A2 =>
                           m2_15, Z => add_1_root_add_0_root_add_101_n193);
   add_1_root_add_0_root_add_101_U237 : NOR2D1 port map( A1 => z1_14_port, A2 
                           => m2_14, Z => add_1_root_add_0_root_add_101_n29);
   add_1_root_add_0_root_add_101_U236 : NAN2DL port map( A1 => z1_13_port, A2 
                           => m2_13, Z => add_1_root_add_0_root_add_101_n39);
   add_1_root_add_0_root_add_101_U235 : NAN2DL port map( A1 => z1_12_port, A2 
                           => m2_12, Z => add_1_root_add_0_root_add_101_n46);
   add_1_root_add_0_root_add_101_U234 : NOR2D1 port map( A1 => z1_13_port, A2 
                           => m2_13, Z => add_1_root_add_0_root_add_101_n38);
   add_1_root_add_0_root_add_101_U233 : NAN2D1 port map( A1 => z1_0_port, A2 =>
                           m2_0, Z => add_1_root_add_0_root_add_101_n117);
   add_1_root_add_0_root_add_101_U232 : NAN2D1 port map( A1 => z1_2_port, A2 =>
                           m2_2, Z => add_1_root_add_0_root_add_101_n111);
   add_1_root_add_0_root_add_101_U231 : NAN2DL port map( A1 => z1_1_port, A2 =>
                           m2_1, Z => add_1_root_add_0_root_add_101_n115);
   add_1_root_add_0_root_add_101_U230 : NOR2D1 port map( A1 => z1_11_port, A2 
                           => m2_11, Z => add_1_root_add_0_root_add_101_n52);
   add_1_root_add_0_root_add_101_U229 : NAN2DL port map( A1 => z1_15_port, A2 
                           => m2_15, Z => add_1_root_add_0_root_add_101_n21);
   add_1_root_add_0_root_add_101_U228 : NAN2D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n193, A2 => 
                           add_1_root_add_0_root_add_101_n21, Z => 
                           add_1_root_add_0_root_add_101_n4);
   add_1_root_add_0_root_add_101_U227 : NOR2D1 port map( A1 => z1_8_port, A2 =>
                           m2_8, Z => add_1_root_add_0_root_add_101_n73);
   add_1_root_add_0_root_add_101_U226 : NOR2D1 port map( A1 => z1_1_port, A2 =>
                           m2_1, Z => add_1_root_add_0_root_add_101_n114);
   add_1_root_add_0_root_add_101_U225 : INVDL port map( A => 
                           add_1_root_add_0_root_add_101_n102, Z => 
                           add_1_root_add_0_root_add_101_n100);
   add_1_root_add_0_root_add_101_U224 : INVDL port map( A => 
                           add_1_root_add_0_root_add_101_n101, Z => 
                           add_1_root_add_0_root_add_101_n99);
   add_1_root_add_0_root_add_101_U223 : INVDL port map( A => 
                           add_1_root_add_0_root_add_101_n107, Z => 
                           add_1_root_add_0_root_add_101_n130);
   add_1_root_add_0_root_add_101_U222 : INVDL port map( A => 
                           add_1_root_add_0_root_add_101_n74, Z => 
                           add_1_root_add_0_root_add_101_n72);
   add_1_root_add_0_root_add_101_U221 : INVDL port map( A => 
                           add_1_root_add_0_root_add_101_n45, Z => 
                           add_1_root_add_0_root_add_101_n44);
   add_1_root_add_0_root_add_101_U220 : INVD1 port map( A => 
                           add_1_root_add_0_root_add_101_n44, Z => 
                           add_1_root_add_0_root_add_101_n43);
   add_1_root_add_0_root_add_101_U219 : INVDL port map( A => 
                           add_1_root_add_0_root_add_101_n59, Z => 
                           add_1_root_add_0_root_add_101_n58);
   add_1_root_add_0_root_add_101_U218 : INVD1 port map( A => 
                           add_1_root_add_0_root_add_101_n58, Z => 
                           add_1_root_add_0_root_add_101_n57);
   add_1_root_add_0_root_add_101_U217 : INVDL port map( A => 
                           add_1_root_add_0_root_add_101_n96, Z => 
                           add_1_root_add_0_root_add_101_n128);
   add_1_root_add_0_root_add_101_U216 : INVDL port map( A => 
                           add_1_root_add_0_root_add_101_n87, Z => 
                           add_1_root_add_0_root_add_101_n86);
   add_1_root_add_0_root_add_101_U215 : INVDL port map( A => 
                           add_1_root_add_0_root_add_101_n80, Z => 
                           add_1_root_add_0_root_add_101_n126);
   add_1_root_add_0_root_add_101_U214 : NOR2D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n73, A2 => 
                           add_1_root_add_0_root_add_101_n68, Z => 
                           add_1_root_add_0_root_add_101_n66);
   add_1_root_add_0_root_add_101_U213 : INVDL port map( A => 
                           add_1_root_add_0_root_add_101_n68, Z => 
                           add_1_root_add_0_root_add_101_n124);
   add_1_root_add_0_root_add_101_U212 : NOR2D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n87, A2 => 
                           add_1_root_add_0_root_add_101_n80, Z => 
                           add_1_root_add_0_root_add_101_n78);
   add_1_root_add_0_root_add_101_U211 : INVD1 port map( A => 
                           add_1_root_add_0_root_add_101_n113, Z => 
                           add_1_root_add_0_root_add_101_n112);
   add_1_root_add_0_root_add_101_U210 : NAN2D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n36, A2 => 
                           add_1_root_add_0_root_add_101_n27, Z => 
                           add_1_root_add_0_root_add_101_n25);
   add_1_root_add_0_root_add_101_U209 : INVD1 port map( A => 
                           add_1_root_add_0_root_add_101_n36, Z => 
                           add_1_root_add_0_root_add_101_n34);
   add_1_root_add_0_root_add_101_U208 : INVD1 port map( A => 
                           add_1_root_add_0_root_add_101_n104, Z => 
                           add_1_root_add_0_root_add_101_n103);
   add_1_root_add_0_root_add_101_U207 : NOR2D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n92, A2 => 
                           add_1_root_add_0_root_add_101_n85, Z => 
                           add_1_root_add_0_root_add_101_n83);
   add_1_root_add_0_root_add_101_U206 : INVDL port map( A => 
                           add_1_root_add_0_root_add_101_n95, Z => 
                           add_1_root_add_0_root_add_101_n93);
   add_1_root_add_0_root_add_101_U205 : INVD1 port map( A => 
                           add_1_root_add_0_root_add_101_n66, Z => 
                           add_1_root_add_0_root_add_101_n64);
   add_1_root_add_0_root_add_101_U204 : INVDL port map( A => 
                           add_1_root_add_0_root_add_101_n67, Z => 
                           add_1_root_add_0_root_add_101_n65);
   add_1_root_add_0_root_add_101_U203 : NOR2D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n3, A2 => 
                           add_1_root_add_0_root_add_101_n43, Z => 
                           add_1_root_add_0_root_add_101_n41);
   add_1_root_add_0_root_add_101_U202 : NAN2D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n66, A2 => 
                           add_1_root_add_0_root_add_101_n50, Z => 
                           add_1_root_add_0_root_add_101_n3);
   add_1_root_add_0_root_add_101_U201 : NAN2D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n94, A2 => 
                           add_1_root_add_0_root_add_101_n78, Z => 
                           add_1_root_add_0_root_add_101_n76);
   add_1_root_add_0_root_add_101_U200 : BUFD4 port map( A => 
                           add_1_root_add_0_root_add_101_n75, Z => 
                           add_1_root_add_0_root_add_101_n1);
   add_1_root_add_0_root_add_101_U199 : INVD1 port map( A => 
                           add_1_root_add_0_root_add_101_n37, Z => 
                           add_1_root_add_0_root_add_101_n35);
   add_1_root_add_0_root_add_101_U198 : INVDL port map( A => 
                           add_1_root_add_0_root_add_101_n2, Z => 
                           add_1_root_add_0_root_add_101_n49);
   add_1_root_add_0_root_add_101_U197 : AND2DL port map( A1 => 
                           add_1_root_add_0_root_add_101_n189, A2 => 
                           add_1_root_add_0_root_add_101_n117, Z => z2_temp_0);
   add_1_root_add_0_root_add_101_U196 : NAN2DL port map( A1 => z1_14_port, A2 
                           => m2_14, Z => add_1_root_add_0_root_add_101_n30);
   add_1_root_add_0_root_add_101_U195 : NAN2D1 port map( A1 => z1_3_port, A2 =>
                           m2_3, Z => add_1_root_add_0_root_add_101_n108);
   add_1_root_add_0_root_add_101_U194 : NAN2D1 port map( A1 => z1_10_port, A2 
                           => m2_10, Z => add_1_root_add_0_root_add_101_n60);
   add_1_root_add_0_root_add_101_U193 : NAN2D1 port map( A1 => z1_9_port, A2 =>
                           m2_9, Z => add_1_root_add_0_root_add_101_n69);
   add_1_root_add_0_root_add_101_U192 : NAN2D1 port map( A1 => z1_5_port, A2 =>
                           m2_5, Z => add_1_root_add_0_root_add_101_n97);
   add_1_root_add_0_root_add_101_U191 : NAN2D1 port map( A1 => z1_7_port, A2 =>
                           m2_7, Z => add_1_root_add_0_root_add_101_n81);
   add_1_root_add_0_root_add_101_U190 : INVDL port map( A => 
                           add_1_root_add_0_root_add_101_n29, Z => 
                           add_1_root_add_0_root_add_101_n27);
   add_1_root_add_0_root_add_101_U189 : OAI21DL port map( A1 => 
                           add_1_root_add_0_root_add_101_n112, A2 => 
                           add_1_root_add_0_root_add_101_n110, B => 
                           add_1_root_add_0_root_add_101_n111, Z => 
                           add_1_root_add_0_root_add_101_n109);
   add_1_root_add_0_root_add_101_U188 : NOR2DL port map( A1 => 
                           add_1_root_add_0_root_add_101_n45, A2 => 
                           add_1_root_add_0_root_add_101_n38, Z => 
                           add_1_root_add_0_root_add_101_n36);
   add_1_root_add_0_root_add_101_U187 : NAN2M1DL port map( A1 => 
                           add_1_root_add_0_root_add_101_n114, A2 => 
                           add_1_root_add_0_root_add_101_n115, Z => 
                           add_1_root_add_0_root_add_101_n18);
   add_1_root_add_0_root_add_101_U186 : OA21M20DL port map( A1 => 
                           add_1_root_add_0_root_add_101_n37, A2 => 
                           add_1_root_add_0_root_add_101_n27, B => 
                           add_1_root_add_0_root_add_101_n30, Z => 
                           add_1_root_add_0_root_add_101_n26);
   add_1_root_add_0_root_add_101_U185 : NAN2M1DL port map( A1 => 
                           add_1_root_add_0_root_add_101_n110, A2 => 
                           add_1_root_add_0_root_add_101_n111, Z => 
                           add_1_root_add_0_root_add_101_n17);
   add_1_root_add_0_root_add_101_U184 : INVDL port map( A => 
                           add_1_root_add_0_root_add_101_n73, Z => 
                           add_1_root_add_0_root_add_101_n71);
   add_1_root_add_0_root_add_101_U183 : NAN2M1DL port map( A1 => 
                           add_1_root_add_0_root_add_101_n101, A2 => 
                           add_1_root_add_0_root_add_101_n102, Z => 
                           add_1_root_add_0_root_add_101_n15);
   add_1_root_add_0_root_add_101_U182 : INVD1 port map( A => 
                           add_1_root_add_0_root_add_101_n86, Z => 
                           add_1_root_add_0_root_add_101_n85);
   add_1_root_add_0_root_add_101_U181 : OAI21DL port map( A1 => 
                           add_1_root_add_0_root_add_101_n107, A2 => 
                           add_1_root_add_0_root_add_101_n111, B => 
                           add_1_root_add_0_root_add_101_n108, Z => 
                           add_1_root_add_0_root_add_101_n191);
   add_1_root_add_0_root_add_101_U180 : NOR2DL port map( A1 => 
                           add_1_root_add_0_root_add_101_n110, A2 => 
                           add_1_root_add_0_root_add_101_n107, Z => 
                           add_1_root_add_0_root_add_101_n190);
   add_1_root_add_0_root_add_101_U179 : AOI21D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n190, A2 => 
                           add_1_root_add_0_root_add_101_n113, B => 
                           add_1_root_add_0_root_add_101_n191, Z => 
                           add_1_root_add_0_root_add_101_n104);
   add_1_root_add_0_root_add_101_U178 : NAN2M1DL port map( A1 => 
                           add_1_root_add_0_root_add_101_n73, A2 => 
                           add_1_root_add_0_root_add_101_n74, Z => 
                           add_1_root_add_0_root_add_101_n11);
   add_1_root_add_0_root_add_101_U177 : NAN2M1DL port map( A1 => 
                           add_1_root_add_0_root_add_101_n45, A2 => 
                           add_1_root_add_0_root_add_101_n46, Z => 
                           add_1_root_add_0_root_add_101_n7);
   add_1_root_add_0_root_add_101_U176 : NAN2M1DL port map( A1 => 
                           add_1_root_add_0_root_add_101_n59, A2 => 
                           add_1_root_add_0_root_add_101_n60, Z => 
                           add_1_root_add_0_root_add_101_n9);
   add_1_root_add_0_root_add_101_U175 : INVDL port map( A => 
                           add_1_root_add_0_root_add_101_n52, Z => 
                           add_1_root_add_0_root_add_101_n122);
   add_1_root_add_0_root_add_101_U174 : NOR2DL port map( A1 => 
                           add_1_root_add_0_root_add_101_n64, A2 => 
                           add_1_root_add_0_root_add_101_n57, Z => 
                           add_1_root_add_0_root_add_101_n55);
   add_1_root_add_0_root_add_101_U173 : NOR2DL port map( A1 => 
                           add_1_root_add_0_root_add_101_n3, A2 => 
                           add_1_root_add_0_root_add_101_n25, Z => 
                           add_1_root_add_0_root_add_101_n23);
   add_1_root_add_0_root_add_101_U172 : NOR2DL port map( A1 => 
                           add_1_root_add_0_root_add_101_n3, A2 => 
                           add_1_root_add_0_root_add_101_n34, Z => 
                           add_1_root_add_0_root_add_101_n32);
   add_1_root_add_0_root_add_101_U171 : INVDL port map( A => 
                           add_1_root_add_0_root_add_101_n64, Z => 
                           add_1_root_add_0_root_add_101_n62);
   add_1_root_add_0_root_add_101_U170 : INVDL port map( A => 
                           add_1_root_add_0_root_add_101_n65, Z => 
                           add_1_root_add_0_root_add_101_n63);
   add_1_root_add_0_root_add_101_U169 : INVDL port map( A => 
                           add_1_root_add_0_root_add_101_n3, Z => 
                           add_1_root_add_0_root_add_101_n48);
   add_1_root_add_0_root_add_101_U168 : AOI21DL port map( A1 => 
                           add_1_root_add_0_root_add_101_n1, A2 => 
                           add_1_root_add_0_root_add_101_n32, B => 
                           add_1_root_add_0_root_add_101_n33, Z => 
                           add_1_root_add_0_root_add_101_n31);
   add_1_root_add_0_root_add_101_U167 : NAN2M1DL port map( A1 => 
                           add_1_root_add_0_root_add_101_n29, A2 => 
                           add_1_root_add_0_root_add_101_n30, Z => 
                           add_1_root_add_0_root_add_101_n5);
   add_1_root_add_0_root_add_101_U166 : AOI21DL port map( A1 => 
                           add_1_root_add_0_root_add_101_n1, A2 => 
                           add_1_root_add_0_root_add_101_n48, B => 
                           add_1_root_add_0_root_add_101_n49, Z => 
                           add_1_root_add_0_root_add_101_n47);
   add_1_root_add_0_root_add_101_U165 : NAN2M1DL port map( A1 => 
                           add_1_root_add_0_root_add_101_n38, A2 => 
                           add_1_root_add_0_root_add_101_n39, Z => 
                           add_1_root_add_0_root_add_101_n6);
   add_1_root_add_0_root_add_101_U164 : NOR2D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n101, A2 => 
                           add_1_root_add_0_root_add_101_n96, Z => 
                           add_1_root_add_0_root_add_101_n94);
   add_1_root_add_0_root_add_101_U163 : INVD1 port map( A => 
                           add_1_root_add_0_root_add_101_n94, Z => 
                           add_1_root_add_0_root_add_101_n92);
   add_1_root_add_0_root_add_101_U162 : NAN2DL port map( A1 => 
                           add_1_root_add_0_root_add_101_n128, A2 => 
                           add_1_root_add_0_root_add_101_n97, Z => 
                           add_1_root_add_0_root_add_101_n14);
   add_1_root_add_0_root_add_101_U161 : NAN2DL port map( A1 => 
                           add_1_root_add_0_root_add_101_n130, A2 => 
                           add_1_root_add_0_root_add_101_n108, Z => 
                           add_1_root_add_0_root_add_101_n16);
   add_1_root_add_0_root_add_101_U160 : NAN2DL port map( A1 => 
                           add_1_root_add_0_root_add_101_n126, A2 => 
                           add_1_root_add_0_root_add_101_n81, Z => 
                           add_1_root_add_0_root_add_101_n12);
   add_1_root_add_0_root_add_101_U159 : NAN2DL port map( A1 => 
                           add_1_root_add_0_root_add_101_n124, A2 => 
                           add_1_root_add_0_root_add_101_n69, Z => 
                           add_1_root_add_0_root_add_101_n10);
   add_1_root_add_0_root_add_101_U158 : NAN2DL port map( A1 => 
                           add_1_root_add_0_root_add_101_n86, A2 => 
                           add_1_root_add_0_root_add_101_n88, Z => 
                           add_1_root_add_0_root_add_101_n13);
   add_1_root_add_0_root_add_101_U157 : NAN2D1 port map( A1 => z1_4_port, A2 =>
                           m2_4, Z => add_1_root_add_0_root_add_101_n102);
   add_1_root_add_0_root_add_101_U156 : NOR2D1 port map( A1 => z1_2_port, A2 =>
                           m2_2, Z => add_1_root_add_0_root_add_101_n110);
   add_1_root_add_0_root_add_101_U155 : NAN2D1 port map( A1 => z1_8_port, A2 =>
                           m2_8, Z => add_1_root_add_0_root_add_101_n74);
   add_1_root_add_0_root_add_101_U154 : NAN2D1 port map( A1 => z1_6_port, A2 =>
                           m2_6, Z => add_1_root_add_0_root_add_101_n88);
   add_1_root_add_0_root_add_101_U153 : OR2DL port map( A1 => z1_0_port, A2 => 
                           m2_0, Z => add_1_root_add_0_root_add_101_n189);
   add_1_root_add_0_root_add_101_U140 : OAI21D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n114, A2 => 
                           add_1_root_add_0_root_add_101_n117, B => 
                           add_1_root_add_0_root_add_101_n115, Z => 
                           add_1_root_add_0_root_add_101_n113);
   add_1_root_add_0_root_add_101_U138 : EXOR2D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n18, A2 => 
                           add_1_root_add_0_root_add_101_n117, Z => z2_temp_1);
   add_1_root_add_0_root_add_101_U132 : EXOR2D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n112, A2 => 
                           add_1_root_add_0_root_add_101_n17, Z => z2_temp_2);
   add_1_root_add_0_root_add_101_U130 : NOR2D2 port map( A1 => z1_3_port, A2 =>
                           m2_3, Z => add_1_root_add_0_root_add_101_n107);
   add_1_root_add_0_root_add_101_U123 : EXNOR2D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n109, A2 => 
                           add_1_root_add_0_root_add_101_n16, Z => z2_temp_3);
   add_1_root_add_0_root_add_101_U121 : NOR2D2 port map( A1 => z1_4_port, A2 =>
                           m2_4, Z => add_1_root_add_0_root_add_101_n101);
   add_1_root_add_0_root_add_101_U116 : AOI21D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n103, A2 => 
                           add_1_root_add_0_root_add_101_n99, B => 
                           add_1_root_add_0_root_add_101_n100, Z => 
                           add_1_root_add_0_root_add_101_n98);
   add_1_root_add_0_root_add_101_U115 : EXNOR2D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n103, A2 => 
                           add_1_root_add_0_root_add_101_n15, Z => z2_temp_4);
   add_1_root_add_0_root_add_101_U113 : NOR2D2 port map( A1 => z1_5_port, A2 =>
                           m2_5, Z => add_1_root_add_0_root_add_101_n96);
   add_1_root_add_0_root_add_101_U110 : OAI21D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n96, A2 => 
                           add_1_root_add_0_root_add_101_n102, B => 
                           add_1_root_add_0_root_add_101_n97, Z => 
                           add_1_root_add_0_root_add_101_n95);
   add_1_root_add_0_root_add_101_U104 : AOI21D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n103, A2 => 
                           add_1_root_add_0_root_add_101_n94, B => 
                           add_1_root_add_0_root_add_101_n95, Z => 
                           add_1_root_add_0_root_add_101_n89);
   add_1_root_add_0_root_add_101_U103 : EXOR2D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n98, A2 => 
                           add_1_root_add_0_root_add_101_n14, Z => z2_temp_5);
   add_1_root_add_0_root_add_101_U101 : NOR2D2 port map( A1 => z1_6_port, A2 =>
                           m2_6, Z => add_1_root_add_0_root_add_101_n87);
   add_1_root_add_0_root_add_101_U96 : OAI21D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n93, A2 => 
                           add_1_root_add_0_root_add_101_n85, B => 
                           add_1_root_add_0_root_add_101_n88, Z => 
                           add_1_root_add_0_root_add_101_n84);
   add_1_root_add_0_root_add_101_U94 : AOI21D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n103, A2 => 
                           add_1_root_add_0_root_add_101_n83, B => 
                           add_1_root_add_0_root_add_101_n84, Z => 
                           add_1_root_add_0_root_add_101_n82);
   add_1_root_add_0_root_add_101_U93 : EXOR2D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n89, A2 => 
                           add_1_root_add_0_root_add_101_n13, Z => z2_temp_6);
   add_1_root_add_0_root_add_101_U91 : NOR2D2 port map( A1 => z1_7_port, A2 => 
                           m2_7, Z => add_1_root_add_0_root_add_101_n80);
   add_1_root_add_0_root_add_101_U88 : OAI21D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n80, A2 => 
                           add_1_root_add_0_root_add_101_n88, B => 
                           add_1_root_add_0_root_add_101_n81, Z => 
                           add_1_root_add_0_root_add_101_n79);
   add_1_root_add_0_root_add_101_U86 : AOI21D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n78, A2 => 
                           add_1_root_add_0_root_add_101_n95, B => 
                           add_1_root_add_0_root_add_101_n79, Z => 
                           add_1_root_add_0_root_add_101_n77);
   add_1_root_add_0_root_add_101_U84 : OAI21D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n104, A2 => 
                           add_1_root_add_0_root_add_101_n76, B => 
                           add_1_root_add_0_root_add_101_n77, Z => 
                           add_1_root_add_0_root_add_101_n75);
   add_1_root_add_0_root_add_101_U83 : EXOR2D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n82, A2 => 
                           add_1_root_add_0_root_add_101_n12, Z => z2_temp_7);
   add_1_root_add_0_root_add_101_U76 : AOI21D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n1, A2 => 
                           add_1_root_add_0_root_add_101_n71, B => 
                           add_1_root_add_0_root_add_101_n72, Z => 
                           add_1_root_add_0_root_add_101_n70);
   add_1_root_add_0_root_add_101_U75 : EXNOR2D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n1, A2 => 
                           add_1_root_add_0_root_add_101_n11, Z => z2_temp_8);
   add_1_root_add_0_root_add_101_U73 : NOR2D2 port map( A1 => z1_9_port, A2 => 
                           m2_9, Z => add_1_root_add_0_root_add_101_n68);
   add_1_root_add_0_root_add_101_U70 : OAI21D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n68, A2 => 
                           add_1_root_add_0_root_add_101_n74, B => 
                           add_1_root_add_0_root_add_101_n69, Z => 
                           add_1_root_add_0_root_add_101_n67);
   add_1_root_add_0_root_add_101_U64 : AOI21D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n1, A2 => 
                           add_1_root_add_0_root_add_101_n62, B => 
                           add_1_root_add_0_root_add_101_n63, Z => 
                           add_1_root_add_0_root_add_101_n61);
   add_1_root_add_0_root_add_101_U63 : EXOR2D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n70, A2 => 
                           add_1_root_add_0_root_add_101_n10, Z => z2_temp_9);
   add_1_root_add_0_root_add_101_U61 : NOR2D2 port map( A1 => z1_10_port, A2 =>
                           m2_10, Z => add_1_root_add_0_root_add_101_n59);
   add_1_root_add_0_root_add_101_U56 : OAI21D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n65, A2 => 
                           add_1_root_add_0_root_add_101_n57, B => 
                           add_1_root_add_0_root_add_101_n60, Z => 
                           add_1_root_add_0_root_add_101_n56);
   add_1_root_add_0_root_add_101_U54 : AOI21D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n1, A2 => 
                           add_1_root_add_0_root_add_101_n55, B => 
                           add_1_root_add_0_root_add_101_n56, Z => 
                           add_1_root_add_0_root_add_101_n54);
   add_1_root_add_0_root_add_101_U53 : EXOR2D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n61, A2 => 
                           add_1_root_add_0_root_add_101_n9, Z => z2_temp_10);
   add_1_root_add_0_root_add_101_U48 : OAI21D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n52, A2 => 
                           add_1_root_add_0_root_add_101_n60, B => 
                           add_1_root_add_0_root_add_101_n53, Z => 
                           add_1_root_add_0_root_add_101_n51);
   add_1_root_add_0_root_add_101_U46 : AOI21D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n50, A2 => 
                           add_1_root_add_0_root_add_101_n67, B => 
                           add_1_root_add_0_root_add_101_n51, Z => 
                           add_1_root_add_0_root_add_101_n2);
   add_1_root_add_0_root_add_101_U41 : EXOR2D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n54, A2 => 
                           add_1_root_add_0_root_add_101_n8, Z => z2_temp_11);
   add_1_root_add_0_root_add_101_U39 : NOR2D2 port map( A1 => z1_12_port, A2 =>
                           m2_12, Z => add_1_root_add_0_root_add_101_n45);
   add_1_root_add_0_root_add_101_U34 : OAI21D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n2, A2 => 
                           add_1_root_add_0_root_add_101_n43, B => 
                           add_1_root_add_0_root_add_101_n46, Z => 
                           add_1_root_add_0_root_add_101_n42);
   add_1_root_add_0_root_add_101_U32 : AOI21D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n1, A2 => 
                           add_1_root_add_0_root_add_101_n41, B => 
                           add_1_root_add_0_root_add_101_n42, Z => 
                           add_1_root_add_0_root_add_101_n40);
   add_1_root_add_0_root_add_101_U31 : EXOR2D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n47, A2 => 
                           add_1_root_add_0_root_add_101_n7, Z => z2_temp_12);
   add_1_root_add_0_root_add_101_U26 : OAI21D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n38, A2 => 
                           add_1_root_add_0_root_add_101_n46, B => 
                           add_1_root_add_0_root_add_101_n39, Z => 
                           add_1_root_add_0_root_add_101_n37);
   add_1_root_add_0_root_add_101_U22 : OAI21D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n2, A2 => 
                           add_1_root_add_0_root_add_101_n34, B => 
                           add_1_root_add_0_root_add_101_n35, Z => 
                           add_1_root_add_0_root_add_101_n33);
   add_1_root_add_0_root_add_101_U19 : EXOR2D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n40, A2 => 
                           add_1_root_add_0_root_add_101_n6, Z => z2_temp_13);
   add_1_root_add_0_root_add_101_U10 : OAI21D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n2, A2 => 
                           add_1_root_add_0_root_add_101_n25, B => 
                           add_1_root_add_0_root_add_101_n26, Z => 
                           add_1_root_add_0_root_add_101_n24);
   add_1_root_add_0_root_add_101_U8 : AOI21D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n1, A2 => 
                           add_1_root_add_0_root_add_101_n23, B => 
                           add_1_root_add_0_root_add_101_n24, Z => 
                           add_1_root_add_0_root_add_101_n22);
   add_1_root_add_0_root_add_101_U7 : EXOR2D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n31, A2 => 
                           add_1_root_add_0_root_add_101_n5, Z => z2_temp_14);
   add_1_root_add_0_root_add_101_U2 : EXOR2D1 port map( A1 => 
                           add_1_root_add_0_root_add_101_n22, A2 => 
                           add_1_root_add_0_root_add_101_n4, Z => z2_temp_15);
   mult_28_C92_U1384 : EXNOR2D4 port map( A1 => coeff_memory_75_port, A2 => 
                           coeff_memory_76_port, Z => mult_28_C92_n40);
   mult_28_C92_U1383 : EXNOR2D4 port map( A1 => coeff_memory_71_port, A2 => 
                           coeff_memory_72_port, Z => mult_28_C92_n28);
   mult_28_C92_U1382 : EXNOR2D4 port map( A1 => coeff_memory_65_port, A2 => 
                           coeff_memory_66_port, Z => mult_28_C92_n9);
   mult_28_C92_U1381 : AOI21DL port map( A1 => mult_28_C92_n128, A2 => 
                           mult_28_C92_net12273, B => mult_28_C92_n129, Z => 
                           mult_28_C92_n127);
   mult_28_C92_U1380 : AOI21DL port map( A1 => mult_28_C92_n135, A2 => 
                           mult_28_C92_net12273, B => mult_28_C92_n136, Z => 
                           mult_28_C92_n134);
   mult_28_C92_U1379 : AOI21DL port map( A1 => mult_28_C92_n106, A2 => 
                           mult_28_C92_net12273, B => mult_28_C92_n107, Z => 
                           mult_28_C92_n105);
   mult_28_C92_U1378 : AOI21DL port map( A1 => mult_28_C92_net12184, A2 => 
                           mult_28_C92_n86, B => mult_28_C92_n87, Z => 
                           mult_28_C92_n85);
   mult_28_C92_U1377 : OAI21DL port map( A1 => mult_28_C92_n1064, A2 => 
                           mult_28_C92_n108, B => mult_28_C92_n109, Z => 
                           mult_28_C92_n107);
   mult_28_C92_U1376 : OAI21DL port map( A1 => mult_28_C92_n1064, A2 => 
                           mult_28_C92_n97, B => mult_28_C92_n100, Z => 
                           mult_28_C92_n96);
   mult_28_C92_U1375 : OAI21DL port map( A1 => mult_28_C92_n1064, A2 => 
                           mult_28_C92_n1148, B => mult_28_C92_n1147, Z => 
                           mult_28_C92_n87);
   mult_28_C92_U1374 : AND2DL port map( A1 => mult_28_C92_n203, A2 => 
                           mult_28_C92_n298, Z => mult_28_C92_n1157);
   mult_28_C92_U1373 : EXNOR2D2 port map( A1 => mult_28_C92_n204, A2 => 
                           mult_28_C92_n1157, Z => m1_2);
   mult_28_C92_U1372 : EXNOR2D2 port map( A1 => mult_28_C92_n195, A2 => 
                           mult_28_C92_net9957, Z => m1_3);
   mult_28_C92_U1371 : EXOR2D1 port map( A1 => mult_28_C92_net12315, A2 => 
                           mult_28_C92_net9959, Z => m1_1);
   mult_28_C92_U1370 : NAN2DL port map( A1 => mult_28_C92_n412, A2 => 
                           mult_28_C92_n425, Z => mult_28_C92_n203);
   mult_28_C92_U1369 : EXNOR2DL port map( A1 => data_in(1), A2 => 
                           coeff_memory_69_port, Z => mult_28_C92_n758);
   mult_28_C92_U1368 : INVDL port map( A => mult_28_C92_n169, Z => 
                           mult_28_C92_n171);
   mult_28_C92_U1367 : INVDL port map( A => coeff_memory_65_port, Z => 
                           mult_28_C92_n842);
   mult_28_C92_U1366 : NAN2M1D2 port map( A1 => mult_28_C92_n1156, A2 => 
                           mult_28_C92_n834, Z => mult_28_C92_n6);
   mult_28_C92_U1365 : NAN2D2 port map( A1 => mult_28_C92_n811, A2 => 
                           mult_28_C92_n46, Z => mult_28_C92_n48);
   mult_28_C92_U1364 : EXNOR2D2 port map( A1 => coeff_memory_77_port, A2 => 
                           coeff_memory_78_port, Z => mult_28_C92_n46);
   mult_28_C92_U1363 : NAN2M1D2 port map( A1 => mult_28_C92_n1155, A2 => 
                           mult_28_C92_n9, Z => mult_28_C92_n12);
   mult_28_C92_U1362 : EXNOR2DL port map( A1 => coeff_memory_75_port, A2 => 
                           coeff_memory_74_port, Z => mult_28_C92_n1154);
   mult_28_C92_U1361 : NAN2M1D2 port map( A1 => mult_28_C92_n1154, A2 => 
                           mult_28_C92_n34, Z => mult_28_C92_n36);
   mult_28_C92_U1360 : NAN2D2 port map( A1 => mult_28_C92_n814, A2 => 
                           mult_28_C92_n28, Z => mult_28_C92_n30);
   mult_28_C92_U1359 : NAN2D2 port map( A1 => mult_28_C92_n812, A2 => 
                           mult_28_C92_n40, Z => mult_28_C92_n42);
   mult_28_C92_U1358 : INVDL port map( A => coeff_memory_79_port, Z => 
                           mult_28_C92_n835);
   mult_28_C92_U1357 : OR2D1 port map( A1 => mult_28_C92_n315, A2 => 
                           mult_28_C92_n942, Z => mult_28_C92_n1153);
   mult_28_C92_U1356 : AO21D1 port map( A1 => mult_28_C92_n42, A2 => 
                           mult_28_C92_n40, B => mult_28_C92_n676, Z => 
                           mult_28_C92_n547);
   mult_28_C92_U1355 : INVDL port map( A => mult_28_C92_n319, Z => 
                           mult_28_C92_n320);
   mult_28_C92_U1354 : AO21D1 port map( A1 => mult_28_C92_n36, A2 => 
                           mult_28_C92_n34, B => mult_28_C92_n693, Z => 
                           mult_28_C92_n563);
   mult_28_C92_U1353 : AO21D1 port map( A1 => mult_28_C92_n30, A2 => 
                           mult_28_C92_n28, B => mult_28_C92_n710, Z => 
                           mult_28_C92_n579);
   mult_28_C92_U1352 : INVD1 port map( A => mult_28_C92_n329, Z => 
                           mult_28_C92_n330);
   mult_28_C92_U1351 : AND2D1 port map( A1 => mult_28_C92_n658, A2 => 
                           mult_28_C92_n530, Z => mult_28_C92_n1152);
   mult_28_C92_U1350 : OR2D1 port map( A1 => mult_28_C92_n657, A2 => 
                           mult_28_C92_n642, Z => mult_28_C92_n1150);
   mult_28_C92_U1349 : NAN2D1 port map( A1 => mult_28_C92_n1153, A2 => 
                           mult_28_C92_n84, Z => mult_28_C92_n54);
   mult_28_C92_U1348 : NAN2DL port map( A1 => mult_28_C92_n522, A2 => 
                           mult_28_C92_n641, Z => mult_28_C92_n276);
   mult_28_C92_U1347 : INVDL port map( A => mult_28_C92_n361, Z => 
                           mult_28_C92_n362);
   mult_28_C92_U1346 : OR2D1 port map( A1 => mult_28_C92_n520, A2 => 
                           mult_28_C92_n521, Z => mult_28_C92_net10919);
   mult_28_C92_U1345 : AO21D1 port map( A1 => mult_28_C92_n24, A2 => 
                           mult_28_C92_n22, B => mult_28_C92_n727, Z => 
                           mult_28_C92_n595);
   mult_28_C92_U1344 : AO21D1 port map( A1 => mult_28_C92_n18, A2 => 
                           mult_28_C92_n16, B => mult_28_C92_n744, Z => 
                           mult_28_C92_n611);
   mult_28_C92_U1343 : OR2D1 port map( A1 => mult_28_C92_n512, A2 => 
                           mult_28_C92_n515, Z => mult_28_C92_net10923);
   mult_28_C92_U1342 : EXNOR2D1 port map( A1 => mult_28_C92_n600, A2 => 
                           mult_28_C92_n558, Z => mult_28_C92_n424);
   mult_28_C92_U1341 : AO21D1 port map( A1 => mult_28_C92_n12, A2 => 
                           mult_28_C92_n9, B => mult_28_C92_n761, Z => 
                           mult_28_C92_n627);
   mult_28_C92_U1340 : INVDL port map( A => mult_28_C92_n383, Z => 
                           mult_28_C92_n384);
   mult_28_C92_U1339 : NAN2DL port map( A1 => mult_28_C92_n317, A2 => 
                           mult_28_C92_n316, Z => mult_28_C92_n93);
   mult_28_C92_U1338 : NOR2D1 port map( A1 => mult_28_C92_n317, A2 => 
                           mult_28_C92_n316, Z => mult_28_C92_n92);
   mult_28_C92_U1337 : NAN2DL port map( A1 => mult_28_C92_n318, A2 => 
                           mult_28_C92_n321, Z => mult_28_C92_n104);
   mult_28_C92_U1336 : NOR2D1 port map( A1 => mult_28_C92_n318, A2 => 
                           mult_28_C92_n321, Z => mult_28_C92_n103);
   mult_28_C92_U1335 : NAN2D1 port map( A1 => mult_28_C92_n325, A2 => 
                           mult_28_C92_n322, Z => mult_28_C92_n113);
   mult_28_C92_U1334 : NOR2D1 port map( A1 => mult_28_C92_n325, A2 => 
                           mult_28_C92_n322, Z => mult_28_C92_n112);
   mult_28_C92_U1333 : INVD2 port map( A => mult_28_C92_n343, Z => 
                           mult_28_C92_n344);
   mult_28_C92_U1332 : OR2D1 port map( A1 => mult_28_C92_n506, A2 => 
                           mult_28_C92_n511, Z => mult_28_C92_n1149);
   mult_28_C92_U1331 : OR2D1 port map( A1 => mult_28_C92_n500, A2 => 
                           mult_28_C92_n505, Z => mult_28_C92_net11021);
   mult_28_C92_U1330 : INVDL port map( A => mult_28_C92_n409, Z => 
                           mult_28_C92_n410);
   mult_28_C92_U1329 : INVD1 port map( A => mult_28_C92_n112, Z => 
                           mult_28_C92_n288);
   mult_28_C92_U1328 : NAN2DL port map( A1 => mult_28_C92_n326, A2 => 
                           mult_28_C92_n331, Z => mult_28_C92_n126);
   mult_28_C92_U1327 : NAN2D1 port map( A1 => mult_28_C92_n332, A2 => 
                           mult_28_C92_n337, Z => mult_28_C92_n133);
   mult_28_C92_U1326 : OA21DL port map( A1 => mult_28_C92_n100, A2 => 
                           mult_28_C92_n92, B => mult_28_C92_n93, Z => 
                           mult_28_C92_n1147);
   mult_28_C92_U1325 : NAN2D1 port map( A1 => mult_28_C92_n338, A2 => 
                           mult_28_C92_n345, Z => mult_28_C92_n146);
   mult_28_C92_U1324 : OR2D1 port map( A1 => mult_28_C92_n338, A2 => 
                           mult_28_C92_n345, Z => mult_28_C92_n1146);
   mult_28_C92_U1323 : NAN2D1 port map( A1 => mult_28_C92_n354, A2 => 
                           mult_28_C92_n363, Z => mult_28_C92_n162);
   mult_28_C92_U1322 : OR2D1 port map( A1 => mult_28_C92_n346, A2 => 
                           mult_28_C92_n353, Z => mult_28_C92_n1145);
   mult_28_C92_U1321 : INVD1 port map( A => mult_28_C92_n103, Z => 
                           mult_28_C92_n287);
   mult_28_C92_U1320 : NOR2DL port map( A1 => mult_28_C92_n53, A2 => 
                           mult_28_C92_n117, Z => mult_28_C92_n115);
   mult_28_C92_U1319 : NAN2DL port map( A1 => mult_28_C92_n119, A2 => 
                           mult_28_C92_n101, Z => mult_28_C92_n97);
   mult_28_C92_U1318 : NOR2DL port map( A1 => mult_28_C92_n53, A2 => 
                           mult_28_C92_n1148, Z => mult_28_C92_n86);
   mult_28_C92_U1317 : NAN2D1 port map( A1 => mult_28_C92_n119, A2 => 
                           mult_28_C92_n288, Z => mult_28_C92_n108);
   mult_28_C92_U1316 : NOR2D1 port map( A1 => mult_28_C92_n130, A2 => 
                           mult_28_C92_n125, Z => mult_28_C92_n119);
   mult_28_C92_U1315 : INVDL port map( A => mult_28_C92_n161, Z => 
                           mult_28_C92_n293);
   mult_28_C92_U1314 : INVD1 port map( A => mult_28_C92_n157, Z => 
                           mult_28_C92_n155);
   mult_28_C92_U1313 : NAN2D1 port map( A1 => mult_28_C92_n1145, A2 => 
                           mult_28_C92_n1146, Z => mult_28_C92_n141);
   mult_28_C92_U1312 : NOR2D1 port map( A1 => mult_28_C92_n141, A2 => 
                           mult_28_C92_n161, Z => mult_28_C92_n139);
   mult_28_C92_U1311 : INVDL port map( A => mult_28_C92_n130, Z => 
                           mult_28_C92_n290);
   mult_28_C92_U1310 : NOR2D1 port map( A1 => mult_28_C92_n170, A2 => 
                           mult_28_C92_n150, Z => mult_28_C92_n148);
   mult_28_C92_U1309 : NOR2DL port map( A1 => mult_28_C92_n53, A2 => 
                           mult_28_C92_n97, Z => mult_28_C92_n95);
   mult_28_C92_U1308 : INVD1 port map( A => mult_28_C92_n168, Z => 
                           mult_28_C92_n170);
   mult_28_C92_U1307 : NOR2DL port map( A1 => mult_28_C92_n53, A2 => 
                           mult_28_C92_n108, Z => mult_28_C92_n106);
   mult_28_C92_U1306 : NAN2D1 port map( A1 => mult_28_C92_n168, A2 => 
                           mult_28_C92_n139, Z => mult_28_C92_n53);
   mult_28_C92_U1305 : INVDL port map( A => mult_28_C92_n1064, Z => 
                           mult_28_C92_n136);
   mult_28_C92_U1304 : INVDL port map( A => mult_28_C92_net12262, Z => 
                           mult_28_C92_n297);
   mult_28_C92_U1303 : EXNOR2DL port map( A1 => coeff_memory_65_port, A2 => 
                           coeff_memory_64_port, Z => mult_28_C92_n1156);
   mult_28_C92_U1302 : EXNOR2DL port map( A1 => coeff_memory_67_port, A2 => 
                           coeff_memory_66_port, Z => mult_28_C92_n1155);
   mult_28_C92_U1301 : EXNOR2DL port map( A1 => data_in(15), A2 => 
                           coeff_memory_79_port, Z => mult_28_C92_n659);
   mult_28_C92_U1300 : EXOR2DL port map( A1 => coeff_memory_69_port, A2 => 
                           coeff_memory_68_port, Z => mult_28_C92_n1143);
   mult_28_C92_U1299 : NAN2D2 port map( A1 => mult_28_C92_n1143, A2 => 
                           mult_28_C92_n16, Z => mult_28_C92_n18);
   mult_28_C92_U1298 : OAI22DL port map( A1 => mult_28_C92_n791, A2 => 
                           mult_28_C92_n6, B1 => mult_28_C92_n790, B2 => 
                           mult_28_C92_n834, Z => mult_28_C92_n656);
   mult_28_C92_U1297 : OAI22DL port map( A1 => mult_28_C92_n789, A2 => 
                           mult_28_C92_n6, B1 => mult_28_C92_n788, B2 => 
                           mult_28_C92_n834, Z => mult_28_C92_n654);
   mult_28_C92_U1296 : OAI22DL port map( A1 => mult_28_C92_n661, A2 => 
                           mult_28_C92_n48, B1 => mult_28_C92_n660, B2 => 
                           mult_28_C92_n46, Z => mult_28_C92_n532);
   mult_28_C92_U1295 : OAI22DL port map( A1 => mult_28_C92_n665, A2 => 
                           mult_28_C92_n48, B1 => mult_28_C92_n664, B2 => 
                           mult_28_C92_n46, Z => mult_28_C92_n536);
   mult_28_C92_U1294 : NAN2DL port map( A1 => mult_28_C92_n315, A2 => 
                           mult_28_C92_n942, Z => mult_28_C92_n84);
   mult_28_C92_U1293 : OAI22DL port map( A1 => mult_28_C92_n698, A2 => 
                           mult_28_C92_n36, B1 => mult_28_C92_n697, B2 => 
                           mult_28_C92_n34, Z => mult_28_C92_n567);
   mult_28_C92_U1292 : OAI22DL port map( A1 => mult_28_C92_n793, A2 => 
                           mult_28_C92_n6, B1 => mult_28_C92_n792, B2 => 
                           mult_28_C92_n834, Z => mult_28_C92_n658);
   mult_28_C92_U1291 : AND2DL port map( A1 => mult_28_C92_n657, A2 => 
                           mult_28_C92_n642, Z => mult_28_C92_n1151);
   mult_28_C92_U1290 : NOR2D1 port map( A1 => mult_28_C92_n522, A2 => 
                           mult_28_C92_n641, Z => mult_28_C92_n275);
   mult_28_C92_U1289 : NOR2D1 port map( A1 => mult_28_C92_n516, A2 => 
                           mult_28_C92_n519, Z => mult_28_C92_n267);
   mult_28_C92_U1288 : OR2DL port map( A1 => mult_28_C92_n97, A2 => 
                           mult_28_C92_n92, Z => mult_28_C92_n1148);
   mult_28_C92_U1287 : NAN2M1DL port map( A1 => mult_28_C92_n92, A2 => 
                           mult_28_C92_n93, Z => mult_28_C92_n55);
   mult_28_C92_U1286 : NAN2DL port map( A1 => mult_28_C92_n346, A2 => 
                           mult_28_C92_n353, Z => mult_28_C92_n157);
   mult_28_C92_U1285 : OA21M20DL port map( A1 => mult_28_C92_n120, A2 => 
                           mult_28_C92_n288, B => mult_28_C92_n113, Z => 
                           mult_28_C92_n109);
   mult_28_C92_U1284 : NAN2DL port map( A1 => mult_28_C92_n288, A2 => 
                           mult_28_C92_n113, Z => mult_28_C92_n57);
   mult_28_C92_U1283 : AND2DL port map( A1 => mult_28_C92_n287, A2 => 
                           mult_28_C92_n104, Z => mult_28_C92_n1142);
   mult_28_C92_U1282 : EXNOR2D2 port map( A1 => mult_28_C92_n105, A2 => 
                           mult_28_C92_n1142, Z => m1_13);
   mult_28_C92_U1281 : NOR2DL port map( A1 => mult_28_C92_n53, A2 => 
                           mult_28_C92_n130, Z => mult_28_C92_n128);
   mult_28_C92_U1280 : NAN2DL port map( A1 => mult_28_C92_n293, A2 => 
                           mult_28_C92_n1145, Z => mult_28_C92_n150);
   mult_28_C92_U1279 : OA21M20DL port map( A1 => mult_28_C92_n155, A2 => 
                           mult_28_C92_n1146, B => mult_28_C92_n146, Z => 
                           mult_28_C92_n142);
   mult_28_C92_U1278 : AOI21DL port map( A1 => mult_28_C92_n164, A2 => 
                           mult_28_C92_n1145, B => mult_28_C92_n155, Z => 
                           mult_28_C92_n151);
   mult_28_C92_U1277 : EXNOR2D2 port map( A1 => mult_28_C92_n127, A2 => 
                           mult_28_C92_n1144, Z => m1_11);
   mult_28_C92_U1276 : AND2DL port map( A1 => mult_28_C92_n289, A2 => 
                           mult_28_C92_n126, Z => mult_28_C92_n1144);
   mult_28_C92_U1275 : EXNOR2D2 port map( A1 => mult_28_C92_n134, A2 => 
                           mult_28_C92_n941, Z => m1_10);
   mult_28_C92_U1274 : NAN2DL port map( A1 => mult_28_C92_n1145, A2 => 
                           mult_28_C92_n157, Z => mult_28_C92_n61);
   mult_28_C92_U1273 : NAN2DL port map( A1 => mult_28_C92_n293, A2 => 
                           mult_28_C92_n162, Z => mult_28_C92_n62);
   mult_28_C92_U1272 : NAN2DL port map( A1 => mult_28_C92_n1146, A2 => 
                           mult_28_C92_n146, Z => mult_28_C92_n60);
   mult_28_C92_U1271 : INVDL port map( A => mult_28_C92_n119, Z => 
                           mult_28_C92_n117);
   mult_28_C92_U1270 : INVDL port map( A => mult_28_C92_n120, Z => 
                           mult_28_C92_n118);
   mult_28_C92_U1269 : EXNOR2D2 port map( A1 => mult_28_C92_n188, A2 => 
                           mult_28_C92_net11247, Z => m1_4);
   mult_28_C92_U1268 : INVDL port map( A => mult_28_C92_n53, Z => 
                           mult_28_C92_n135);
   mult_28_C92_U1267 : EXNOR2DL port map( A1 => mult_28_C92_n215, A2 => 
                           mult_28_C92_n69, Z => m1_0);
   mult_28_C92_U1266 : INVDL port map( A => mult_28_C92_n162, Z => 
                           mult_28_C92_n164);
   mult_28_C92_U1265 : EXNOR2D4 port map( A1 => coeff_memory_67_port, A2 => 
                           coeff_memory_68_port, Z => mult_28_C92_n16);
   mult_28_C92_U1264 : NAN2D2 port map( A1 => mult_28_C92_n1140, A2 => 
                           mult_28_C92_n1141, Z => mult_28_C92_n619);
   mult_28_C92_U1263 : NAN3D2 port map( A1 => mult_28_C92_n1137, A2 => 
                           mult_28_C92_n1139, A3 => mult_28_C92_n1138, Z => 
                           mult_28_C92_n479);
   mult_28_C92_U1262 : NAN2D1 port map( A1 => mult_28_C92_n577, A2 => 
                           mult_28_C92_n648, Z => mult_28_C92_n1139);
   mult_28_C92_U1261 : NAN2D1 port map( A1 => mult_28_C92_n619, A2 => 
                           mult_28_C92_n648, Z => mult_28_C92_n1138);
   mult_28_C92_U1260 : NAN2D1 port map( A1 => mult_28_C92_n619, A2 => 
                           mult_28_C92_n577, Z => mult_28_C92_n1137);
   mult_28_C92_U1259 : NOR2DL port map( A1 => mult_28_C92_n112, A2 => 
                           mult_28_C92_n103, Z => mult_28_C92_n101);
   mult_28_C92_U1258 : AOI21D1 port map( A1 => mult_28_C92_net12273, A2 => 
                           mult_28_C92_n168, B => mult_28_C92_n169, Z => 
                           mult_28_C92_n167);
   mult_28_C92_U1257 : EXOR2D2 port map( A1 => mult_28_C92_n167, A2 => 
                           mult_28_C92_n62, Z => m1_7);
   mult_28_C92_U1256 : EXOR2D4 port map( A1 => mult_28_C92_n943, A2 => 
                           mult_28_C92_n524, Z => mult_28_C92_n462);
   mult_28_C92_U1255 : NAN3D1 port map( A1 => mult_28_C92_n1134, A2 => 
                           mult_28_C92_n1135, A3 => mult_28_C92_n1136, Z => 
                           mult_28_C92_n439);
   mult_28_C92_U1254 : NAN2DL port map( A1 => mult_28_C92_n444, A2 => 
                           mult_28_C92_n442, Z => mult_28_C92_n1136);
   mult_28_C92_U1253 : NAN2DL port map( A1 => mult_28_C92_n453, A2 => 
                           mult_28_C92_n442, Z => mult_28_C92_n1135);
   mult_28_C92_U1252 : NAN2DL port map( A1 => mult_28_C92_n453, A2 => 
                           mult_28_C92_n444, Z => mult_28_C92_n1134);
   mult_28_C92_U1251 : NAN2DL port map( A1 => mult_28_C92_n446, A2 => 
                           mult_28_C92_n448, Z => mult_28_C92_n1133);
   mult_28_C92_U1250 : EXOR3D2 port map( A1 => mult_28_C92_n619, A2 => 
                           mult_28_C92_n648, A3 => mult_28_C92_n577, Z => 
                           mult_28_C92_n480);
   mult_28_C92_U1249 : INVDL port map( A => mult_28_C92_n1006, Z => 
                           mult_28_C92_n296);
   mult_28_C92_U1248 : NAN3D1 port map( A1 => mult_28_C92_n1130, A2 => 
                           mult_28_C92_n1132, A3 => mult_28_C92_n1131, Z => 
                           mult_28_C92_n391);
   mult_28_C92_U1247 : NAN2D1 port map( A1 => mult_28_C92_n407, A2 => 
                           mult_28_C92_n584, Z => mult_28_C92_n1130);
   mult_28_C92_U1246 : EXOR2D1 port map( A1 => mult_28_C92_n1129, A2 => 
                           mult_28_C92_n407, Z => mult_28_C92_n392);
   mult_28_C92_U1245 : EXNOR2DL port map( A1 => data_in(7), A2 => 
                           coeff_memory_65_port, Z => mult_28_C92_n786);
   mult_28_C92_U1244 : EXNOR2DL port map( A1 => data_in(7), A2 => 
                           coeff_memory_79_port, Z => mult_28_C92_n667);
   mult_28_C92_U1243 : EXNOR2DL port map( A1 => data_in(7), A2 => 
                           coeff_memory_67_port, Z => mult_28_C92_n769);
   mult_28_C92_U1242 : EXNOR2DL port map( A1 => data_in(7), A2 => 
                           coeff_memory_77_port, Z => mult_28_C92_n684);
   mult_28_C92_U1241 : NAN2DL port map( A1 => mult_28_C92_n416, A2 => 
                           mult_28_C92_n414, Z => mult_28_C92_n1125);
   mult_28_C92_U1240 : NAN2DL port map( A1 => mult_28_C92_n1103, A2 => 
                           mult_28_C92_n414, Z => mult_28_C92_n1124);
   mult_28_C92_U1239 : NAN2DL port map( A1 => mult_28_C92_n1103, A2 => 
                           mult_28_C92_n416, Z => mult_28_C92_n1123);
   mult_28_C92_U1238 : NAN3D2 port map( A1 => mult_28_C92_n1120, A2 => 
                           mult_28_C92_n1121, A3 => mult_28_C92_n1122, Z => 
                           mult_28_C92_n413);
   mult_28_C92_U1237 : NAN2D1 port map( A1 => mult_28_C92_n431, A2 => 
                           mult_28_C92_n418, Z => mult_28_C92_n1122);
   mult_28_C92_U1236 : NAN2D1 port map( A1 => mult_28_C92_n429, A2 => 
                           mult_28_C92_n418, Z => mult_28_C92_n1121);
   mult_28_C92_U1235 : NAN3D2 port map( A1 => mult_28_C92_n1117, A2 => 
                           mult_28_C92_n1119, A3 => mult_28_C92_n1118, Z => 
                           mult_28_C92_n429);
   mult_28_C92_U1234 : NAN2D1 port map( A1 => mult_28_C92_n445, A2 => 
                           mult_28_C92_n447, Z => mult_28_C92_n1119);
   mult_28_C92_U1233 : NAN2D1 port map( A1 => mult_28_C92_n434, A2 => 
                           mult_28_C92_n447, Z => mult_28_C92_n1118);
   mult_28_C92_U1232 : NAN2D1 port map( A1 => mult_28_C92_n434, A2 => 
                           mult_28_C92_n445, Z => mult_28_C92_n1117);
   mult_28_C92_U1231 : AOI21DL port map( A1 => mult_28_C92_n115, A2 => 
                           mult_28_C92_net12273, B => mult_28_C92_n116, Z => 
                           mult_28_C92_n114);
   mult_28_C92_U1230 : NAN3D1 port map( A1 => mult_28_C92_n1114, A2 => 
                           mult_28_C92_n1116, A3 => mult_28_C92_n1115, Z => 
                           mult_28_C92_n425);
   mult_28_C92_U1229 : NAN2DL port map( A1 => mult_28_C92_n430, A2 => 
                           mult_28_C92_n441, Z => mult_28_C92_n1116);
   mult_28_C92_U1228 : NAN2DL port map( A1 => mult_28_C92_n428, A2 => 
                           mult_28_C92_n430, Z => mult_28_C92_n1114);
   mult_28_C92_U1227 : NAN2D1 port map( A1 => data_in(7), A2 => 
                           coeff_memory_73_port, Z => mult_28_C92_n1127);
   mult_28_C92_U1226 : OAI22D1 port map( A1 => mult_28_C92_n671, A2 => 
                           mult_28_C92_n48, B1 => mult_28_C92_n670, B2 => 
                           mult_28_C92_n46, Z => mult_28_C92_n542);
   mult_28_C92_U1225 : EXNOR2DL port map( A1 => data_in(10), A2 => 
                           coeff_memory_65_port, Z => mult_28_C92_n1109);
   mult_28_C92_U1224 : NAN2D1 port map( A1 => data_in(3), A2 => 
                           coeff_memory_73_port, Z => mult_28_C92_n1111);
   mult_28_C92_U1223 : EXNOR2DL port map( A1 => data_in(7), A2 => 
                           coeff_memory_69_port, Z => mult_28_C92_n1108);
   mult_28_C92_U1222 : EXNOR2DL port map( A1 => data_in(11), A2 => 
                           coeff_memory_65_port, Z => mult_28_C92_n782);
   mult_28_C92_U1221 : EXNOR2DL port map( A1 => data_in(11), A2 => 
                           coeff_memory_65_port, Z => mult_28_C92_n1107);
   mult_28_C92_U1220 : EXNOR2DL port map( A1 => data_in(4), A2 => 
                           coeff_memory_73_port, Z => mult_28_C92_n1106);
   mult_28_C92_U1219 : EXNOR2DL port map( A1 => data_in(8), A2 => 
                           coeff_memory_69_port, Z => mult_28_C92_n1105);
   mult_28_C92_U1218 : OAI22DL port map( A1 => mult_28_C92_n785, A2 => 
                           mult_28_C92_n6, B1 => mult_28_C92_n784, B2 => 
                           mult_28_C92_n834, Z => mult_28_C92_n650);
   mult_28_C92_U1217 : OAI22D1 port map( A1 => mult_28_C92_n784, A2 => 
                           mult_28_C92_n6, B1 => mult_28_C92_n1109, B2 => 
                           mult_28_C92_n834, Z => mult_28_C92_n649);
   mult_28_C92_U1216 : EXOR2D1 port map( A1 => mult_28_C92_n147, A2 => 
                           mult_28_C92_n60, Z => m1_9);
   mult_28_C92_U1215 : EXNOR2DL port map( A1 => data_in(6), A2 => 
                           coeff_memory_69_port, Z => mult_28_C92_n1104);
   mult_28_C92_U1214 : INVDL port map( A => mult_28_C92_n1102, Z => 
                           mult_28_C92_n1103);
   mult_28_C92_U1213 : INVDL port map( A => mult_28_C92_n427, Z => 
                           mult_28_C92_n1102);
   mult_28_C92_U1212 : OAI22D2 port map( A1 => mult_28_C92_n764, A2 => 
                           mult_28_C92_n12, B1 => mult_28_C92_n1091, B2 => 
                           mult_28_C92_n9, Z => mult_28_C92_n629);
   mult_28_C92_U1211 : NAN3D1 port map( A1 => mult_28_C92_n1099, A2 => 
                           mult_28_C92_n1101, A3 => mult_28_C92_n1100, Z => 
                           mult_28_C92_n459);
   mult_28_C92_U1210 : NAN2DL port map( A1 => mult_28_C92_n646, A2 => 
                           mult_28_C92_n1083, Z => mult_28_C92_n1101);
   mult_28_C92_U1209 : NAN2DL port map( A1 => mult_28_C92_n1065, A2 => 
                           mult_28_C92_n1083, Z => mult_28_C92_n1100);
   mult_28_C92_U1208 : NAN2DL port map( A1 => mult_28_C92_n1065, A2 => 
                           mult_28_C92_n646, Z => mult_28_C92_n1099);
   mult_28_C92_U1207 : EXOR3D2 port map( A1 => mult_28_C92_n603, A2 => 
                           mult_28_C92_n631, A3 => mult_28_C92_n646, Z => 
                           mult_28_C92_n460);
   mult_28_C92_U1206 : NAN2D2 port map( A1 => mult_28_C92_n1127, A2 => 
                           mult_28_C92_n1128, Z => mult_28_C92_n718);
   mult_28_C92_U1205 : NAN2DL port map( A1 => mult_28_C92_n407, A2 => 
                           mult_28_C92_n570, Z => mult_28_C92_n1131);
   mult_28_C92_U1204 : NAN2DL port map( A1 => mult_28_C92_n584, A2 => 
                           mult_28_C92_n570, Z => mult_28_C92_n1132);
   mult_28_C92_U1203 : EXOR2DL port map( A1 => mult_28_C92_n570, A2 => 
                           mult_28_C92_n584, Z => mult_28_C92_n1129);
   mult_28_C92_U1202 : OAI22DL port map( A1 => mult_28_C92_n687, A2 => 
                           mult_28_C92_n42, B1 => mult_28_C92_n686, B2 => 
                           mult_28_C92_n40, Z => mult_28_C92_n557);
   mult_28_C92_U1201 : NAN2DL port map( A1 => mult_28_C92_n557, A2 => 
                           mult_28_C92_n585, Z => mult_28_C92_n1098);
   mult_28_C92_U1200 : NAN2DL port map( A1 => mult_28_C92_n599, A2 => 
                           mult_28_C92_n585, Z => mult_28_C92_n1097);
   mult_28_C92_U1199 : NAN2DL port map( A1 => mult_28_C92_n599, A2 => 
                           mult_28_C92_n557, Z => mult_28_C92_n1096);
   mult_28_C92_U1198 : NAN3D1 port map( A1 => mult_28_C92_n1094, A2 => 
                           mult_28_C92_n1095, A3 => mult_28_C92_n1093, Z => 
                           mult_28_C92_n401);
   mult_28_C92_U1197 : NAN2DL port map( A1 => mult_28_C92_n406, A2 => 
                           mult_28_C92_n419, Z => mult_28_C92_n1094);
   mult_28_C92_U1196 : NAN2DL port map( A1 => mult_28_C92_n406, A2 => 
                           mult_28_C92_n408, Z => mult_28_C92_n1093);
   mult_28_C92_U1195 : EXNOR2DL port map( A1 => data_in(13), A2 => 
                           coeff_memory_67_port, Z => mult_28_C92_n1091);
   mult_28_C92_U1194 : INVD16 port map( A => data_in(7), Z => mult_28_C92_n1126
                           );
   mult_28_C92_U1193 : NAN2D2 port map( A1 => mult_28_C92_n1126, A2 => 
                           mult_28_C92_n1056, Z => mult_28_C92_n1128);
   mult_28_C92_U1192 : EXNOR2DL port map( A1 => data_in(5), A2 => 
                           coeff_memory_73_port, Z => mult_28_C92_n720);
   mult_28_C92_U1191 : EXNOR2DL port map( A1 => data_in(5), A2 => 
                           coeff_memory_69_port, Z => mult_28_C92_n754);
   mult_28_C92_U1190 : EXNOR2DL port map( A1 => data_in(5), A2 => 
                           coeff_memory_79_port, Z => mult_28_C92_n669);
   mult_28_C92_U1189 : NAN2DL port map( A1 => mult_28_C92_n408, A2 => 
                           mult_28_C92_n419, Z => mult_28_C92_n1095);
   mult_28_C92_U1188 : EXOR3D1 port map( A1 => mult_28_C92_n419, A2 => 
                           mult_28_C92_n1052, A3 => mult_28_C92_n408, Z => 
                           mult_28_C92_n402);
   mult_28_C92_U1187 : EXNOR2DL port map( A1 => data_in(11), A2 => 
                           coeff_memory_69_port, Z => mult_28_C92_n1090);
   mult_28_C92_U1186 : EXOR3D2 port map( A1 => mult_28_C92_n434, A2 => 
                           mult_28_C92_n447, A3 => mult_28_C92_n445, Z => 
                           mult_28_C92_n430);
   mult_28_C92_U1185 : OAI22DL port map( A1 => mult_28_C92_n720, A2 => 
                           mult_28_C92_n30, B1 => mult_28_C92_n719, B2 => 
                           mult_28_C92_n28, Z => mult_28_C92_n588);
   mult_28_C92_U1184 : EXOR2D1 port map( A1 => data_in(1), A2 => 
                           mult_28_C92_n835, Z => mult_28_C92_n1089);
   mult_28_C92_U1183 : NAN2D2 port map( A1 => mult_28_C92_n1126, A2 => 
                           mult_28_C92_net12088, Z => mult_28_C92_n1088);
   mult_28_C92_U1182 : NAN2D1 port map( A1 => data_in(7), A2 => 
                           coeff_memory_69_port, Z => mult_28_C92_n1087);
   mult_28_C92_U1181 : EXNOR2D1 port map( A1 => data_in(6), A2 => 
                           coeff_memory_71_port, Z => mult_28_C92_n736);
   mult_28_C92_U1180 : EXOR2D1 port map( A1 => data_in(2), A2 => 
                           mult_28_C92_net11946, Z => mult_28_C92_n706);
   mult_28_C92_U1179 : NAN2D1 port map( A1 => mult_28_C92_n1085, A2 => 
                           mult_28_C92_n1086, Z => mult_28_C92_n705);
   mult_28_C92_U1178 : NAN3D2 port map( A1 => mult_28_C92_net11942, A2 => 
                           mult_28_C92_net11943, A3 => mult_28_C92_net11944, Z 
                           => mult_28_C92_n467);
   mult_28_C92_U1177 : OAI22D2 port map( A1 => mult_28_C92_n690, A2 => 
                           mult_28_C92_n42, B1 => mult_28_C92_n1045, B2 => 
                           mult_28_C92_n40, Z => mult_28_C92_n560);
   mult_28_C92_U1176 : OAI22D2 port map( A1 => mult_28_C92_n724, A2 => 
                           mult_28_C92_n30, B1 => mult_28_C92_n917, B2 => 
                           mult_28_C92_n28, Z => mult_28_C92_n592);
   mult_28_C92_U1175 : ADFULD2 port map( A => mult_28_C92_n592, B => 
                           mult_28_C92_n634, CI => mult_28_C92_n620, CO => 
                           mult_28_C92_n487, S => mult_28_C92_n488);
   mult_28_C92_U1174 : NAN2D2 port map( A1 => mult_28_C92_n1110, A2 => 
                           mult_28_C92_n1056, Z => mult_28_C92_n1112);
   mult_28_C92_U1173 : OAI22DL port map( A1 => mult_28_C92_n1066, A2 => 
                           mult_28_C92_n12, B1 => mult_28_C92_n765, B2 => 
                           mult_28_C92_n9, Z => mult_28_C92_n1083);
   mult_28_C92_U1172 : EXNOR2D1 port map( A1 => data_in(9), A2 => 
                           coeff_memory_69_port, Z => mult_28_C92_n750);
   mult_28_C92_U1171 : EXNOR2DL port map( A1 => data_in(14), A2 => 
                           coeff_memory_65_port, Z => mult_28_C92_n779);
   mult_28_C92_U1170 : EXNOR2DL port map( A1 => data_in(14), A2 => 
                           coeff_memory_65_port, Z => mult_28_C92_n1082);
   mult_28_C92_U1169 : NAN2D1 port map( A1 => data_in(3), A2 => 
                           coeff_memory_75_port, Z => mult_28_C92_n1085);
   mult_28_C92_U1168 : EXOR2D1 port map( A1 => data_in(1), A2 => 
                           mult_28_C92_n1056, Z => mult_28_C92_n724);
   mult_28_C92_U1167 : EXNOR2D1 port map( A1 => data_in(9), A2 => 
                           coeff_memory_65_port, Z => mult_28_C92_n784);
   mult_28_C92_U1166 : EXNOR2D2 port map( A1 => data_in(9), A2 => 
                           coeff_memory_71_port, Z => mult_28_C92_n733);
   mult_28_C92_U1165 : EXNOR2DL port map( A1 => data_in(9), A2 => 
                           coeff_memory_79_port, Z => mult_28_C92_n665);
   mult_28_C92_U1164 : ADFULDL port map( A => mult_28_C92_n383, B => 
                           mult_28_C92_n540, CI => mult_28_C92_n611, CO => 
                           mult_28_C92_n371, S => mult_28_C92_n372);
   mult_28_C92_U1163 : EXNOR2D1 port map( A1 => data_in(7), A2 => 
                           coeff_memory_71_port, Z => mult_28_C92_n735);
   mult_28_C92_U1162 : BUFDL port map( A => mult_28_C92_net12262, Z => 
                           mult_28_C92_net12005);
   mult_28_C92_U1161 : AOI21D1 port map( A1 => mult_28_C92_net11686, A2 => 
                           mult_28_C92_n189, B => mult_28_C92_n190, Z => 
                           mult_28_C92_n188);
   mult_28_C92_U1160 : NAN2D2 port map( A1 => mult_28_C92_n1084, A2 => 
                           mult_28_C92_net11946, Z => mult_28_C92_n1086);
   mult_28_C92_U1159 : NAN2D1 port map( A1 => mult_28_C92_n1085, A2 => 
                           mult_28_C92_n1086, Z => mult_28_C92_n1080);
   mult_28_C92_U1158 : INVDL port map( A => mult_28_C92_n441, Z => 
                           mult_28_C92_n1076);
   mult_28_C92_U1157 : NAN2D1 port map( A1 => mult_28_C92_n1076, A2 => 
                           mult_28_C92_n430, Z => mult_28_C92_n1079);
   mult_28_C92_U1156 : NAN2D1 port map( A1 => mult_28_C92_n1077, A2 => 
                           mult_28_C92_n441, Z => mult_28_C92_n1078);
   mult_28_C92_U1155 : INVD2 port map( A => data_in(8), Z => mult_28_C92_n1072)
                           ;
   mult_28_C92_U1154 : NAN2D1 port map( A1 => mult_28_C92_net11021, A2 => 
                           mult_28_C92_n1149, Z => mult_28_C92_net11339);
   mult_28_C92_U1153 : EXNOR2D1 port map( A1 => data_in(4), A2 => 
                           coeff_memory_73_port, Z => mult_28_C92_n721);
   mult_28_C92_U1152 : NAN3D2 port map( A1 => mult_28_C92_n1070, A2 => 
                           mult_28_C92_net12114, A3 => mult_28_C92_n1071, Z => 
                           mult_28_C92_n471);
   mult_28_C92_U1151 : NAN2DL port map( A1 => mult_28_C92_n590, A2 => 
                           mult_28_C92_n562, Z => mult_28_C92_n1071);
   mult_28_C92_U1150 : EXNOR2D1 port map( A1 => data_in(5), A2 => 
                           coeff_memory_77_port, Z => mult_28_C92_n686);
   mult_28_C92_U1149 : EXNOR2D1 port map( A1 => data_in(10), A2 => 
                           coeff_memory_67_port, Z => mult_28_C92_n766);
   mult_28_C92_U1148 : EXNOR2D2 port map( A1 => data_in(1), A2 => 
                           coeff_memory_75_port, Z => mult_28_C92_n707);
   mult_28_C92_U1147 : EXNOR2DL port map( A1 => data_in(3), A2 => 
                           coeff_memory_71_port, Z => mult_28_C92_n1069);
   mult_28_C92_U1146 : EXNOR2D2 port map( A1 => data_in(4), A2 => 
                           coeff_memory_69_port, Z => mult_28_C92_n755);
   mult_28_C92_U1145 : OAI22D1 port map( A1 => mult_28_C92_n781, A2 => 
                           mult_28_C92_n6, B1 => mult_28_C92_n780, B2 => 
                           mult_28_C92_n834, Z => mult_28_C92_n646);
   mult_28_C92_U1144 : OAI22DL port map( A1 => mult_28_C92_n758, A2 => 
                           mult_28_C92_n18, B1 => mult_28_C92_n757, B2 => 
                           mult_28_C92_n16, Z => mult_28_C92_n624);
   mult_28_C92_U1143 : INVD20 port map( A => data_in(3), Z => mult_28_C92_n1084
                           );
   mult_28_C92_U1142 : NAN2M1D1 port map( A1 => data_in(0), A2 => 
                           coeff_memory_77_port, Z => mult_28_C92_n692);
   mult_28_C92_U1141 : EXNOR2D1 port map( A1 => data_in(2), A2 => 
                           coeff_memory_69_port, Z => mult_28_C92_n757);
   mult_28_C92_U1140 : EXNOR2DL port map( A1 => data_in(10), A2 => 
                           coeff_memory_67_port, Z => mult_28_C92_n1066);
   mult_28_C92_U1139 : OAI22DL port map( A1 => mult_28_C92_n916, A2 => 
                           mult_28_C92_n24, B1 => mult_28_C92_n735, B2 => 
                           mult_28_C92_n22, Z => mult_28_C92_n1065);
   mult_28_C92_U1138 : OAI22D2 port map( A1 => mult_28_C92_n674, A2 => 
                           mult_28_C92_n48, B1 => mult_28_C92_n1089, B2 => 
                           mult_28_C92_n46, Z => mult_28_C92_n545);
   mult_28_C92_U1137 : BUFDL port map( A => mult_28_C92_net12273, Z => 
                           mult_28_C92_net12184);
   mult_28_C92_U1136 : OAI22D1 port map( A1 => mult_28_C92_n740, A2 => 
                           mult_28_C92_n24, B1 => mult_28_C92_n1069, B2 => 
                           mult_28_C92_n22, Z => mult_28_C92_n607);
   mult_28_C92_U1135 : ADFULD2 port map( A => mult_28_C92_n593, B => 
                           mult_28_C92_n621, CI => mult_28_C92_n635, CO => 
                           mult_28_C92_n495, S => mult_28_C92_n496);
   mult_28_C92_U1134 : NAN2D1 port map( A1 => mult_28_C92_n590, A2 => 
                           mult_28_C92_n647, Z => mult_28_C92_n1070);
   mult_28_C92_U1133 : AOI21DL port map( A1 => mult_28_C92_n169, A2 => 
                           mult_28_C92_n139, B => mult_28_C92_n140, Z => 
                           mult_28_C92_n52);
   mult_28_C92_U1132 : INVDL port map( A => coeff_memory_77_port, Z => 
                           mult_28_C92_n1061);
   mult_28_C92_U1131 : NAN2D1 port map( A1 => mult_28_C92_n1062, A2 => 
                           mult_28_C92_n1063, Z => mult_28_C92_n691);
   mult_28_C92_U1130 : NAN2D1 port map( A1 => mult_28_C92_net12321, A2 => 
                           mult_28_C92_n1061, Z => mult_28_C92_n1063);
   mult_28_C92_U1129 : NAN2DL port map( A1 => data_in(0), A2 => 
                           coeff_memory_77_port, Z => mult_28_C92_n1062);
   mult_28_C92_U1128 : INVD1 port map( A => mult_28_C92_n835, Z => 
                           mult_28_C92_n1058);
   mult_28_C92_U1127 : NAN2D1 port map( A1 => mult_28_C92_n1059, A2 => 
                           mult_28_C92_n1060, Z => mult_28_C92_n673);
   mult_28_C92_U1126 : NAN2D1 port map( A1 => mult_28_C92_n957, A2 => 
                           mult_28_C92_n835, Z => mult_28_C92_n1060);
   mult_28_C92_U1125 : NAN2D1 port map( A1 => data_in(1), A2 => 
                           mult_28_C92_n1058, Z => mult_28_C92_n1059);
   mult_28_C92_U1124 : EXOR2D1 port map( A1 => mult_28_C92_n158, A2 => 
                           mult_28_C92_n61, Z => m1_8);
   mult_28_C92_U1123 : NAN3D1 port map( A1 => mult_28_C92_n1133, A2 => 
                           mult_28_C92_net11523, A3 => mult_28_C92_net11524, Z 
                           => mult_28_C92_n441);
   mult_28_C92_U1122 : EXOR2D1 port map( A1 => data_in(8), A2 => 
                           mult_28_C92_n1056, Z => mult_28_C92_n717);
   mult_28_C92_U1121 : NOR2DL port map( A1 => mult_28_C92_n398, A2 => 
                           mult_28_C92_n411, Z => mult_28_C92_net12262);
   mult_28_C92_U1120 : INVD4 port map( A => data_in(14), Z => mult_28_C92_n1053
                           );
   mult_28_C92_U1119 : NAN2D2 port map( A1 => mult_28_C92_n1054, A2 => 
                           mult_28_C92_n1055, Z => mult_28_C92_n762);
   mult_28_C92_U1118 : NAN2D2 port map( A1 => mult_28_C92_n1053, A2 => 
                           mult_28_C92_net12160, Z => mult_28_C92_n1055);
   mult_28_C92_U1117 : NAN2D1 port map( A1 => data_in(14), A2 => 
                           coeff_memory_67_port, Z => mult_28_C92_n1054);
   mult_28_C92_U1116 : AOI21D1 port map( A1 => mult_28_C92_net12184, A2 => 
                           mult_28_C92_n95, B => mult_28_C92_n96, Z => 
                           mult_28_C92_n94);
   mult_28_C92_U1115 : EXNOR2DL port map( A1 => data_in(10), A2 => 
                           coeff_memory_75_port, Z => mult_28_C92_n698);
   mult_28_C92_U1114 : INVDL port map( A => mult_28_C92_n207, Z => 
                           mult_28_C92_n299);
   mult_28_C92_U1113 : INVD1 port map( A => mult_28_C92_n1051, Z => 
                           mult_28_C92_n1052);
   mult_28_C92_U1112 : INVDL port map( A => mult_28_C92_n406, Z => 
                           mult_28_C92_n1051);
   mult_28_C92_U1111 : NAN2D1 port map( A1 => mult_28_C92_n435, A2 => 
                           mult_28_C92_n437, Z => mult_28_C92_n1050);
   mult_28_C92_U1110 : NAN2DL port map( A1 => mult_28_C92_n424, A2 => 
                           mult_28_C92_n437, Z => mult_28_C92_n1049);
   mult_28_C92_U1109 : INVD16 port map( A => data_in(0), Z => 
                           mult_28_C92_net12321);
   mult_28_C92_U1108 : NAN2D1 port map( A1 => mult_28_C92_n1046, A2 => 
                           mult_28_C92_n1047, Z => mult_28_C92_n674);
   mult_28_C92_U1107 : NAN2D2 port map( A1 => mult_28_C92_net12321, A2 => 
                           mult_28_C92_n835, Z => mult_28_C92_n1047);
   mult_28_C92_U1106 : NAN2D1 port map( A1 => data_in(0), A2 => 
                           coeff_memory_79_port, Z => mult_28_C92_n1046);
   mult_28_C92_U1105 : EXNOR2D4 port map( A1 => coeff_memory_73_port, A2 => 
                           coeff_memory_74_port, Z => mult_28_C92_n34);
   mult_28_C92_U1104 : OAI22D1 port map( A1 => mult_28_C92_n34, A2 => 
                           mult_28_C92_n701, B1 => mult_28_C92_n702, B2 => 
                           mult_28_C92_n36, Z => mult_28_C92_n571);
   mult_28_C92_U1103 : EXNOR2DL port map( A1 => data_in(2), A2 => 
                           coeff_memory_77_port, Z => mult_28_C92_n1045);
   mult_28_C92_U1102 : EXNOR2D1 port map( A1 => mult_28_C92_net12273, A2 => 
                           mult_28_C92_n64, Z => m1_5);
   mult_28_C92_U1101 : NAN2D1 port map( A1 => data_in(8), A2 => 
                           coeff_memory_69_port, Z => mult_28_C92_n1073);
   mult_28_C92_U1100 : EXNOR2D4 port map( A1 => coeff_memory_69_port, A2 => 
                           coeff_memory_70_port, Z => mult_28_C92_n22);
   mult_28_C92_U1099 : EXOR2DL port map( A1 => coeff_memory_71_port, A2 => 
                           coeff_memory_70_port, Z => mult_28_C92_n1041);
   mult_28_C92_U1098 : NAN2D2 port map( A1 => mult_28_C92_n1041, A2 => 
                           mult_28_C92_n22, Z => mult_28_C92_n24);
   mult_28_C92_U1097 : NAN2D1 port map( A1 => data_in(5), A2 => 
                           coeff_memory_71_port, Z => mult_28_C92_n1043);
   mult_28_C92_U1096 : INVDL port map( A => coeff_memory_71_port, Z => 
                           mult_28_C92_net11920);
   mult_28_C92_U1095 : INVDL port map( A => mult_28_C92_n202, Z => 
                           mult_28_C92_n298);
   mult_28_C92_U1094 : INVDL port map( A => mult_28_C92_n954, Z => 
                           mult_28_C92_n206);
   mult_28_C92_U1093 : AND2D1 port map( A1 => mult_28_C92_n299, A2 => 
                           mult_28_C92_n954, Z => mult_28_C92_net9959);
   mult_28_C92_U1092 : NAN2DL port map( A1 => mult_28_C92_n386, A2 => 
                           mult_28_C92_n397, Z => mult_28_C92_n187);
   mult_28_C92_U1091 : INVDL port map( A => mult_28_C92_n400, Z => 
                           mult_28_C92_n1039);
   mult_28_C92_U1090 : INVD1 port map( A => mult_28_C92_n1039, Z => 
                           mult_28_C92_n1040);
   mult_28_C92_U1089 : EXOR3D1 port map( A1 => mult_28_C92_n413, A2 => 
                           mult_28_C92_n402, A3 => mult_28_C92_n1040, Z => 
                           mult_28_C92_n1038);
   mult_28_C92_U1088 : NAN2D1 port map( A1 => mult_28_C92_n300, A2 => 
                           mult_28_C92_n214, Z => mult_28_C92_n69);
   mult_28_C92_U1087 : INVDL port map( A => mult_28_C92_n213, Z => 
                           mult_28_C92_n300);
   mult_28_C92_U1086 : NOR2D1 port map( A1 => mult_28_C92_n213, A2 => 
                           mult_28_C92_n216, Z => mult_28_C92_n211);
   mult_28_C92_U1085 : INVDL port map( A => mult_28_C92_net11981, Z => 
                           mult_28_C92_net11982);
   mult_28_C92_U1084 : NAN3D1 port map( A1 => mult_28_C92_net9976, A2 => 
                           mult_28_C92_net9974, A3 => mult_28_C92_net9975, Z =>
                           mult_28_C92_n469);
   mult_28_C92_U1083 : NAN2DL port map( A1 => mult_28_C92_n446, A2 => 
                           mult_28_C92_n455, Z => mult_28_C92_net11523);
   mult_28_C92_U1082 : NAN2DL port map( A1 => mult_28_C92_n448, A2 => 
                           mult_28_C92_n455, Z => mult_28_C92_net11524);
   mult_28_C92_U1081 : EXOR3D1 port map( A1 => mult_28_C92_n446, A2 => 
                           mult_28_C92_n448, A3 => mult_28_C92_n455, Z => 
                           mult_28_C92_n442);
   mult_28_C92_U1080 : NAN3D2 port map( A1 => mult_28_C92_net9968, A2 => 
                           mult_28_C92_net9967, A3 => mult_28_C92_net9969, Z =>
                           mult_28_C92_n465);
   mult_28_C92_U1079 : NAN3M1D1 port map( A1 => mult_28_C92_net11961, A2 => 
                           mult_28_C92_net9971, A3 => mult_28_C92_net9972, Z =>
                           mult_28_C92_n463);
   mult_28_C92_U1078 : NAN2D1 port map( A1 => mult_28_C92_n440, A2 => 
                           mult_28_C92_n451, Z => mult_28_C92_n214);
   mult_28_C92_U1077 : ADFULDL port map( A => mult_28_C92_n465, B => 
                           mult_28_C92_n456, CI => mult_28_C92_n454, CO => 
                           mult_28_C92_n451, S => mult_28_C92_n452);
   mult_28_C92_U1076 : NAN3M1DL port map( A1 => mult_28_C92_net11961, A2 => 
                           mult_28_C92_net9971, A3 => mult_28_C92_net9972, Z =>
                           mult_28_C92_n1037);
   mult_28_C92_U1075 : NAN2D1 port map( A1 => mult_28_C92_n452, A2 => 
                           mult_28_C92_n1037, Z => mult_28_C92_n221);
   mult_28_C92_U1074 : AOI21DL port map( A1 => mult_28_C92_net12350, A2 => 
                           mult_28_C92_n218, B => mult_28_C92_n219, Z => 
                           mult_28_C92_net12187);
   mult_28_C92_U1073 : OAI21D1 port map( A1 => mult_28_C92_n217, A2 => 
                           mult_28_C92_n213, B => mult_28_C92_n214, Z => 
                           mult_28_C92_n212);
   mult_28_C92_U1072 : EXOR3D1 port map( A1 => mult_28_C92_n487, A2 => 
                           mult_28_C92_n489, A3 => mult_28_C92_n480, Z => 
                           mult_28_C92_n476);
   mult_28_C92_U1071 : NAN2D1 port map( A1 => mult_28_C92_n479, A2 => 
                           mult_28_C92_n618, Z => mult_28_C92_net11943);
   mult_28_C92_U1070 : NAN2D1 port map( A1 => mult_28_C92_n487, A2 => 
                           mult_28_C92_n489, Z => mult_28_C92_n1034);
   mult_28_C92_U1069 : NAN2D1 port map( A1 => mult_28_C92_n487, A2 => 
                           mult_28_C92_n480, Z => mult_28_C92_n1035);
   mult_28_C92_U1068 : NAN2D1 port map( A1 => mult_28_C92_n489, A2 => 
                           mult_28_C92_n480, Z => mult_28_C92_n1036);
   mult_28_C92_U1067 : NAN3D2 port map( A1 => mult_28_C92_n1034, A2 => 
                           mult_28_C92_n1035, A3 => mult_28_C92_n1036, Z => 
                           mult_28_C92_n475);
   mult_28_C92_U1066 : BUFDL port map( A => mult_28_C92_n479, Z => 
                           mult_28_C92_net12148);
   mult_28_C92_U1065 : EXOR2D1 port map( A1 => mult_28_C92_net11941, A2 => 
                           mult_28_C92_net12148, Z => mult_28_C92_n468);
   mult_28_C92_U1064 : NOR2M1DL port map( A1 => mult_28_C92_n955, A2 => 
                           mult_28_C92_net12005, Z => mult_28_C92_n189);
   mult_28_C92_U1063 : AND2DL port map( A1 => mult_28_C92_n296, A2 => 
                           mult_28_C92_n187, Z => mult_28_C92_net11247);
   mult_28_C92_U1062 : OAI21DL port map( A1 => mult_28_C92_n199, A2 => 
                           mult_28_C92_net12005, B => mult_28_C92_n1010, Z => 
                           mult_28_C92_n190);
   mult_28_C92_U1061 : NOR2D1 port map( A1 => mult_28_C92_n374, A2 => 
                           mult_28_C92_n385, Z => mult_28_C92_n179);
   mult_28_C92_U1060 : NOR2D1 port map( A1 => mult_28_C92_n191, A2 => 
                           mult_28_C92_n186, Z => mult_28_C92_n184);
   mult_28_C92_U1059 : AND2D1 port map( A1 => mult_28_C92_n184, A2 => 
                           mult_28_C92_n196, Z => mult_28_C92_net12274);
   mult_28_C92_U1058 : NOR2DL port map( A1 => mult_28_C92_n191, A2 => 
                           mult_28_C92_n186, Z => mult_28_C92_n1033);
   mult_28_C92_U1057 : OAI21DL port map( A1 => mult_28_C92_n194, A2 => 
                           mult_28_C92_n186, B => mult_28_C92_n187, Z => 
                           mult_28_C92_n185);
   mult_28_C92_U1056 : NOR2D1 port map( A1 => mult_28_C92_n179, A2 => 
                           mult_28_C92_n174, Z => mult_28_C92_n168);
   mult_28_C92_U1055 : NOR2D2 port map( A1 => mult_28_C92_n364, A2 => 
                           mult_28_C92_n373, Z => mult_28_C92_n174);
   mult_28_C92_U1054 : NAN2D1 port map( A1 => mult_28_C92_n364, A2 => 
                           mult_28_C92_n373, Z => mult_28_C92_n175);
   mult_28_C92_U1053 : NAN2DL port map( A1 => mult_28_C92_n295, A2 => 
                           mult_28_C92_n180, Z => mult_28_C92_n64);
   mult_28_C92_U1052 : INVDL port map( A => mult_28_C92_n179, Z => 
                           mult_28_C92_n295);
   mult_28_C92_U1051 : INVDL port map( A => mult_28_C92_n180, Z => 
                           mult_28_C92_n178);
   mult_28_C92_U1050 : AOI21D1 port map( A1 => mult_28_C92_net12273, A2 => 
                           mult_28_C92_n295, B => mult_28_C92_n178, Z => 
                           mult_28_C92_n176);
   mult_28_C92_U1049 : INVDL port map( A => mult_28_C92_n174, Z => 
                           mult_28_C92_n294);
   mult_28_C92_U1048 : EXOR2D2 port map( A1 => mult_28_C92_n176, A2 => 
                           mult_28_C92_n63, Z => m1_6);
   mult_28_C92_U1047 : NAN2DL port map( A1 => data_in(9), A2 => 
                           coeff_memory_67_port, Z => mult_28_C92_n1031);
   mult_28_C92_U1046 : NAN2D1 port map( A1 => mult_28_C92_net11996, A2 => 
                           mult_28_C92_net12160, Z => mult_28_C92_n1032);
   mult_28_C92_U1045 : NAN2D1 port map( A1 => mult_28_C92_n1031, A2 => 
                           mult_28_C92_n1032, Z => mult_28_C92_n767);
   mult_28_C92_U1044 : EXNOR2DL port map( A1 => coeff_memory_75_port, A2 => 
                           data_in(2), Z => mult_28_C92_n1029);
   mult_28_C92_U1043 : OAI22D1 port map( A1 => mult_28_C92_n707, A2 => 
                           mult_28_C92_n36, B1 => mult_28_C92_n1029, B2 => 
                           mult_28_C92_n34, Z => mult_28_C92_n576);
   mult_28_C92_U1042 : AND2D1 port map( A1 => mult_28_C92_n520, A2 => 
                           mult_28_C92_n521, Z => mult_28_C92_n1018);
   mult_28_C92_U1041 : NAN2DL port map( A1 => mult_28_C92_n516, A2 => 
                           mult_28_C92_n519, Z => mult_28_C92_n268);
   mult_28_C92_U1040 : AND2DL port map( A1 => mult_28_C92_n512, A2 => 
                           mult_28_C92_n515, Z => mult_28_C92_n1019);
   mult_28_C92_U1039 : AND2DL port map( A1 => mult_28_C92_n506, A2 => 
                           mult_28_C92_n511, Z => mult_28_C92_n1024);
   mult_28_C92_U1038 : AND2DL port map( A1 => mult_28_C92_n500, A2 => 
                           mult_28_C92_n505, Z => mult_28_C92_n1022);
   mult_28_C92_U1037 : OAI21D1 port map( A1 => mult_28_C92_net11339, A2 => 
                           mult_28_C92_n261, B => mult_28_C92_n250, Z => 
                           mult_28_C92_n248);
   mult_28_C92_U1036 : OR2D1 port map( A1 => mult_28_C92_n492, A2 => 
                           mult_28_C92_n499, Z => mult_28_C92_n1021);
   mult_28_C92_U1035 : AND2D1 port map( A1 => mult_28_C92_n492, A2 => 
                           mult_28_C92_n499, Z => mult_28_C92_n1020);
   mult_28_C92_U1034 : INVDL port map( A => mult_28_C92_n235, Z => 
                           mult_28_C92_n233);
   mult_28_C92_U1033 : EXOR3DL port map( A1 => mult_28_C92_n493, A2 => 
                           mult_28_C92_n488, A3 => mult_28_C92_n486, Z => 
                           mult_28_C92_n1026);
   mult_28_C92_U1032 : OR2D1 port map( A1 => mult_28_C92_n1026, A2 => 
                           mult_28_C92_n491, Z => mult_28_C92_n1023);
   mult_28_C92_U1031 : NAN2D1 port map( A1 => mult_28_C92_n233, A2 => 
                           mult_28_C92_n1023, Z => mult_28_C92_n231);
   mult_28_C92_U1030 : NAN2D1 port map( A1 => mult_28_C92_n484, A2 => 
                           mult_28_C92_n491, Z => mult_28_C92_n1025);
   mult_28_C92_U1029 : NAN2DL port map( A1 => mult_28_C92_n474, A2 => 
                           mult_28_C92_n483, Z => mult_28_C92_n1027);
   mult_28_C92_U1028 : AO21D1 port map( A1 => mult_28_C92_n230, A2 => 
                           mult_28_C92_n211, B => mult_28_C92_n212, Z => 
                           mult_28_C92_net12315);
   mult_28_C92_U1027 : OAI21D1 port map( A1 => mult_28_C92_n243, A2 => 
                           mult_28_C92_n231, B => mult_28_C92_n1028, Z => 
                           mult_28_C92_n230);
   mult_28_C92_U1026 : BUFDL port map( A => mult_28_C92_net12275, Z => 
                           mult_28_C92_net11686);
   mult_28_C92_U1025 : OAI21M20D2 port map( A1 => mult_28_C92_net12274, A2 => 
                           mult_28_C92_net12275, B => mult_28_C92_n183, Z => 
                           mult_28_C92_net12273);
   mult_28_C92_U1024 : AOI21DL port map( A1 => mult_28_C92_net12275, A2 => 
                           mult_28_C92_n956, B => mult_28_C92_n926, Z => 
                           mult_28_C92_n195);
   mult_28_C92_U1023 : NAN2D1 port map( A1 => mult_28_C92_n647, A2 => 
                           mult_28_C92_n562, Z => mult_28_C92_net12114);
   mult_28_C92_U1022 : NAN2DL port map( A1 => mult_28_C92_net11982, A2 => 
                           mult_28_C92_n632, Z => mult_28_C92_net9976);
   mult_28_C92_U1021 : NAN2DL port map( A1 => mult_28_C92_n576, A2 => 
                           mult_28_C92_n632, Z => mult_28_C92_net9974);
   mult_28_C92_U1020 : NAN2DL port map( A1 => mult_28_C92_net11982, A2 => 
                           mult_28_C92_n576, Z => mult_28_C92_net9975);
   mult_28_C92_U1019 : OAI22DL port map( A1 => mult_28_C92_n738, A2 => 
                           mult_28_C92_n24, B1 => mult_28_C92_n737, B2 => 
                           mult_28_C92_n22, Z => mult_28_C92_n605);
   mult_28_C92_U1018 : EXNOR2DL port map( A1 => data_in(9), A2 => 
                           coeff_memory_67_port, Z => mult_28_C92_n1017);
   mult_28_C92_U1017 : OAI22DL port map( A1 => mult_28_C92_n768, A2 => 
                           mult_28_C92_n12, B1 => mult_28_C92_n1017, B2 => 
                           mult_28_C92_n9, Z => mult_28_C92_n633);
   mult_28_C92_U1016 : OAI22D1 port map( A1 => mult_28_C92_n28, A2 => 
                           mult_28_C92_n722, B1 => mult_28_C92_n723, B2 => 
                           mult_28_C92_n30, Z => mult_28_C92_n591);
   mult_28_C92_U1015 : EXOR2DL port map( A1 => mult_28_C92_n618, A2 => 
                           mult_28_C92_n481, Z => mult_28_C92_net11941);
   mult_28_C92_U1014 : NAN2DL port map( A1 => mult_28_C92_n481, A2 => 
                           mult_28_C92_n618, Z => mult_28_C92_net11944);
   mult_28_C92_U1013 : NAN2D1 port map( A1 => mult_28_C92_n479, A2 => 
                           mult_28_C92_n481, Z => mult_28_C92_net11942);
   mult_28_C92_U1012 : EXOR3D1 port map( A1 => mult_28_C92_n562, A2 => 
                           mult_28_C92_n590, A3 => mult_28_C92_n647, Z => 
                           mult_28_C92_n472);
   mult_28_C92_U1011 : EXOR2D1 port map( A1 => mult_28_C92_n632, A2 => 
                           mult_28_C92_n604, Z => mult_28_C92_net11337);
   mult_28_C92_U1010 : NAN2DL port map( A1 => mult_28_C92_n477, A2 => 
                           mult_28_C92_n470, Z => mult_28_C92_net9968);
   mult_28_C92_U1009 : NAN2DL port map( A1 => mult_28_C92_n470, A2 => 
                           mult_28_C92_n472, Z => mult_28_C92_net9967);
   mult_28_C92_U1008 : EXOR2D2 port map( A1 => mult_28_C92_net11337, A2 => 
                           mult_28_C92_n576, Z => mult_28_C92_n470);
   mult_28_C92_U1007 : EXOR2D1 port map( A1 => mult_28_C92_net11797, A2 => 
                           mult_28_C92_n476, Z => mult_28_C92_n474);
   mult_28_C92_U1006 : AND2DL port map( A1 => mult_28_C92_n468, A2 => 
                           mult_28_C92_n475, Z => mult_28_C92_net11961);
   mult_28_C92_U1005 : NAN2DL port map( A1 => mult_28_C92_n475, A2 => 
                           mult_28_C92_n466, Z => mult_28_C92_net9972);
   mult_28_C92_U1004 : NAN2DL port map( A1 => mult_28_C92_n468, A2 => 
                           mult_28_C92_n466, Z => mult_28_C92_net9971);
   mult_28_C92_U1003 : NAN2DL port map( A1 => mult_28_C92_n476, A2 => 
                           mult_28_C92_n911, Z => mult_28_C92_n1015);
   mult_28_C92_U1002 : NAN2DL port map( A1 => mult_28_C92_n478, A2 => 
                           mult_28_C92_n476, Z => mult_28_C92_net11803);
   mult_28_C92_U1001 : EXNOR2D1 port map( A1 => mult_28_C92_n468, A2 => 
                           mult_28_C92_n475, Z => mult_28_C92_net11020);
   mult_28_C92_U1000 : EXOR3D1 port map( A1 => mult_28_C92_n470, A2 => 
                           mult_28_C92_n472, A3 => mult_28_C92_n477, Z => 
                           mult_28_C92_n466);
   mult_28_C92_U999 : INVDL port map( A => mult_28_C92_n466, Z => 
                           mult_28_C92_n1012);
   mult_28_C92_U998 : INVD1 port map( A => mult_28_C92_net11020, Z => 
                           mult_28_C92_n1011);
   mult_28_C92_U997 : NAN2D1 port map( A1 => mult_28_C92_n1013, A2 => 
                           mult_28_C92_n1014, Z => mult_28_C92_n464);
   mult_28_C92_U996 : NAN2D1 port map( A1 => mult_28_C92_n1011, A2 => 
                           mult_28_C92_n1012, Z => mult_28_C92_n1014);
   mult_28_C92_U995 : NAN2DL port map( A1 => mult_28_C92_net11020, A2 => 
                           mult_28_C92_n466, Z => mult_28_C92_n1013);
   mult_28_C92_U994 : NAN2D2 port map( A1 => mult_28_C92_n1042, A2 => 
                           mult_28_C92_net11920, Z => mult_28_C92_n1044);
   mult_28_C92_U993 : NAN2DL port map( A1 => mult_28_C92_n1038, A2 => 
                           mult_28_C92_n411, Z => mult_28_C92_n194);
   mult_28_C92_U992 : NAN2DL port map( A1 => mult_28_C92_n1038, A2 => 
                           mult_28_C92_n411, Z => mult_28_C92_n1010);
   mult_28_C92_U991 : INVD2 port map( A => mult_28_C92_n220, Z => 
                           mult_28_C92_n218);
   mult_28_C92_U990 : OR2D1 port map( A1 => mult_28_C92_n753, A2 => 
                           mult_28_C92_n18, Z => mult_28_C92_n1140);
   mult_28_C92_U989 : INVD2 port map( A => data_in(6), Z => mult_28_C92_n1007);
   mult_28_C92_U988 : NAN2D1 port map( A1 => mult_28_C92_n1008, A2 => 
                           mult_28_C92_n1009, Z => mult_28_C92_n753);
   mult_28_C92_U987 : NAN2D1 port map( A1 => mult_28_C92_n1007, A2 => 
                           mult_28_C92_net12088, Z => mult_28_C92_n1009);
   mult_28_C92_U986 : NAN2DL port map( A1 => data_in(6), A2 => 
                           coeff_memory_69_port, Z => mult_28_C92_n1008);
   mult_28_C92_U985 : OAI22D1 port map( A1 => mult_28_C92_n701, A2 => 
                           mult_28_C92_n36, B1 => mult_28_C92_n700, B2 => 
                           mult_28_C92_n34, Z => mult_28_C92_n570);
   mult_28_C92_U984 : NOR2DL port map( A1 => mult_28_C92_n397, A2 => 
                           mult_28_C92_n386, Z => mult_28_C92_n1006);
   mult_28_C92_U983 : INVD4 port map( A => data_in(7), Z => mult_28_C92_n1003);
   mult_28_C92_U982 : NAN2D2 port map( A1 => mult_28_C92_n1004, A2 => 
                           mult_28_C92_n1005, Z => mult_28_C92_n701);
   mult_28_C92_U981 : NAN2D2 port map( A1 => mult_28_C92_n1003, A2 => 
                           mult_28_C92_net11946, Z => mult_28_C92_n1005);
   mult_28_C92_U980 : NAN2D1 port map( A1 => data_in(7), A2 => 
                           coeff_memory_75_port, Z => mult_28_C92_n1004);
   mult_28_C92_U979 : EXNOR2D1 port map( A1 => data_in(2), A2 => 
                           coeff_memory_73_port, Z => mult_28_C92_n723);
   mult_28_C92_U978 : AO21M10DL port map( A2 => mult_28_C92_n230, A1 => 
                           mult_28_C92_n216, B => mult_28_C92_n1002, Z => 
                           mult_28_C92_n215);
   mult_28_C92_U977 : NAN3M1D1 port map( A1 => mult_28_C92_n940, A2 => 
                           mult_28_C92_n1015, A3 => mult_28_C92_net11803, Z => 
                           mult_28_C92_n473);
   mult_28_C92_U976 : INVDL port map( A => mult_28_C92_n527, Z => 
                           mult_28_C92_n1000);
   mult_28_C92_U975 : NAN2M1D1 port map( A1 => mult_28_C92_n1000, A2 => 
                           mult_28_C92_n623, Z => mult_28_C92_n1001);
   mult_28_C92_U974 : OAI21M10DL port map( A1 => mult_28_C92_n119, A2 => 
                           mult_28_C92_n52, B => mult_28_C92_n118, Z => 
                           mult_28_C92_n116);
   mult_28_C92_U973 : OAI21D1 port map( A1 => mult_28_C92_n235, A2 => 
                           mult_28_C92_n1025, B => mult_28_C92_n1027, Z => 
                           mult_28_C92_n999);
   mult_28_C92_U972 : OAI22D1 port map( A1 => mult_28_C92_n36, A2 => 
                           mult_28_C92_n705, B1 => mult_28_C92_n704, B2 => 
                           mult_28_C92_n34, Z => mult_28_C92_n574);
   mult_28_C92_U971 : INVDL port map( A => mult_28_C92_n473, Z => 
                           mult_28_C92_n998);
   mult_28_C92_U970 : INVDL port map( A => mult_28_C92_n464, Z => 
                           mult_28_C92_n997);
   mult_28_C92_U969 : OAI21M20D1 port map( A1 => mult_28_C92_n997, A2 => 
                           mult_28_C92_n998, B => mult_28_C92_n218, Z => 
                           mult_28_C92_n216);
   mult_28_C92_U968 : EXOR3D1 port map( A1 => mult_28_C92_n599, A2 => 
                           mult_28_C92_n585, A3 => mult_28_C92_n557, Z => 
                           mult_28_C92_n406);
   mult_28_C92_U967 : INVD1 port map( A => mult_28_C92_n212, Z => 
                           mult_28_C92_n996);
   mult_28_C92_U966 : OAI21M20D2 port map( A1 => mult_28_C92_n230, A2 => 
                           mult_28_C92_n211, B => mult_28_C92_n996, Z => 
                           mult_28_C92_net12275);
   mult_28_C92_U965 : OAI22D1 port map( A1 => mult_28_C92_n716, A2 => 
                           mult_28_C92_n28, B1 => mult_28_C92_n30, B2 => 
                           mult_28_C92_n1092, Z => mult_28_C92_n585);
   mult_28_C92_U964 : INVD20 port map( A => data_in(13), Z => mult_28_C92_n1067
                           );
   mult_28_C92_U963 : OAI21D1 port map( A1 => mult_28_C92_n1067, A2 => 
                           mult_28_C92_net12160, B => mult_28_C92_n1068, Z => 
                           mult_28_C92_n763);
   mult_28_C92_U962 : EXOR3D2 port map( A1 => mult_28_C92_n429, A2 => 
                           mult_28_C92_n431, A3 => mult_28_C92_n418, Z => 
                           mult_28_C92_n414);
   mult_28_C92_U961 : OAI22DL port map( A1 => mult_28_C92_n42, A2 => 
                           mult_28_C92_n1061, B1 => mult_28_C92_n692, B2 => 
                           mult_28_C92_n40, Z => mult_28_C92_n524);
   mult_28_C92_U960 : NAN3D2 port map( A1 => mult_28_C92_n1123, A2 => 
                           mult_28_C92_n1124, A3 => mult_28_C92_n1125, Z => 
                           mult_28_C92_n411);
   mult_28_C92_U959 : NAN2DL port map( A1 => mult_28_C92_n428, A2 => 
                           mult_28_C92_n441, Z => mult_28_C92_n1115);
   mult_28_C92_U958 : EXNOR2D1 port map( A1 => data_in(2), A2 => 
                           coeff_memory_79_port, Z => mult_28_C92_n1057);
   mult_28_C92_U957 : OAI22DL port map( A1 => mult_28_C92_n979, A2 => 
                           mult_28_C92_n18, B1 => mult_28_C92_n749, B2 => 
                           mult_28_C92_n16, Z => mult_28_C92_n616);
   mult_28_C92_U956 : NAN3D1 port map( A1 => mult_28_C92_n992, A2 => 
                           mult_28_C92_n990, A3 => mult_28_C92_n991, Z => 
                           mult_28_C92_n421);
   mult_28_C92_U955 : NAN2DL port map( A1 => mult_28_C92_n586, A2 => 
                           mult_28_C92_n643, Z => mult_28_C92_n992);
   mult_28_C92_U954 : NAN2DL port map( A1 => mult_28_C92_n544, A2 => 
                           mult_28_C92_n643, Z => mult_28_C92_n991);
   mult_28_C92_U953 : NAN2DL port map( A1 => mult_28_C92_n544, A2 => 
                           mult_28_C92_n586, Z => mult_28_C92_n990);
   mult_28_C92_U952 : EXOR2D1 port map( A1 => mult_28_C92_n485, A2 => 
                           mult_28_C92_n478, Z => mult_28_C92_net11797);
   mult_28_C92_U951 : OAI21DL port map( A1 => mult_28_C92_n52, A2 => 
                           mult_28_C92_n130, B => mult_28_C92_n133, Z => 
                           mult_28_C92_n129);
   mult_28_C92_U950 : EXNOR2D2 port map( A1 => data_in(6), A2 => 
                           coeff_memory_73_port, Z => mult_28_C92_n719);
   mult_28_C92_U949 : EXNOR2D1 port map( A1 => mult_28_C92_n453, A2 => 
                           mult_28_C92_n444, Z => mult_28_C92_n989);
   mult_28_C92_U948 : EXNOR2D2 port map( A1 => mult_28_C92_n989, A2 => 
                           mult_28_C92_n442, Z => mult_28_C92_n440);
   mult_28_C92_U947 : NAN2D2 port map( A1 => mult_28_C92_n987, A2 => 
                           mult_28_C92_n988, Z => mult_28_C92_n732);
   mult_28_C92_U946 : NAN2D2 port map( A1 => mult_28_C92_n986, A2 => 
                           mult_28_C92_net11920, Z => mult_28_C92_n988);
   mult_28_C92_U945 : NAN2D1 port map( A1 => data_in(10), A2 => 
                           coeff_memory_71_port, Z => mult_28_C92_n987);
   mult_28_C92_U944 : OAI22D1 port map( A1 => mult_28_C92_n28, A2 => 
                           mult_28_C92_n718, B1 => mult_28_C92_n719, B2 => 
                           mult_28_C92_n30, Z => mult_28_C92_n587);
   mult_28_C92_U943 : NAN3D1 port map( A1 => mult_28_C92_n983, A2 => 
                           mult_28_C92_n985, A3 => mult_28_C92_n984, Z => 
                           mult_28_C92_n445);
   mult_28_C92_U942 : NAN2D1 port map( A1 => mult_28_C92_n939, A2 => 
                           mult_28_C92_n602, Z => mult_28_C92_n985);
   mult_28_C92_U941 : NAN2DL port map( A1 => mult_28_C92_n616, A2 => 
                           mult_28_C92_n602, Z => mult_28_C92_n984);
   mult_28_C92_U940 : NAN2DL port map( A1 => mult_28_C92_n616, A2 => 
                           mult_28_C92_n939, Z => mult_28_C92_n983);
   mult_28_C92_U939 : EXOR3D1 port map( A1 => mult_28_C92_n602, A2 => 
                           mult_28_C92_n616, A3 => mult_28_C92_n939, Z => 
                           mult_28_C92_n446);
   mult_28_C92_U938 : INVD2 port map( A => data_in(12), Z => mult_28_C92_n980);
   mult_28_C92_U937 : NAN2D2 port map( A1 => mult_28_C92_n981, A2 => 
                           mult_28_C92_n982, Z => mult_28_C92_n747);
   mult_28_C92_U936 : NAN2D2 port map( A1 => mult_28_C92_n980, A2 => 
                           mult_28_C92_net12088, Z => mult_28_C92_n982);
   mult_28_C92_U935 : NAN2D1 port map( A1 => data_in(12), A2 => 
                           coeff_memory_69_port, Z => mult_28_C92_n981);
   mult_28_C92_U934 : AND2D1 port map( A1 => mult_28_C92_n297, A2 => 
                           mult_28_C92_n1010, Z => mult_28_C92_net9957);
   mult_28_C92_U933 : NAN2D1 port map( A1 => mult_28_C92_n994, A2 => 
                           mult_28_C92_n995, Z => mult_28_C92_n748);
   mult_28_C92_U932 : EXNOR2DL port map( A1 => data_in(9), A2 => 
                           coeff_memory_69_port, Z => mult_28_C92_n979);
   mult_28_C92_U931 : INVDL port map( A => mult_28_C92_n604, Z => 
                           mult_28_C92_net11981);
   mult_28_C92_U930 : INVD16 port map( A => data_in(5), Z => mult_28_C92_n1042)
                           ;
   mult_28_C92_U929 : NAN3D1 port map( A1 => mult_28_C92_n976, A2 => 
                           mult_28_C92_n977, A3 => mult_28_C92_n978, Z => 
                           mult_28_C92_n373);
   mult_28_C92_U928 : NAN2DL port map( A1 => mult_28_C92_n378, A2 => 
                           mult_28_C92_n376, Z => mult_28_C92_n978);
   mult_28_C92_U927 : NAN2DL port map( A1 => mult_28_C92_n387, A2 => 
                           mult_28_C92_n376, Z => mult_28_C92_n977);
   mult_28_C92_U926 : NAN2DL port map( A1 => mult_28_C92_n387, A2 => 
                           mult_28_C92_n378, Z => mult_28_C92_n976);
   mult_28_C92_U925 : NAN3D2 port map( A1 => mult_28_C92_n973, A2 => 
                           mult_28_C92_n974, A3 => mult_28_C92_n975, Z => 
                           mult_28_C92_n375);
   mult_28_C92_U924 : NAN2D1 port map( A1 => mult_28_C92_n380, A2 => 
                           mult_28_C92_n389, Z => mult_28_C92_n975);
   mult_28_C92_U923 : NAN2D1 port map( A1 => mult_28_C92_n391, A2 => 
                           mult_28_C92_n389, Z => mult_28_C92_n974);
   mult_28_C92_U922 : NAN2DL port map( A1 => mult_28_C92_n391, A2 => 
                           mult_28_C92_n380, Z => mult_28_C92_n973);
   mult_28_C92_U921 : EXOR2D1 port map( A1 => mult_28_C92_n972, A2 => 
                           mult_28_C92_n376, Z => mult_28_C92_n374);
   mult_28_C92_U920 : EXOR2D2 port map( A1 => mult_28_C92_n387, A2 => 
                           mult_28_C92_n378, Z => mult_28_C92_n972);
   mult_28_C92_U919 : EXOR3D1 port map( A1 => mult_28_C92_n391, A2 => 
                           mult_28_C92_n380, A3 => mult_28_C92_n389, Z => 
                           mult_28_C92_n376);
   mult_28_C92_U918 : NAN3D2 port map( A1 => mult_28_C92_n969, A2 => 
                           mult_28_C92_n971, A3 => mult_28_C92_n970, Z => 
                           mult_28_C92_n389);
   mult_28_C92_U917 : NAN2D1 port map( A1 => mult_28_C92_n396, A2 => 
                           mult_28_C92_n405, Z => mult_28_C92_n971);
   mult_28_C92_U916 : NAN2D1 port map( A1 => mult_28_C92_n394, A2 => 
                           mult_28_C92_n405, Z => mult_28_C92_n970);
   mult_28_C92_U915 : NAN2D1 port map( A1 => mult_28_C92_n394, A2 => 
                           mult_28_C92_n396, Z => mult_28_C92_n969);
   mult_28_C92_U914 : NAN2D1 port map( A1 => mult_28_C92_n429, A2 => 
                           mult_28_C92_n431, Z => mult_28_C92_n1120);
   mult_28_C92_U913 : INVD2 port map( A => mult_28_C92_n414, Z => 
                           mult_28_C92_n966);
   mult_28_C92_U912 : INVD2 port map( A => mult_28_C92_n1081, Z => 
                           mult_28_C92_n965);
   mult_28_C92_U911 : NAN2D2 port map( A1 => mult_28_C92_n967, A2 => 
                           mult_28_C92_n968, Z => mult_28_C92_n412);
   mult_28_C92_U910 : NAN2D2 port map( A1 => mult_28_C92_n965, A2 => 
                           mult_28_C92_n966, Z => mult_28_C92_n968);
   mult_28_C92_U909 : NAN2D1 port map( A1 => mult_28_C92_n1081, A2 => 
                           mult_28_C92_n414, Z => mult_28_C92_n967);
   mult_28_C92_U908 : INVD20 port map( A => data_in(11), Z => mult_28_C92_n993)
                           ;
   mult_28_C92_U907 : NAN2D2 port map( A1 => mult_28_C92_n993, A2 => 
                           mult_28_C92_net12088, Z => mult_28_C92_n995);
   mult_28_C92_U906 : NAN2D1 port map( A1 => mult_28_C92_n374, A2 => 
                           mult_28_C92_n385, Z => mult_28_C92_n180);
   mult_28_C92_U905 : NAN3D2 port map( A1 => mult_28_C92_n1048, A2 => 
                           mult_28_C92_n1050, A3 => mult_28_C92_n1049, Z => 
                           mult_28_C92_n417);
   mult_28_C92_U904 : OAI22D1 port map( A1 => mult_28_C92_n716, A2 => 
                           mult_28_C92_n30, B1 => mult_28_C92_n715, B2 => 
                           mult_28_C92_n28, Z => mult_28_C92_n584);
   mult_28_C92_U903 : INVD2 port map( A => data_in(9), Z => mult_28_C92_n962);
   mult_28_C92_U902 : NAN2D1 port map( A1 => mult_28_C92_n963, A2 => 
                           mult_28_C92_n964, Z => mult_28_C92_n716);
   mult_28_C92_U901 : NAN2D2 port map( A1 => mult_28_C92_n962, A2 => 
                           mult_28_C92_n1056, Z => mult_28_C92_n964);
   mult_28_C92_U900 : NAN2D1 port map( A1 => data_in(9), A2 => 
                           coeff_memory_73_port, Z => mult_28_C92_n963);
   mult_28_C92_U899 : OAI22DL port map( A1 => mult_28_C92_n765, A2 => 
                           mult_28_C92_n12, B1 => mult_28_C92_n764, B2 => 
                           mult_28_C92_n9, Z => mult_28_C92_n630);
   mult_28_C92_U898 : NAN2D2 port map( A1 => mult_28_C92_n960, A2 => 
                           mult_28_C92_n961, Z => mult_28_C92_n765);
   mult_28_C92_U897 : NAN2D2 port map( A1 => mult_28_C92_n993, A2 => 
                           mult_28_C92_net12160, Z => mult_28_C92_n961);
   mult_28_C92_U896 : NAN2D1 port map( A1 => data_in(11), A2 => 
                           coeff_memory_67_port, Z => mult_28_C92_n960);
   mult_28_C92_U895 : EXNOR2DL port map( A1 => data_in(2), A2 => 
                           coeff_memory_79_port, Z => mult_28_C92_n672);
   mult_28_C92_U894 : OAI22D1 port map( A1 => mult_28_C92_n672, A2 => 
                           mult_28_C92_n48, B1 => mult_28_C92_n671, B2 => 
                           mult_28_C92_n46, Z => mult_28_C92_n543);
   mult_28_C92_U893 : NAN2D2 port map( A1 => mult_28_C92_n1111, A2 => 
                           mult_28_C92_n1112, Z => mult_28_C92_n722);
   mult_28_C92_U892 : NAN2D2 port map( A1 => mult_28_C92_n1067, A2 => 
                           mult_28_C92_net12160, Z => mult_28_C92_n1068);
   mult_28_C92_U891 : INVD4 port map( A => data_in(1), Z => mult_28_C92_n957);
   mult_28_C92_U890 : NAN2D2 port map( A1 => mult_28_C92_n958, A2 => 
                           mult_28_C92_n959, Z => mult_28_C92_n690);
   mult_28_C92_U889 : NAN2D2 port map( A1 => mult_28_C92_n957, A2 => 
                           mult_28_C92_n1061, Z => mult_28_C92_n959);
   mult_28_C92_U888 : NAN2D1 port map( A1 => data_in(1), A2 => 
                           coeff_memory_77_port, Z => mult_28_C92_n958);
   mult_28_C92_U887 : NOR2DL port map( A1 => mult_28_C92_n202, A2 => 
                           mult_28_C92_n207, Z => mult_28_C92_n196);
   mult_28_C92_U886 : NOR2DL port map( A1 => mult_28_C92_n202, A2 => 
                           mult_28_C92_n207, Z => mult_28_C92_n956);
   mult_28_C92_U885 : NOR2DL port map( A1 => mult_28_C92_n202, A2 => 
                           mult_28_C92_n207, Z => mult_28_C92_n955);
   mult_28_C92_U884 : INVD2 port map( A => mult_28_C92_n1001, Z => 
                           mult_28_C92_n509);
   mult_28_C92_U883 : INVDL port map( A => mult_28_C92_n999, Z => 
                           mult_28_C92_n1028);
   mult_28_C92_U882 : NAN2DL port map( A1 => mult_28_C92_n426, A2 => 
                           mult_28_C92_n439, Z => mult_28_C92_n208);
   mult_28_C92_U881 : NAN2D1 port map( A1 => mult_28_C92_n1043, A2 => 
                           mult_28_C92_n1044, Z => mult_28_C92_n737);
   mult_28_C92_U880 : NAN3D2 port map( A1 => mult_28_C92_n951, A2 => 
                           mult_28_C92_n952, A3 => mult_28_C92_n953, Z => 
                           mult_28_C92_n443);
   mult_28_C92_U879 : NAN2D1 port map( A1 => mult_28_C92_n459, A2 => 
                           mult_28_C92_n450, Z => mult_28_C92_n953);
   mult_28_C92_U878 : NAN2D1 port map( A1 => mult_28_C92_n457, A2 => 
                           mult_28_C92_n450, Z => mult_28_C92_n952);
   mult_28_C92_U877 : NAN2DL port map( A1 => mult_28_C92_n457, A2 => 
                           mult_28_C92_n459, Z => mult_28_C92_n951);
   mult_28_C92_U876 : NAN3D2 port map( A1 => mult_28_C92_n948, A2 => 
                           mult_28_C92_n949, A3 => mult_28_C92_n950, Z => 
                           mult_28_C92_n449);
   mult_28_C92_U875 : NAN2D1 port map( A1 => mult_28_C92_n546, A2 => 
                           mult_28_C92_n645, Z => mult_28_C92_n950);
   mult_28_C92_U874 : NAN2D1 port map( A1 => mult_28_C92_n574, A2 => 
                           mult_28_C92_n645, Z => mult_28_C92_n949);
   mult_28_C92_U873 : NAN2D1 port map( A1 => mult_28_C92_n574, A2 => 
                           mult_28_C92_n546, Z => mult_28_C92_n948);
   mult_28_C92_U872 : EXOR2D1 port map( A1 => mult_28_C92_n457, A2 => 
                           mult_28_C92_n459, Z => mult_28_C92_n947);
   mult_28_C92_U871 : EXOR3D2 port map( A1 => mult_28_C92_n574, A2 => 
                           mult_28_C92_n546, A3 => mult_28_C92_n645, Z => 
                           mult_28_C92_n450);
   mult_28_C92_U870 : EXOR3D1 port map( A1 => mult_28_C92_n643, A2 => 
                           mult_28_C92_n544, A3 => mult_28_C92_n586, Z => 
                           mult_28_C92_n422);
   mult_28_C92_U869 : NAN3D1 port map( A1 => mult_28_C92_n944, A2 => 
                           mult_28_C92_n946, A3 => mult_28_C92_n945, Z => 
                           mult_28_C92_n415);
   mult_28_C92_U868 : NAN2D1 port map( A1 => mult_28_C92_n420, A2 => 
                           mult_28_C92_n433, Z => mult_28_C92_n946);
   mult_28_C92_U867 : NAN2DL port map( A1 => mult_28_C92_n422, A2 => 
                           mult_28_C92_n433, Z => mult_28_C92_n945);
   mult_28_C92_U866 : NAN2DL port map( A1 => mult_28_C92_n422, A2 => 
                           mult_28_C92_n420, Z => mult_28_C92_n944);
   mult_28_C92_U865 : NAN2D2 port map( A1 => mult_28_C92_n1072, A2 => 
                           mult_28_C92_net12088, Z => mult_28_C92_n1074);
   mult_28_C92_U864 : EXOR2D1 port map( A1 => mult_28_C92_n947, A2 => 
                           mult_28_C92_n450, Z => mult_28_C92_n444);
   mult_28_C92_U863 : EXNOR2D1 port map( A1 => data_in(4), A2 => 
                           coeff_memory_75_port, Z => mult_28_C92_n704);
   mult_28_C92_U862 : OAI22DL port map( A1 => mult_28_C92_n704, A2 => 
                           mult_28_C92_n36, B1 => mult_28_C92_n703, B2 => 
                           mult_28_C92_n34, Z => mult_28_C92_n573);
   mult_28_C92_U861 : EXNOR2D1 port map( A1 => data_in(8), A2 => 
                           coeff_memory_73_port, Z => mult_28_C92_n1092);
   mult_28_C92_U860 : OAI22D1 port map( A1 => mult_28_C92_n706, A2 => 
                           mult_28_C92_n36, B1 => mult_28_C92_n1080, B2 => 
                           mult_28_C92_n34, Z => mult_28_C92_n943);
   mult_28_C92_U859 : EXOR2D1 port map( A1 => mult_28_C92_n623, A2 => 
                           mult_28_C92_n527, Z => mult_28_C92_n510);
   mult_28_C92_U858 : EXNOR2D1 port map( A1 => data_in(12), A2 => 
                           coeff_memory_65_port, Z => mult_28_C92_n781);
   mult_28_C92_U857 : OA22DL port map( A1 => mult_28_C92_n660, A2 => 
                           mult_28_C92_n48, B1 => mult_28_C92_n659, B2 => 
                           mult_28_C92_n46, Z => mult_28_C92_n942);
   mult_28_C92_U856 : AND2DL port map( A1 => mult_28_C92_n290, A2 => 
                           mult_28_C92_n133, Z => mult_28_C92_n941);
   mult_28_C92_U855 : AND2DL port map( A1 => mult_28_C92_n911, A2 => 
                           mult_28_C92_n478, Z => mult_28_C92_n940);
   mult_28_C92_U854 : AND2D1 port map( A1 => mult_28_C92_n943, A2 => 
                           mult_28_C92_n524, Z => mult_28_C92_n939);
   mult_28_C92_U853 : INVDL port map( A => coeff_memory_67_port, Z => 
                           mult_28_C92_net12160);
   mult_28_C92_U852 : INVDL port map( A => coeff_memory_75_port, Z => 
                           mult_28_C92_net11946);
   mult_28_C92_U851 : INVD1 port map( A => coeff_memory_73_port, Z => 
                           mult_28_C92_n1056);
   mult_28_C92_U850 : INVD1 port map( A => coeff_memory_69_port, Z => 
                           mult_28_C92_net12088);
   mult_28_C92_U849 : NAN2DL port map( A1 => mult_28_C92_n294, A2 => 
                           mult_28_C92_n175, Z => mult_28_C92_n63);
   mult_28_C92_U848 : NOR2D1 port map( A1 => mult_28_C92_n332, A2 => 
                           mult_28_C92_n337, Z => mult_28_C92_n130);
   mult_28_C92_U847 : OAI22DL port map( A1 => mult_28_C92_n754, A2 => 
                           mult_28_C92_n18, B1 => mult_28_C92_n1104, B2 => 
                           mult_28_C92_n16, Z => mult_28_C92_n620);
   mult_28_C92_U846 : OAI22D1 port map( A1 => mult_28_C92_n1108, A2 => 
                           mult_28_C92_n18, B1 => mult_28_C92_n1105, B2 => 
                           mult_28_C92_n16, Z => mult_28_C92_n618);
   mult_28_C92_U845 : INVD1 port map( A => coeff_memory_64_port, Z => 
                           mult_28_C92_n834);
   mult_28_C92_U844 : NAN3D1 port map( A1 => mult_28_C92_n1096, A2 => 
                           mult_28_C92_n1098, A3 => mult_28_C92_n1097, Z => 
                           mult_28_C92_n405);
   mult_28_C92_U843 : INVD16 port map( A => data_in(3), Z => mult_28_C92_n1110)
                           ;
   mult_28_C92_U842 : NAN2D1 port map( A1 => mult_28_C92_n1087, A2 => 
                           mult_28_C92_n1088, Z => mult_28_C92_n752);
   mult_28_C92_U841 : OR2D1 port map( A1 => mult_28_C92_n752, A2 => 
                           mult_28_C92_n16, Z => mult_28_C92_n1141);
   mult_28_C92_U840 : INVD1 port map( A => mult_28_C92_n842, Z => 
                           mult_28_C92_n1075);
   mult_28_C92_U839 : NAN2DL port map( A1 => data_in(11), A2 => 
                           coeff_memory_69_port, Z => mult_28_C92_n994);
   mult_28_C92_U838 : EXOR2D1 port map( A1 => mult_28_C92_n57, A2 => 
                           mult_28_C92_n114, Z => m1_12);
   mult_28_C92_U837 : INVDL port map( A => mult_28_C92_n125, Z => 
                           mult_28_C92_n289);
   mult_28_C92_U836 : NOR2DL port map( A1 => mult_28_C92_n170, A2 => 
                           mult_28_C92_n161, Z => mult_28_C92_n159);
   mult_28_C92_U835 : NAN2D2 port map( A1 => mult_28_C92_n1078, A2 => 
                           mult_28_C92_n1079, Z => mult_28_C92_n1113);
   mult_28_C92_U834 : INVD16 port map( A => data_in(10), Z => mult_28_C92_n986)
                           ;
   mult_28_C92_U833 : EXNOR2DL port map( A1 => data_in(10), A2 => 
                           coeff_memory_69_port, Z => mult_28_C92_n749);
   mult_28_C92_U832 : EXNOR2DL port map( A1 => data_in(10), A2 => 
                           coeff_memory_79_port, Z => mult_28_C92_n664);
   mult_28_C92_U831 : INVD1 port map( A => mult_28_C92_n1075, Z => 
                           mult_28_C92_n936);
   mult_28_C92_U830 : INVD1 port map( A => data_in(10), Z => mult_28_C92_n935);
   mult_28_C92_U829 : NAN2D1 port map( A1 => mult_28_C92_n937, A2 => 
                           mult_28_C92_n938, Z => mult_28_C92_n783);
   mult_28_C92_U828 : NAN2D1 port map( A1 => mult_28_C92_n935, A2 => 
                           mult_28_C92_n936, Z => mult_28_C92_n938);
   mult_28_C92_U827 : NAN2D1 port map( A1 => data_in(10), A2 => 
                           mult_28_C92_n1075, Z => mult_28_C92_n937);
   mult_28_C92_U826 : INVD2 port map( A => data_in(9), Z => 
                           mult_28_C92_net11996);
   mult_28_C92_U825 : OAI21D1 port map( A1 => mult_28_C92_n141, A2 => 
                           mult_28_C92_n162, B => mult_28_C92_n142, Z => 
                           mult_28_C92_n140);
   mult_28_C92_U824 : INVD2 port map( A => mult_28_C92_n430, Z => 
                           mult_28_C92_n1077);
   mult_28_C92_U823 : NOR2D1 port map( A1 => mult_28_C92_n386, A2 => 
                           mult_28_C92_n397, Z => mult_28_C92_n186);
   mult_28_C92_U822 : EXOR3D1 port map( A1 => mult_28_C92_n405, A2 => 
                           mult_28_C92_n394, A3 => mult_28_C92_n396, Z => 
                           mult_28_C92_n390);
   mult_28_C92_U821 : NAN3D1 port map( A1 => mult_28_C92_n932, A2 => 
                           mult_28_C92_n934, A3 => mult_28_C92_n933, Z => 
                           mult_28_C92_n385);
   mult_28_C92_U820 : NAN2DL port map( A1 => mult_28_C92_n388, A2 => 
                           mult_28_C92_n390, Z => mult_28_C92_n934);
   mult_28_C92_U819 : NAN2DL port map( A1 => mult_28_C92_n399, A2 => 
                           mult_28_C92_n390, Z => mult_28_C92_n933);
   mult_28_C92_U818 : NAN2DL port map( A1 => mult_28_C92_n399, A2 => 
                           mult_28_C92_n388, Z => mult_28_C92_n932);
   mult_28_C92_U817 : EXOR3D1 port map( A1 => mult_28_C92_n399, A2 => 
                           mult_28_C92_n390, A3 => mult_28_C92_n388, Z => 
                           mult_28_C92_n386);
   mult_28_C92_U816 : INVDL port map( A => mult_28_C92_net12187, Z => 
                           mult_28_C92_n1002);
   mult_28_C92_U815 : AOI21D1 port map( A1 => mult_28_C92_n169, A2 => 
                           mult_28_C92_n139, B => mult_28_C92_n140, Z => 
                           mult_28_C92_n1064);
   mult_28_C92_U814 : AND2D1 port map( A1 => mult_28_C92_n464, A2 => 
                           mult_28_C92_n473, Z => mult_28_C92_net12350);
   mult_28_C92_U813 : EXNOR2DL port map( A1 => data_in(15), A2 => 
                           coeff_memory_65_port, Z => mult_28_C92_n931);
   mult_28_C92_U812 : INVD1 port map( A => mult_28_C92_n221, Z => 
                           mult_28_C92_n219);
   mult_28_C92_U811 : INVDL port map( A => coeff_memory_71_port, Z => 
                           mult_28_C92_n928);
   mult_28_C92_U810 : INVD1 port map( A => data_in(6), Z => mult_28_C92_n927);
   mult_28_C92_U809 : NAN2D1 port map( A1 => mult_28_C92_n929, A2 => 
                           mult_28_C92_n930, Z => mult_28_C92_n1016);
   mult_28_C92_U808 : NAN2D1 port map( A1 => mult_28_C92_n927, A2 => 
                           mult_28_C92_n928, Z => mult_28_C92_n930);
   mult_28_C92_U807 : NAN2DL port map( A1 => data_in(6), A2 => 
                           coeff_memory_71_port, Z => mult_28_C92_n929);
   mult_28_C92_U806 : INVD1 port map( A => mult_28_C92_n197, Z => 
                           mult_28_C92_n199);
   mult_28_C92_U805 : INVD1 port map( A => mult_28_C92_n199, Z => 
                           mult_28_C92_n926);
   mult_28_C92_U804 : NOR2D1 port map( A1 => mult_28_C92_n426, A2 => 
                           mult_28_C92_n439, Z => mult_28_C92_n207);
   mult_28_C92_U803 : NAN2D1 port map( A1 => mult_28_C92_n426, A2 => 
                           mult_28_C92_n439, Z => mult_28_C92_n954);
   mult_28_C92_U802 : INVDL port map( A => mult_28_C92_n428, Z => 
                           mult_28_C92_n923);
   mult_28_C92_U801 : INVD2 port map( A => mult_28_C92_n1113, Z => 
                           mult_28_C92_n922);
   mult_28_C92_U800 : NAN2D2 port map( A1 => mult_28_C92_n924, A2 => 
                           mult_28_C92_n925, Z => mult_28_C92_n426);
   mult_28_C92_U799 : NAN2D1 port map( A1 => mult_28_C92_n922, A2 => 
                           mult_28_C92_n428, Z => mult_28_C92_n925);
   mult_28_C92_U798 : NAN2D1 port map( A1 => mult_28_C92_n1113, A2 => 
                           mult_28_C92_n923, Z => mult_28_C92_n924);
   mult_28_C92_U797 : EXNOR2D1 port map( A1 => data_in(10), A2 => 
                           coeff_memory_67_port, Z => mult_28_C92_n1030);
   mult_28_C92_U796 : INVDL port map( A => coeff_memory_77_port, Z => 
                           mult_28_C92_n919);
   mult_28_C92_U795 : INVD2 port map( A => data_in(3), Z => mult_28_C92_n918);
   mult_28_C92_U794 : NAN2D2 port map( A1 => mult_28_C92_n920, A2 => 
                           mult_28_C92_n921, Z => mult_28_C92_n688);
   mult_28_C92_U793 : NAN2D2 port map( A1 => mult_28_C92_n918, A2 => 
                           mult_28_C92_n919, Z => mult_28_C92_n921);
   mult_28_C92_U792 : NAN2D1 port map( A1 => data_in(3), A2 => 
                           coeff_memory_77_port, Z => mult_28_C92_n920);
   mult_28_C92_U791 : NAN2D1 port map( A1 => mult_28_C92_n424, A2 => 
                           mult_28_C92_n435, Z => mult_28_C92_n1048);
   mult_28_C92_U790 : EXNOR2D1 port map( A1 => data_in(2), A2 => 
                           coeff_memory_73_port, Z => mult_28_C92_n917);
   mult_28_C92_U789 : EXNOR2DL port map( A1 => data_in(6), A2 => 
                           coeff_memory_71_port, Z => mult_28_C92_n916);
   mult_28_C92_U788 : NAN2D2 port map( A1 => mult_28_C92_n1073, A2 => 
                           mult_28_C92_n1074, Z => mult_28_C92_n751);
   mult_28_C92_U787 : EXOR3D2 port map( A1 => mult_28_C92_n465, A2 => 
                           mult_28_C92_n456, A3 => mult_28_C92_n454, Z => 
                           mult_28_C92_net11792);
   mult_28_C92_U786 : EXOR3D2 port map( A1 => mult_28_C92_n433, A2 => 
                           mult_28_C92_n422, A3 => mult_28_C92_n420, Z => 
                           mult_28_C92_n416);
   mult_28_C92_U785 : INVDL port map( A => mult_28_C92_n416, Z => 
                           mult_28_C92_n913);
   mult_28_C92_U784 : INVD1 port map( A => mult_28_C92_n427, Z => 
                           mult_28_C92_n912);
   mult_28_C92_U783 : NAN2D2 port map( A1 => mult_28_C92_n914, A2 => 
                           mult_28_C92_n915, Z => mult_28_C92_n1081);
   mult_28_C92_U782 : NAN2D2 port map( A1 => mult_28_C92_n912, A2 => 
                           mult_28_C92_n913, Z => mult_28_C92_n915);
   mult_28_C92_U781 : NAN2D1 port map( A1 => mult_28_C92_n427, A2 => 
                           mult_28_C92_n416, Z => mult_28_C92_n914);
   mult_28_C92_U780 : EXOR3D2 port map( A1 => mult_28_C92_n437, A2 => 
                           mult_28_C92_n424, A3 => mult_28_C92_n435, Z => 
                           mult_28_C92_n418);
   mult_28_C92_U779 : NAN2DL port map( A1 => mult_28_C92_n472, A2 => 
                           mult_28_C92_n477, Z => mult_28_C92_net9969);
   mult_28_C92_U778 : INVDL port map( A => mult_28_C92_n910, Z => 
                           mult_28_C92_n911);
   mult_28_C92_U777 : INVDL port map( A => mult_28_C92_n485, Z => 
                           mult_28_C92_n910);
   mult_28_C92_U237 : AOI21D1 port map( A1 => mult_28_C92_n218, A2 => 
                           mult_28_C92_net12350, B => mult_28_C92_n219, Z => 
                           mult_28_C92_n217);
   mult_28_C92_U599 : OAI22D1 port map( A1 => mult_28_C92_n737, A2 => 
                           mult_28_C92_n24, B1 => mult_28_C92_n1016, B2 => 
                           mult_28_C92_n22, Z => mult_28_C92_n604);
   mult_28_C92_U426 : ADFULD1 port map( A => mult_28_C92_n605, B => 
                           mult_28_C92_n633, CI => mult_28_C92_n482, CO => 
                           mult_28_C92_n477, S => mult_28_C92_n478);
   mult_28_C92_U428 : ADHALFD1 port map( A => mult_28_C92_n525, B => 
                           mult_28_C92_n591, CO => mult_28_C92_n481, S => 
                           mult_28_C92_n482);
   mult_28_C92_U518 : OAI22D1 port map( A1 => mult_28_C92_n36, A2 => 
                           mult_28_C92_net11946, B1 => mult_28_C92_n709, B2 => 
                           mult_28_C92_n34, Z => mult_28_C92_n525);
   mult_28_C92_U552 : NAN2M1D1 port map( A1 => data_in(0), A2 => 
                           coeff_memory_75_port, Z => mult_28_C92_n709);
   mult_28_C92_U218 : AOI21D1 port map( A1 => mult_28_C92_n299, A2 => 
                           mult_28_C92_net12275, B => mult_28_C92_n206, Z => 
                           mult_28_C92_n204);
   mult_28_C92_U429 : ADFULD1 port map( A => mult_28_C92_n493, B => 
                           mult_28_C92_n488, CI => mult_28_C92_n486, CO => 
                           mult_28_C92_n483, S => mult_28_C92_n484);
   mult_28_C92_U263 : NOR2D2 port map( A1 => mult_28_C92_n474, A2 => 
                           mult_28_C92_n483, Z => mult_28_C92_n235);
   mult_28_C92_U275 : AOI21D1 port map( A1 => mult_28_C92_n248, A2 => 
                           mult_28_C92_n1021, B => mult_28_C92_n1020, Z => 
                           mult_28_C92_n243);
   mult_28_C92_U285 : AOI21D1 port map( A1 => mult_28_C92_net11021, A2 => 
                           mult_28_C92_n1024, B => mult_28_C92_n1022, Z => 
                           mult_28_C92_n250);
   mult_28_C92_U302 : AOI21D1 port map( A1 => mult_28_C92_net10923, A2 => 
                           mult_28_C92_n266, B => mult_28_C92_n1019, Z => 
                           mult_28_C92_n261);
   mult_28_C92_U310 : OAI21D1 port map( A1 => mult_28_C92_n267, A2 => 
                           mult_28_C92_n269, B => mult_28_C92_n268, Z => 
                           mult_28_C92_n266);
   mult_28_C92_U316 : AOI21D1 port map( A1 => mult_28_C92_net10919, A2 => 
                           mult_28_C92_n274, B => mult_28_C92_n1018, Z => 
                           mult_28_C92_n269);
   mult_28_C92_U665 : OAI22D1 port map( A1 => mult_28_C92_n767, A2 => 
                           mult_28_C92_n12, B1 => mult_28_C92_n1030, B2 => 
                           mult_28_C92_n9, Z => mult_28_C92_n632);
   mult_28_C92_U534 : OAI22D1 port map( A1 => mult_28_C92_n708, A2 => 
                           mult_28_C92_n36, B1 => mult_28_C92_n707, B2 => 
                           mult_28_C92_n34, Z => mult_28_C92_n577);
   mult_28_C92_U172 : OAI21D1 port map( A1 => mult_28_C92_n174, A2 => 
                           mult_28_C92_n180, B => mult_28_C92_n175, Z => 
                           mult_28_C92_n169);
   mult_28_C92_U188 : AOI21D1 port map( A1 => mult_28_C92_n197, A2 => 
                           mult_28_C92_n1033, B => mult_28_C92_n185, Z => 
                           mult_28_C92_n183);
   mult_28_C92_U232 : NOR2D2 port map( A1 => mult_28_C92_n440, A2 => 
                           mult_28_C92_n451, Z => mult_28_C92_n213);
   mult_28_C92_U415 : ADFULD1 port map( A => mult_28_C92_n462, B => 
                           mult_28_C92_n471, CI => mult_28_C92_n469, CO => 
                           mult_28_C92_n455, S => mult_28_C92_n456);
   mult_28_C92_U212 : OAI21D1 port map( A1 => mult_28_C92_n208, A2 => 
                           mult_28_C92_n202, B => mult_28_C92_n203, Z => 
                           mult_28_C92_n197);
   mult_28_C92_U203 : NOR2D2 port map( A1 => mult_28_C92_n398, A2 => 
                           mult_28_C92_n411, Z => mult_28_C92_n191);
   mult_28_C92_U761 : EXOR2D1 port map( A1 => coeff_memory_73_port, A2 => 
                           coeff_memory_72_port, Z => mult_28_C92_n814);
   mult_28_C92_U755 : EXOR2D1 port map( A1 => coeff_memory_77_port, A2 => 
                           coeff_memory_76_port, Z => mult_28_C92_n812);
   mult_28_C92_U752 : EXOR2D1 port map( A1 => coeff_memory_78_port, A2 => 
                           coeff_memory_79_port, Z => mult_28_C92_n811);
   mult_28_C92_U727 : NAN2M1D1 port map( A1 => data_in(0), A2 => 
                           coeff_memory_65_port, Z => mult_28_C92_n794);
   mult_28_C92_U726 : EXNOR2D1 port map( A1 => data_in(0), A2 => 
                           coeff_memory_65_port, Z => mult_28_C92_n793);
   mult_28_C92_U725 : EXNOR2D1 port map( A1 => data_in(1), A2 => 
                           coeff_memory_65_port, Z => mult_28_C92_n792);
   mult_28_C92_U724 : EXNOR2D1 port map( A1 => data_in(2), A2 => 
                           coeff_memory_65_port, Z => mult_28_C92_n791);
   mult_28_C92_U723 : EXNOR2D1 port map( A1 => data_in(3), A2 => 
                           coeff_memory_65_port, Z => mult_28_C92_n790);
   mult_28_C92_U722 : EXNOR2D1 port map( A1 => data_in(4), A2 => 
                           coeff_memory_65_port, Z => mult_28_C92_n789);
   mult_28_C92_U721 : EXNOR2D1 port map( A1 => data_in(5), A2 => 
                           coeff_memory_65_port, Z => mult_28_C92_n788);
   mult_28_C92_U720 : EXNOR2D1 port map( A1 => data_in(6), A2 => 
                           coeff_memory_65_port, Z => mult_28_C92_n787);
   mult_28_C92_U718 : EXNOR2D1 port map( A1 => data_in(8), A2 => 
                           coeff_memory_65_port, Z => mult_28_C92_n785);
   mult_28_C92_U713 : EXNOR2D1 port map( A1 => data_in(13), A2 => 
                           coeff_memory_65_port, Z => mult_28_C92_n780);
   mult_28_C92_U711 : EXNOR2D1 port map( A1 => data_in(15), A2 => 
                           coeff_memory_65_port, Z => mult_28_C92_n778);
   mult_28_C92_U708 : OAI22D1 port map( A1 => mult_28_C92_n792, A2 => 
                           mult_28_C92_n6, B1 => mult_28_C92_n791, B2 => 
                           mult_28_C92_n834, Z => mult_28_C92_n657);
   mult_28_C92_U706 : OAI22D1 port map( A1 => mult_28_C92_n790, A2 => 
                           mult_28_C92_n6, B1 => mult_28_C92_n789, B2 => 
                           mult_28_C92_n834, Z => mult_28_C92_n655);
   mult_28_C92_U704 : OAI22D1 port map( A1 => mult_28_C92_n788, A2 => 
                           mult_28_C92_n6, B1 => mult_28_C92_n787, B2 => 
                           mult_28_C92_n834, Z => mult_28_C92_n653);
   mult_28_C92_U703 : OAI22D1 port map( A1 => mult_28_C92_n787, A2 => 
                           mult_28_C92_n6, B1 => mult_28_C92_n786, B2 => 
                           mult_28_C92_n834, Z => mult_28_C92_n652);
   mult_28_C92_U702 : OAI22D1 port map( A1 => mult_28_C92_n786, A2 => 
                           mult_28_C92_n6, B1 => mult_28_C92_n785, B2 => 
                           mult_28_C92_n834, Z => mult_28_C92_n651);
   mult_28_C92_U699 : OAI22D1 port map( A1 => mult_28_C92_n783, A2 => 
                           mult_28_C92_n6, B1 => mult_28_C92_n782, B2 => 
                           mult_28_C92_n834, Z => mult_28_C92_n648);
   mult_28_C92_U698 : OAI22D1 port map( A1 => mult_28_C92_n1107, A2 => 
                           mult_28_C92_n6, B1 => mult_28_C92_n781, B2 => 
                           mult_28_C92_n834, Z => mult_28_C92_n647);
   mult_28_C92_U696 : OAI22D1 port map( A1 => mult_28_C92_n780, A2 => 
                           mult_28_C92_n6, B1 => mult_28_C92_n1082, B2 => 
                           mult_28_C92_n834, Z => mult_28_C92_n645);
   mult_28_C92_U695 : OAI22D1 port map( A1 => mult_28_C92_n779, A2 => 
                           mult_28_C92_n6, B1 => mult_28_C92_n931, B2 => 
                           mult_28_C92_n834, Z => mult_28_C92_n644);
   mult_28_C92_U694 : AO21D2 port map( A1 => mult_28_C92_n6, A2 => 
                           mult_28_C92_n834, B => mult_28_C92_n778, Z => 
                           mult_28_C92_n643);
   mult_28_C92_U693 : OAI22D1 port map( A1 => mult_28_C92_n6, A2 => 
                           mult_28_C92_n842, B1 => mult_28_C92_n794, B2 => 
                           mult_28_C92_n834, Z => mult_28_C92_n530);
   mult_28_C92_U692 : NAN2M1D1 port map( A1 => data_in(0), A2 => 
                           coeff_memory_67_port, Z => mult_28_C92_n777);
   mult_28_C92_U691 : EXNOR2D1 port map( A1 => data_in(0), A2 => 
                           coeff_memory_67_port, Z => mult_28_C92_n776);
   mult_28_C92_U690 : EXNOR2D1 port map( A1 => data_in(1), A2 => 
                           coeff_memory_67_port, Z => mult_28_C92_n775);
   mult_28_C92_U689 : EXNOR2D1 port map( A1 => data_in(2), A2 => 
                           coeff_memory_67_port, Z => mult_28_C92_n774);
   mult_28_C92_U688 : EXNOR2D1 port map( A1 => data_in(3), A2 => 
                           coeff_memory_67_port, Z => mult_28_C92_n773);
   mult_28_C92_U687 : EXNOR2D1 port map( A1 => data_in(4), A2 => 
                           coeff_memory_67_port, Z => mult_28_C92_n772);
   mult_28_C92_U686 : EXNOR2D1 port map( A1 => data_in(5), A2 => 
                           coeff_memory_67_port, Z => mult_28_C92_n771);
   mult_28_C92_U685 : EXNOR2D1 port map( A1 => data_in(6), A2 => 
                           coeff_memory_67_port, Z => mult_28_C92_n770);
   mult_28_C92_U683 : EXNOR2D1 port map( A1 => data_in(8), A2 => 
                           coeff_memory_67_port, Z => mult_28_C92_n768);
   mult_28_C92_U679 : EXNOR2D1 port map( A1 => data_in(12), A2 => 
                           coeff_memory_67_port, Z => mult_28_C92_n764);
   mult_28_C92_U676 : EXNOR2D1 port map( A1 => data_in(15), A2 => 
                           coeff_memory_67_port, Z => mult_28_C92_n761);
   mult_28_C92_U675 : NOR2M1D1 port map( A1 => data_in(0), A2 => mult_28_C92_n9
                           , Z => mult_28_C92_n642);
   mult_28_C92_U674 : OAI22D1 port map( A1 => mult_28_C92_n776, A2 => 
                           mult_28_C92_n12, B1 => mult_28_C92_n775, B2 => 
                           mult_28_C92_n9, Z => mult_28_C92_n641);
   mult_28_C92_U673 : OAI22D1 port map( A1 => mult_28_C92_n775, A2 => 
                           mult_28_C92_n12, B1 => mult_28_C92_n774, B2 => 
                           mult_28_C92_n9, Z => mult_28_C92_n640);
   mult_28_C92_U672 : OAI22D1 port map( A1 => mult_28_C92_n774, A2 => 
                           mult_28_C92_n12, B1 => mult_28_C92_n773, B2 => 
                           mult_28_C92_n9, Z => mult_28_C92_n639);
   mult_28_C92_U671 : OAI22D1 port map( A1 => mult_28_C92_n773, A2 => 
                           mult_28_C92_n12, B1 => mult_28_C92_n772, B2 => 
                           mult_28_C92_n9, Z => mult_28_C92_n638);
   mult_28_C92_U670 : OAI22D1 port map( A1 => mult_28_C92_n772, A2 => 
                           mult_28_C92_n12, B1 => mult_28_C92_n771, B2 => 
                           mult_28_C92_n9, Z => mult_28_C92_n637);
   mult_28_C92_U669 : OAI22D1 port map( A1 => mult_28_C92_n771, A2 => 
                           mult_28_C92_n12, B1 => mult_28_C92_n770, B2 => 
                           mult_28_C92_n9, Z => mult_28_C92_n636);
   mult_28_C92_U668 : OAI22D1 port map( A1 => mult_28_C92_n770, A2 => 
                           mult_28_C92_n12, B1 => mult_28_C92_n769, B2 => 
                           mult_28_C92_n9, Z => mult_28_C92_n635);
   mult_28_C92_U667 : OAI22D1 port map( A1 => mult_28_C92_n769, A2 => 
                           mult_28_C92_n12, B1 => mult_28_C92_n768, B2 => 
                           mult_28_C92_n9, Z => mult_28_C92_n634);
   mult_28_C92_U664 : OAI22D1 port map( A1 => mult_28_C92_n766, A2 => 
                           mult_28_C92_n12, B1 => mult_28_C92_n765, B2 => 
                           mult_28_C92_n9, Z => mult_28_C92_n631);
   mult_28_C92_U661 : OAI22D1 port map( A1 => mult_28_C92_n763, A2 => 
                           mult_28_C92_n12, B1 => mult_28_C92_n762, B2 => 
                           mult_28_C92_n9, Z => mult_28_C92_n628);
   mult_28_C92_U660 : OAI22D1 port map( A1 => mult_28_C92_n762, A2 => 
                           mult_28_C92_n12, B1 => mult_28_C92_n761, B2 => 
                           mult_28_C92_n9, Z => mult_28_C92_n409);
   mult_28_C92_U658 : OAI22D1 port map( A1 => mult_28_C92_n12, A2 => 
                           mult_28_C92_net12160, B1 => mult_28_C92_n777, B2 => 
                           mult_28_C92_n9, Z => mult_28_C92_n529);
   mult_28_C92_U657 : NAN2M1D1 port map( A1 => data_in(0), A2 => 
                           coeff_memory_69_port, Z => mult_28_C92_n760);
   mult_28_C92_U656 : EXNOR2D1 port map( A1 => data_in(0), A2 => 
                           coeff_memory_69_port, Z => mult_28_C92_n759);
   mult_28_C92_U653 : EXNOR2D1 port map( A1 => data_in(3), A2 => 
                           coeff_memory_69_port, Z => mult_28_C92_n756);
   mult_28_C92_U643 : EXNOR2D1 port map( A1 => data_in(13), A2 => 
                           coeff_memory_69_port, Z => mult_28_C92_n746);
   mult_28_C92_U642 : EXNOR2D1 port map( A1 => data_in(14), A2 => 
                           coeff_memory_69_port, Z => mult_28_C92_n745);
   mult_28_C92_U641 : EXNOR2D1 port map( A1 => data_in(15), A2 => 
                           coeff_memory_69_port, Z => mult_28_C92_n744);
   mult_28_C92_U640 : NOR2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C92_n16, Z => mult_28_C92_n626);
   mult_28_C92_U639 : OAI22D1 port map( A1 => mult_28_C92_n759, A2 => 
                           mult_28_C92_n18, B1 => mult_28_C92_n758, B2 => 
                           mult_28_C92_n16, Z => mult_28_C92_n625);
   mult_28_C92_U637 : OAI22D1 port map( A1 => mult_28_C92_n757, A2 => 
                           mult_28_C92_n18, B1 => mult_28_C92_n756, B2 => 
                           mult_28_C92_n16, Z => mult_28_C92_n623);
   mult_28_C92_U636 : OAI22D1 port map( A1 => mult_28_C92_n756, A2 => 
                           mult_28_C92_n18, B1 => mult_28_C92_n755, B2 => 
                           mult_28_C92_n16, Z => mult_28_C92_n622);
   mult_28_C92_U635 : OAI22D1 port map( A1 => mult_28_C92_n755, A2 => 
                           mult_28_C92_n18, B1 => mult_28_C92_n754, B2 => 
                           mult_28_C92_n16, Z => mult_28_C92_n621);
   mult_28_C92_U631 : OAI22D1 port map( A1 => mult_28_C92_n751, A2 => 
                           mult_28_C92_n18, B1 => mult_28_C92_n750, B2 => 
                           mult_28_C92_n16, Z => mult_28_C92_n617);
   mult_28_C92_U629 : OAI22D1 port map( A1 => mult_28_C92_n749, A2 => 
                           mult_28_C92_n18, B1 => mult_28_C92_n1090, B2 => 
                           mult_28_C92_n16, Z => mult_28_C92_n615);
   mult_28_C92_U628 : OAI22D1 port map( A1 => mult_28_C92_n748, A2 => 
                           mult_28_C92_n18, B1 => mult_28_C92_n747, B2 => 
                           mult_28_C92_n16, Z => mult_28_C92_n614);
   mult_28_C92_U627 : OAI22D1 port map( A1 => mult_28_C92_n747, A2 => 
                           mult_28_C92_n18, B1 => mult_28_C92_n746, B2 => 
                           mult_28_C92_n16, Z => mult_28_C92_n613);
   mult_28_C92_U626 : OAI22D1 port map( A1 => mult_28_C92_n746, A2 => 
                           mult_28_C92_n18, B1 => mult_28_C92_n745, B2 => 
                           mult_28_C92_n16, Z => mult_28_C92_n612);
   mult_28_C92_U625 : OAI22D1 port map( A1 => mult_28_C92_n745, A2 => 
                           mult_28_C92_n18, B1 => mult_28_C92_n744, B2 => 
                           mult_28_C92_n16, Z => mult_28_C92_n383);
   mult_28_C92_U623 : OAI22D1 port map( A1 => mult_28_C92_n18, A2 => 
                           mult_28_C92_net12088, B1 => mult_28_C92_n760, B2 => 
                           mult_28_C92_n16, Z => mult_28_C92_n528);
   mult_28_C92_U622 : NAN2M1D1 port map( A1 => data_in(0), A2 => 
                           coeff_memory_71_port, Z => mult_28_C92_n743);
   mult_28_C92_U621 : EXNOR2D1 port map( A1 => data_in(0), A2 => 
                           coeff_memory_71_port, Z => mult_28_C92_n742);
   mult_28_C92_U620 : EXNOR2D1 port map( A1 => data_in(1), A2 => 
                           coeff_memory_71_port, Z => mult_28_C92_n741);
   mult_28_C92_U619 : EXNOR2D1 port map( A1 => data_in(2), A2 => 
                           coeff_memory_71_port, Z => mult_28_C92_n740);
   mult_28_C92_U618 : EXNOR2D1 port map( A1 => data_in(3), A2 => 
                           coeff_memory_71_port, Z => mult_28_C92_n739);
   mult_28_C92_U617 : EXNOR2D1 port map( A1 => data_in(4), A2 => 
                           coeff_memory_71_port, Z => mult_28_C92_n738);
   mult_28_C92_U613 : EXNOR2D1 port map( A1 => data_in(8), A2 => 
                           coeff_memory_71_port, Z => mult_28_C92_n734);
   mult_28_C92_U610 : EXNOR2D1 port map( A1 => data_in(11), A2 => 
                           coeff_memory_71_port, Z => mult_28_C92_n731);
   mult_28_C92_U609 : EXNOR2D1 port map( A1 => data_in(12), A2 => 
                           coeff_memory_71_port, Z => mult_28_C92_n730);
   mult_28_C92_U608 : EXNOR2D1 port map( A1 => data_in(13), A2 => 
                           coeff_memory_71_port, Z => mult_28_C92_n729);
   mult_28_C92_U607 : EXNOR2D1 port map( A1 => data_in(14), A2 => 
                           coeff_memory_71_port, Z => mult_28_C92_n728);
   mult_28_C92_U606 : EXNOR2D1 port map( A1 => data_in(15), A2 => 
                           coeff_memory_71_port, Z => mult_28_C92_n727);
   mult_28_C92_U605 : NOR2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C92_n22, Z => mult_28_C92_n610);
   mult_28_C92_U604 : OAI22D1 port map( A1 => mult_28_C92_n742, A2 => 
                           mult_28_C92_n24, B1 => mult_28_C92_n741, B2 => 
                           mult_28_C92_n22, Z => mult_28_C92_n609);
   mult_28_C92_U603 : OAI22D1 port map( A1 => mult_28_C92_n741, A2 => 
                           mult_28_C92_n24, B1 => mult_28_C92_n740, B2 => 
                           mult_28_C92_n22, Z => mult_28_C92_n608);
   mult_28_C92_U601 : OAI22D1 port map( A1 => mult_28_C92_n739, A2 => 
                           mult_28_C92_n24, B1 => mult_28_C92_n738, B2 => 
                           mult_28_C92_n22, Z => mult_28_C92_n606);
   mult_28_C92_U598 : OAI22D1 port map( A1 => mult_28_C92_n736, A2 => 
                           mult_28_C92_n24, B1 => mult_28_C92_n735, B2 => 
                           mult_28_C92_n22, Z => mult_28_C92_n603);
   mult_28_C92_U597 : OAI22D1 port map( A1 => mult_28_C92_n735, A2 => 
                           mult_28_C92_n24, B1 => mult_28_C92_n734, B2 => 
                           mult_28_C92_n22, Z => mult_28_C92_n602);
   mult_28_C92_U596 : OAI22D1 port map( A1 => mult_28_C92_n734, A2 => 
                           mult_28_C92_n24, B1 => mult_28_C92_n733, B2 => 
                           mult_28_C92_n22, Z => mult_28_C92_n601);
   mult_28_C92_U595 : OAI22D1 port map( A1 => mult_28_C92_n733, A2 => 
                           mult_28_C92_n24, B1 => mult_28_C92_n732, B2 => 
                           mult_28_C92_n22, Z => mult_28_C92_n600);
   mult_28_C92_U594 : OAI22D1 port map( A1 => mult_28_C92_n732, A2 => 
                           mult_28_C92_n24, B1 => mult_28_C92_n731, B2 => 
                           mult_28_C92_n22, Z => mult_28_C92_n599);
   mult_28_C92_U593 : OAI22D1 port map( A1 => mult_28_C92_n731, A2 => 
                           mult_28_C92_n24, B1 => mult_28_C92_n730, B2 => 
                           mult_28_C92_n22, Z => mult_28_C92_n598);
   mult_28_C92_U592 : OAI22D1 port map( A1 => mult_28_C92_n730, A2 => 
                           mult_28_C92_n24, B1 => mult_28_C92_n729, B2 => 
                           mult_28_C92_n22, Z => mult_28_C92_n597);
   mult_28_C92_U591 : OAI22D1 port map( A1 => mult_28_C92_n729, A2 => 
                           mult_28_C92_n24, B1 => mult_28_C92_n728, B2 => 
                           mult_28_C92_n22, Z => mult_28_C92_n596);
   mult_28_C92_U590 : OAI22D1 port map( A1 => mult_28_C92_n728, A2 => 
                           mult_28_C92_n24, B1 => mult_28_C92_n727, B2 => 
                           mult_28_C92_n22, Z => mult_28_C92_n361);
   mult_28_C92_U588 : OAI22D1 port map( A1 => mult_28_C92_n24, A2 => 
                           mult_28_C92_net11920, B1 => mult_28_C92_n743, B2 => 
                           mult_28_C92_n22, Z => mult_28_C92_n527);
   mult_28_C92_U587 : NAN2M1D1 port map( A1 => data_in(0), A2 => 
                           coeff_memory_73_port, Z => mult_28_C92_n726);
   mult_28_C92_U586 : EXNOR2D1 port map( A1 => data_in(0), A2 => 
                           coeff_memory_73_port, Z => mult_28_C92_n725);
   mult_28_C92_U576 : EXNOR2D1 port map( A1 => data_in(10), A2 => 
                           coeff_memory_73_port, Z => mult_28_C92_n715);
   mult_28_C92_U575 : EXNOR2D1 port map( A1 => data_in(11), A2 => 
                           coeff_memory_73_port, Z => mult_28_C92_n714);
   mult_28_C92_U574 : EXNOR2D1 port map( A1 => data_in(12), A2 => 
                           coeff_memory_73_port, Z => mult_28_C92_n713);
   mult_28_C92_U573 : EXNOR2D1 port map( A1 => data_in(13), A2 => 
                           coeff_memory_73_port, Z => mult_28_C92_n712);
   mult_28_C92_U572 : EXNOR2D1 port map( A1 => data_in(14), A2 => 
                           coeff_memory_73_port, Z => mult_28_C92_n711);
   mult_28_C92_U571 : EXNOR2D1 port map( A1 => data_in(15), A2 => 
                           coeff_memory_73_port, Z => mult_28_C92_n710);
   mult_28_C92_U570 : NOR2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C92_n28, Z => mult_28_C92_n594);
   mult_28_C92_U569 : OAI22D1 port map( A1 => mult_28_C92_n725, A2 => 
                           mult_28_C92_n30, B1 => mult_28_C92_n724, B2 => 
                           mult_28_C92_n28, Z => mult_28_C92_n593);
   mult_28_C92_U566 : OAI22D1 port map( A1 => mult_28_C92_n722, A2 => 
                           mult_28_C92_n30, B1 => mult_28_C92_n721, B2 => 
                           mult_28_C92_n28, Z => mult_28_C92_n590);
   mult_28_C92_U565 : OAI22D1 port map( A1 => mult_28_C92_n1106, A2 => 
                           mult_28_C92_n30, B1 => mult_28_C92_n720, B2 => 
                           mult_28_C92_n28, Z => mult_28_C92_n589);
   mult_28_C92_U562 : OAI22D1 port map( A1 => mult_28_C92_n718, A2 => 
                           mult_28_C92_n30, B1 => mult_28_C92_n717, B2 => 
                           mult_28_C92_n28, Z => mult_28_C92_n586);
   mult_28_C92_U559 : OAI22D1 port map( A1 => mult_28_C92_n715, A2 => 
                           mult_28_C92_n30, B1 => mult_28_C92_n714, B2 => 
                           mult_28_C92_n28, Z => mult_28_C92_n583);
   mult_28_C92_U558 : OAI22D1 port map( A1 => mult_28_C92_n714, A2 => 
                           mult_28_C92_n30, B1 => mult_28_C92_n713, B2 => 
                           mult_28_C92_n28, Z => mult_28_C92_n582);
   mult_28_C92_U557 : OAI22D1 port map( A1 => mult_28_C92_n713, A2 => 
                           mult_28_C92_n30, B1 => mult_28_C92_n712, B2 => 
                           mult_28_C92_n28, Z => mult_28_C92_n581);
   mult_28_C92_U556 : OAI22D1 port map( A1 => mult_28_C92_n712, A2 => 
                           mult_28_C92_n30, B1 => mult_28_C92_n711, B2 => 
                           mult_28_C92_n28, Z => mult_28_C92_n580);
   mult_28_C92_U555 : OAI22D1 port map( A1 => mult_28_C92_n711, A2 => 
                           mult_28_C92_n30, B1 => mult_28_C92_n710, B2 => 
                           mult_28_C92_n28, Z => mult_28_C92_n343);
   mult_28_C92_U553 : OAI22D1 port map( A1 => mult_28_C92_n30, A2 => 
                           mult_28_C92_n1056, B1 => mult_28_C92_n726, B2 => 
                           mult_28_C92_n28, Z => mult_28_C92_n526);
   mult_28_C92_U551 : EXNOR2D1 port map( A1 => data_in(0), A2 => 
                           coeff_memory_75_port, Z => mult_28_C92_n708);
   mult_28_C92_U546 : EXNOR2D1 port map( A1 => data_in(5), A2 => 
                           coeff_memory_75_port, Z => mult_28_C92_n703);
   mult_28_C92_U545 : EXNOR2D1 port map( A1 => data_in(6), A2 => 
                           coeff_memory_75_port, Z => mult_28_C92_n702);
   mult_28_C92_U543 : EXNOR2D1 port map( A1 => data_in(8), A2 => 
                           coeff_memory_75_port, Z => mult_28_C92_n700);
   mult_28_C92_U542 : EXNOR2D1 port map( A1 => data_in(9), A2 => 
                           coeff_memory_75_port, Z => mult_28_C92_n699);
   mult_28_C92_U540 : EXNOR2D1 port map( A1 => data_in(11), A2 => 
                           coeff_memory_75_port, Z => mult_28_C92_n697);
   mult_28_C92_U539 : EXNOR2D1 port map( A1 => data_in(12), A2 => 
                           coeff_memory_75_port, Z => mult_28_C92_n696);
   mult_28_C92_U538 : EXNOR2D1 port map( A1 => data_in(13), A2 => 
                           coeff_memory_75_port, Z => mult_28_C92_n695);
   mult_28_C92_U537 : EXNOR2D1 port map( A1 => data_in(14), A2 => 
                           coeff_memory_75_port, Z => mult_28_C92_n694);
   mult_28_C92_U536 : EXNOR2D1 port map( A1 => data_in(15), A2 => 
                           coeff_memory_75_port, Z => mult_28_C92_n693);
   mult_28_C92_U535 : NOR2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C92_n34, Z => mult_28_C92_n578);
   mult_28_C92_U529 : OAI22D1 port map( A1 => mult_28_C92_n703, A2 => 
                           mult_28_C92_n36, B1 => mult_28_C92_n702, B2 => 
                           mult_28_C92_n34, Z => mult_28_C92_n572);
   mult_28_C92_U526 : OAI22D1 port map( A1 => mult_28_C92_n700, A2 => 
                           mult_28_C92_n36, B1 => mult_28_C92_n699, B2 => 
                           mult_28_C92_n34, Z => mult_28_C92_n569);
   mult_28_C92_U525 : OAI22D1 port map( A1 => mult_28_C92_n699, A2 => 
                           mult_28_C92_n36, B1 => mult_28_C92_n698, B2 => 
                           mult_28_C92_n34, Z => mult_28_C92_n568);
   mult_28_C92_U523 : OAI22D1 port map( A1 => mult_28_C92_n697, A2 => 
                           mult_28_C92_n36, B1 => mult_28_C92_n696, B2 => 
                           mult_28_C92_n34, Z => mult_28_C92_n566);
   mult_28_C92_U522 : OAI22D1 port map( A1 => mult_28_C92_n696, A2 => 
                           mult_28_C92_n36, B1 => mult_28_C92_n695, B2 => 
                           mult_28_C92_n34, Z => mult_28_C92_n565);
   mult_28_C92_U521 : OAI22D1 port map( A1 => mult_28_C92_n695, A2 => 
                           mult_28_C92_n36, B1 => mult_28_C92_n694, B2 => 
                           mult_28_C92_n34, Z => mult_28_C92_n564);
   mult_28_C92_U520 : OAI22D1 port map( A1 => mult_28_C92_n694, A2 => 
                           mult_28_C92_n36, B1 => mult_28_C92_n693, B2 => 
                           mult_28_C92_n34, Z => mult_28_C92_n329);
   mult_28_C92_U514 : EXNOR2D1 port map( A1 => data_in(2), A2 => 
                           coeff_memory_77_port, Z => mult_28_C92_n689);
   mult_28_C92_U512 : EXNOR2D1 port map( A1 => data_in(4), A2 => 
                           coeff_memory_77_port, Z => mult_28_C92_n687);
   mult_28_C92_U510 : EXNOR2D1 port map( A1 => data_in(6), A2 => 
                           coeff_memory_77_port, Z => mult_28_C92_n685);
   mult_28_C92_U508 : EXNOR2D1 port map( A1 => data_in(8), A2 => 
                           coeff_memory_77_port, Z => mult_28_C92_n683);
   mult_28_C92_U507 : EXNOR2D1 port map( A1 => data_in(9), A2 => 
                           coeff_memory_77_port, Z => mult_28_C92_n682);
   mult_28_C92_U506 : EXNOR2D1 port map( A1 => data_in(10), A2 => 
                           coeff_memory_77_port, Z => mult_28_C92_n681);
   mult_28_C92_U505 : EXNOR2D1 port map( A1 => data_in(11), A2 => 
                           coeff_memory_77_port, Z => mult_28_C92_n680);
   mult_28_C92_U504 : EXNOR2D1 port map( A1 => data_in(12), A2 => 
                           coeff_memory_77_port, Z => mult_28_C92_n679);
   mult_28_C92_U503 : EXNOR2D1 port map( A1 => data_in(13), A2 => 
                           coeff_memory_77_port, Z => mult_28_C92_n678);
   mult_28_C92_U502 : EXNOR2D1 port map( A1 => data_in(14), A2 => 
                           coeff_memory_77_port, Z => mult_28_C92_n677);
   mult_28_C92_U501 : EXNOR2D1 port map( A1 => data_in(15), A2 => 
                           coeff_memory_77_port, Z => mult_28_C92_n676);
   mult_28_C92_U500 : NOR2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C92_n40, Z => mult_28_C92_n562);
   mult_28_C92_U499 : OAI22D1 port map( A1 => mult_28_C92_n691, A2 => 
                           mult_28_C92_n42, B1 => mult_28_C92_n690, B2 => 
                           mult_28_C92_n40, Z => mult_28_C92_n561);
   mult_28_C92_U497 : OAI22D1 port map( A1 => mult_28_C92_n689, A2 => 
                           mult_28_C92_n42, B1 => mult_28_C92_n688, B2 => 
                           mult_28_C92_n40, Z => mult_28_C92_n559);
   mult_28_C92_U496 : OAI22D1 port map( A1 => mult_28_C92_n688, A2 => 
                           mult_28_C92_n42, B1 => mult_28_C92_n687, B2 => 
                           mult_28_C92_n40, Z => mult_28_C92_n558);
   mult_28_C92_U494 : OAI22D1 port map( A1 => mult_28_C92_n686, A2 => 
                           mult_28_C92_n42, B1 => mult_28_C92_n685, B2 => 
                           mult_28_C92_n40, Z => mult_28_C92_n556);
   mult_28_C92_U493 : OAI22D1 port map( A1 => mult_28_C92_n685, A2 => 
                           mult_28_C92_n42, B1 => mult_28_C92_n684, B2 => 
                           mult_28_C92_n40, Z => mult_28_C92_n555);
   mult_28_C92_U492 : OAI22D1 port map( A1 => mult_28_C92_n684, A2 => 
                           mult_28_C92_n42, B1 => mult_28_C92_n683, B2 => 
                           mult_28_C92_n40, Z => mult_28_C92_n554);
   mult_28_C92_U491 : OAI22D1 port map( A1 => mult_28_C92_n683, A2 => 
                           mult_28_C92_n42, B1 => mult_28_C92_n682, B2 => 
                           mult_28_C92_n40, Z => mult_28_C92_n553);
   mult_28_C92_U490 : OAI22D1 port map( A1 => mult_28_C92_n682, A2 => 
                           mult_28_C92_n42, B1 => mult_28_C92_n681, B2 => 
                           mult_28_C92_n40, Z => mult_28_C92_n552);
   mult_28_C92_U489 : OAI22D1 port map( A1 => mult_28_C92_n681, A2 => 
                           mult_28_C92_n42, B1 => mult_28_C92_n680, B2 => 
                           mult_28_C92_n40, Z => mult_28_C92_n551);
   mult_28_C92_U488 : OAI22D1 port map( A1 => mult_28_C92_n680, A2 => 
                           mult_28_C92_n42, B1 => mult_28_C92_n679, B2 => 
                           mult_28_C92_n40, Z => mult_28_C92_n550);
   mult_28_C92_U487 : OAI22D1 port map( A1 => mult_28_C92_n679, A2 => 
                           mult_28_C92_n42, B1 => mult_28_C92_n678, B2 => 
                           mult_28_C92_n40, Z => mult_28_C92_n549);
   mult_28_C92_U486 : OAI22D1 port map( A1 => mult_28_C92_n678, A2 => 
                           mult_28_C92_n42, B1 => mult_28_C92_n677, B2 => 
                           mult_28_C92_n40, Z => mult_28_C92_n548);
   mult_28_C92_U485 : OAI22D1 port map( A1 => mult_28_C92_n677, A2 => 
                           mult_28_C92_n42, B1 => mult_28_C92_n676, B2 => 
                           mult_28_C92_n40, Z => mult_28_C92_n319);
   mult_28_C92_U482 : NAN2M1D1 port map( A1 => data_in(0), A2 => 
                           coeff_memory_79_port, Z => mult_28_C92_n675);
   mult_28_C92_U478 : EXNOR2D1 port map( A1 => data_in(3), A2 => 
                           coeff_memory_79_port, Z => mult_28_C92_n671);
   mult_28_C92_U477 : EXNOR2D1 port map( A1 => data_in(4), A2 => 
                           coeff_memory_79_port, Z => mult_28_C92_n670);
   mult_28_C92_U475 : EXNOR2D1 port map( A1 => data_in(6), A2 => 
                           coeff_memory_79_port, Z => mult_28_C92_n668);
   mult_28_C92_U473 : EXNOR2D1 port map( A1 => data_in(8), A2 => 
                           coeff_memory_79_port, Z => mult_28_C92_n666);
   mult_28_C92_U470 : EXNOR2D1 port map( A1 => data_in(11), A2 => 
                           coeff_memory_79_port, Z => mult_28_C92_n663);
   mult_28_C92_U469 : EXNOR2D1 port map( A1 => data_in(12), A2 => 
                           coeff_memory_79_port, Z => mult_28_C92_n662);
   mult_28_C92_U468 : EXNOR2D1 port map( A1 => data_in(13), A2 => 
                           coeff_memory_79_port, Z => mult_28_C92_n661);
   mult_28_C92_U467 : EXNOR2D1 port map( A1 => data_in(14), A2 => 
                           coeff_memory_79_port, Z => mult_28_C92_n660);
   mult_28_C92_U465 : NOR2M1D1 port map( A1 => data_in(0), A2 => 
                           mult_28_C92_n46, Z => mult_28_C92_n546);
   mult_28_C92_U463 : OAI22D1 port map( A1 => mult_28_C92_n673, A2 => 
                           mult_28_C92_n48, B1 => mult_28_C92_n1057, B2 => 
                           mult_28_C92_n46, Z => mult_28_C92_n544);
   mult_28_C92_U460 : OAI22D1 port map( A1 => mult_28_C92_n670, A2 => 
                           mult_28_C92_n48, B1 => mult_28_C92_n669, B2 => 
                           mult_28_C92_n46, Z => mult_28_C92_n541);
   mult_28_C92_U459 : OAI22D1 port map( A1 => mult_28_C92_n669, A2 => 
                           mult_28_C92_n48, B1 => mult_28_C92_n668, B2 => 
                           mult_28_C92_n46, Z => mult_28_C92_n540);
   mult_28_C92_U458 : OAI22D1 port map( A1 => mult_28_C92_n668, A2 => 
                           mult_28_C92_n48, B1 => mult_28_C92_n667, B2 => 
                           mult_28_C92_n46, Z => mult_28_C92_n539);
   mult_28_C92_U457 : OAI22D1 port map( A1 => mult_28_C92_n667, A2 => 
                           mult_28_C92_n48, B1 => mult_28_C92_n666, B2 => 
                           mult_28_C92_n46, Z => mult_28_C92_n538);
   mult_28_C92_U456 : OAI22D1 port map( A1 => mult_28_C92_n666, A2 => 
                           mult_28_C92_n48, B1 => mult_28_C92_n665, B2 => 
                           mult_28_C92_n46, Z => mult_28_C92_n537);
   mult_28_C92_U454 : OAI22D1 port map( A1 => mult_28_C92_n664, A2 => 
                           mult_28_C92_n48, B1 => mult_28_C92_n663, B2 => 
                           mult_28_C92_n46, Z => mult_28_C92_n535);
   mult_28_C92_U453 : OAI22D1 port map( A1 => mult_28_C92_n663, A2 => 
                           mult_28_C92_n48, B1 => mult_28_C92_n662, B2 => 
                           mult_28_C92_n46, Z => mult_28_C92_n534);
   mult_28_C92_U452 : OAI22D1 port map( A1 => mult_28_C92_n662, A2 => 
                           mult_28_C92_n48, B1 => mult_28_C92_n661, B2 => 
                           mult_28_C92_n46, Z => mult_28_C92_n533);
   mult_28_C92_U449 : OAI22D1 port map( A1 => mult_28_C92_n48, A2 => 
                           mult_28_C92_n835, B1 => mult_28_C92_n675, B2 => 
                           mult_28_C92_n46, Z => mult_28_C92_n523);
   mult_28_C92_U448 : ADHALFD1 port map( A => mult_28_C92_n656, B => 
                           mult_28_C92_n529, CO => mult_28_C92_n521, S => 
                           mult_28_C92_n522);
   mult_28_C92_U447 : ADFULD1 port map( A => mult_28_C92_n655, B => 
                           mult_28_C92_n626, CI => mult_28_C92_n640, CO => 
                           mult_28_C92_n519, S => mult_28_C92_n520);
   mult_28_C92_U446 : ADHALFD1 port map( A => mult_28_C92_n654, B => 
                           mult_28_C92_n528, CO => mult_28_C92_n517, S => 
                           mult_28_C92_n518);
   mult_28_C92_U445 : ADFULD1 port map( A => mult_28_C92_n625, B => 
                           mult_28_C92_n639, CI => mult_28_C92_n518, CO => 
                           mult_28_C92_n515, S => mult_28_C92_n516);
   mult_28_C92_U444 : ADFULD1 port map( A => mult_28_C92_n653, B => 
                           mult_28_C92_n610, CI => mult_28_C92_n638, CO => 
                           mult_28_C92_n513, S => mult_28_C92_n514);
   mult_28_C92_U443 : ADFULD1 port map( A => mult_28_C92_n517, B => 
                           mult_28_C92_n624, CI => mult_28_C92_n514, CO => 
                           mult_28_C92_n511, S => mult_28_C92_n512);
   mult_28_C92_U441 : ADFULD1 port map( A => mult_28_C92_n609, B => 
                           mult_28_C92_n652, CI => mult_28_C92_n637, CO => 
                           mult_28_C92_n507, S => mult_28_C92_n508);
   mult_28_C92_U440 : ADFULD1 port map( A => mult_28_C92_n513, B => 
                           mult_28_C92_n510, CI => mult_28_C92_n508, CO => 
                           mult_28_C92_n505, S => mult_28_C92_n506);
   mult_28_C92_U439 : ADFULD1 port map( A => mult_28_C92_n622, B => 
                           mult_28_C92_n594, CI => mult_28_C92_n651, CO => 
                           mult_28_C92_n503, S => mult_28_C92_n504);
   mult_28_C92_U438 : ADFULD1 port map( A => mult_28_C92_n608, B => 
                           mult_28_C92_n636, CI => mult_28_C92_n509, CO => 
                           mult_28_C92_n501, S => mult_28_C92_n502);
   mult_28_C92_U437 : ADFULD1 port map( A => mult_28_C92_n504, B => 
                           mult_28_C92_n507, CI => mult_28_C92_n502, CO => 
                           mult_28_C92_n499, S => mult_28_C92_n500);
   mult_28_C92_U436 : ADHALFD1 port map( A => mult_28_C92_n607, B => 
                           mult_28_C92_n526, CO => mult_28_C92_n497, S => 
                           mult_28_C92_n498);
   mult_28_C92_U434 : ADFULD1 port map( A => mult_28_C92_n498, B => 
                           mult_28_C92_n650, CI => mult_28_C92_n503, CO => 
                           mult_28_C92_n493, S => mult_28_C92_n494);
   mult_28_C92_U433 : ADFULD1 port map( A => mult_28_C92_n496, B => 
                           mult_28_C92_n501, CI => mult_28_C92_n494, CO => 
                           mult_28_C92_n491, S => mult_28_C92_n492);
   mult_28_C92_U432 : ADFULD1 port map( A => mult_28_C92_n606, B => 
                           mult_28_C92_n578, CI => mult_28_C92_n649, CO => 
                           mult_28_C92_n489, S => mult_28_C92_n490);
   mult_28_C92_U430 : ADFULD1 port map( A => mult_28_C92_n495, B => 
                           mult_28_C92_n497, CI => mult_28_C92_n490, CO => 
                           mult_28_C92_n485, S => mult_28_C92_n486);
   mult_28_C92_U416 : ADFULD1 port map( A => mult_28_C92_n561, B => 
                           mult_28_C92_n617, CI => mult_28_C92_n589, CO => 
                           mult_28_C92_n457, S => mult_28_C92_n458);
   mult_28_C92_U414 : ADFULD1 port map( A => mult_28_C92_n458, B => 
                           mult_28_C92_n460, CI => mult_28_C92_n467, CO => 
                           mult_28_C92_n453, S => mult_28_C92_n454);
   mult_28_C92_U411 : ADFULD1 port map( A => mult_28_C92_n560, B => 
                           mult_28_C92_n630, CI => mult_28_C92_n588, CO => 
                           mult_28_C92_n447, S => mult_28_C92_n448);
   mult_28_C92_U406 : ADHALFD1 port map( A => mult_28_C92_n559, B => 
                           mult_28_C92_n523, CO => mult_28_C92_n437, S => 
                           mult_28_C92_n438);
   mult_28_C92_U405 : ADFULD1 port map( A => mult_28_C92_n545, B => 
                           mult_28_C92_n601, CI => mult_28_C92_n573, CO => 
                           mult_28_C92_n435, S => mult_28_C92_n436);
   mult_28_C92_U404 : ADFULD1 port map( A => mult_28_C92_n644, B => 
                           mult_28_C92_n587, CI => mult_28_C92_n615, CO => 
                           mult_28_C92_n433, S => mult_28_C92_n434);
   mult_28_C92_U403 : ADFULD1 port map( A => mult_28_C92_n438, B => 
                           mult_28_C92_n629, CI => mult_28_C92_n449, CO => 
                           mult_28_C92_n431, S => mult_28_C92_n432);
   mult_28_C92_U401 : ADFULD1 port map( A => mult_28_C92_n432, B => 
                           mult_28_C92_n436, CI => mult_28_C92_n443, CO => 
                           mult_28_C92_n427, S => mult_28_C92_n428);
   mult_28_C92_U399 : OR2D1 port map( A1 => mult_28_C92_n600, A2 => 
                           mult_28_C92_n558, Z => mult_28_C92_n423);
   mult_28_C92_U396 : ADFULD1 port map( A => mult_28_C92_n614, B => 
                           mult_28_C92_n628, CI => mult_28_C92_n572, CO => 
                           mult_28_C92_n419, S => mult_28_C92_n420);
   mult_28_C92_U390 : ADFULD1 port map( A => mult_28_C92_n613, B => 
                           mult_28_C92_n571, CI => mult_28_C92_n543, CO => 
                           mult_28_C92_n407, S => mult_28_C92_n408);
   mult_28_C92_U388 : ADFULD1 port map( A => mult_28_C92_n423, B => 
                           mult_28_C92_n410, CI => mult_28_C92_n421, CO => 
                           mult_28_C92_n403, S => mult_28_C92_n404);
   mult_28_C92_U386 : ADFULD1 port map( A => mult_28_C92_n404, B => 
                           mult_28_C92_n417, CI => mult_28_C92_n415, CO => 
                           mult_28_C92_n399, S => mult_28_C92_n400);
   mult_28_C92_U385 : ADFULD1 port map( A => mult_28_C92_n413, B => 
                           mult_28_C92_n402, CI => mult_28_C92_n400, CO => 
                           mult_28_C92_n397, S => mult_28_C92_n398);
   mult_28_C92_U384 : ADFULD1 port map( A => mult_28_C92_n409, B => 
                           mult_28_C92_n542, CI => mult_28_C92_n627, CO => 
                           mult_28_C92_n395, S => mult_28_C92_n396);
   mult_28_C92_U383 : ADFULD1 port map( A => mult_28_C92_n612, B => 
                           mult_28_C92_n556, CI => mult_28_C92_n598, CO => 
                           mult_28_C92_n393, S => mult_28_C92_n394);
   mult_28_C92_U380 : ADFULD1 port map( A => mult_28_C92_n392, B => 
                           mult_28_C92_n403, CI => mult_28_C92_n401, CO => 
                           mult_28_C92_n387, S => mult_28_C92_n388);
   mult_28_C92_U377 : ADFULD1 port map( A => mult_28_C92_n597, B => 
                           mult_28_C92_n569, CI => mult_28_C92_n583, CO => 
                           mult_28_C92_n381, S => mult_28_C92_n382);
   mult_28_C92_U376 : ADFULD1 port map( A => mult_28_C92_n541, B => 
                           mult_28_C92_n555, CI => mult_28_C92_n384, CO => 
                           mult_28_C92_n379, S => mult_28_C92_n380);
   mult_28_C92_U375 : ADFULD1 port map( A => mult_28_C92_n393, B => 
                           mult_28_C92_n395, CI => mult_28_C92_n382, CO => 
                           mult_28_C92_n377, S => mult_28_C92_n378);
   mult_28_C92_U371 : ADFULD1 port map( A => mult_28_C92_n554, B => 
                           mult_28_C92_n596, CI => mult_28_C92_n568, CO => 
                           mult_28_C92_n369, S => mult_28_C92_n370);
   mult_28_C92_U370 : ADFULD1 port map( A => mult_28_C92_n381, B => 
                           mult_28_C92_n582, CI => mult_28_C92_n379, CO => 
                           mult_28_C92_n367, S => mult_28_C92_n368);
   mult_28_C92_U369 : ADFULD1 port map( A => mult_28_C92_n372, B => 
                           mult_28_C92_n370, CI => mult_28_C92_n377, CO => 
                           mult_28_C92_n365, S => mult_28_C92_n366);
   mult_28_C92_U368 : ADFULD1 port map( A => mult_28_C92_n375, B => 
                           mult_28_C92_n368, CI => mult_28_C92_n366, CO => 
                           mult_28_C92_n363, S => mult_28_C92_n364);
   mult_28_C92_U366 : ADFULD1 port map( A => mult_28_C92_n581, B => 
                           mult_28_C92_n553, CI => mult_28_C92_n539, CO => 
                           mult_28_C92_n359, S => mult_28_C92_n360);
   mult_28_C92_U365 : ADFULD1 port map( A => mult_28_C92_n362, B => 
                           mult_28_C92_n567, CI => mult_28_C92_n371, CO => 
                           mult_28_C92_n357, S => mult_28_C92_n358);
   mult_28_C92_U364 : ADFULD1 port map( A => mult_28_C92_n360, B => 
                           mult_28_C92_n369, CI => mult_28_C92_n367, CO => 
                           mult_28_C92_n355, S => mult_28_C92_n356);
   mult_28_C92_U363 : ADFULD1 port map( A => mult_28_C92_n365, B => 
                           mult_28_C92_n358, CI => mult_28_C92_n356, CO => 
                           mult_28_C92_n353, S => mult_28_C92_n354);
   mult_28_C92_U362 : ADFULD1 port map( A => mult_28_C92_n580, B => 
                           mult_28_C92_n538, CI => mult_28_C92_n595, CO => 
                           mult_28_C92_n351, S => mult_28_C92_n352);
   mult_28_C92_U361 : ADFULD1 port map( A => mult_28_C92_n552, B => 
                           mult_28_C92_n361, CI => mult_28_C92_n566, CO => 
                           mult_28_C92_n349, S => mult_28_C92_n350);
   mult_28_C92_U360 : ADFULD1 port map( A => mult_28_C92_n350, B => 
                           mult_28_C92_n359, CI => mult_28_C92_n352, CO => 
                           mult_28_C92_n347, S => mult_28_C92_n348);
   mult_28_C92_U359 : ADFULD1 port map( A => mult_28_C92_n348, B => 
                           mult_28_C92_n357, CI => mult_28_C92_n355, CO => 
                           mult_28_C92_n345, S => mult_28_C92_n346);
   mult_28_C92_U357 : ADFULD1 port map( A => mult_28_C92_n537, B => 
                           mult_28_C92_n551, CI => mult_28_C92_n565, CO => 
                           mult_28_C92_n341, S => mult_28_C92_n342);
   mult_28_C92_U356 : ADFULD1 port map( A => mult_28_C92_n351, B => 
                           mult_28_C92_n344, CI => mult_28_C92_n349, CO => 
                           mult_28_C92_n339, S => mult_28_C92_n340);
   mult_28_C92_U355 : ADFULD1 port map( A => mult_28_C92_n347, B => 
                           mult_28_C92_n342, CI => mult_28_C92_n340, CO => 
                           mult_28_C92_n337, S => mult_28_C92_n338);
   mult_28_C92_U354 : ADFULD1 port map( A => mult_28_C92_n550, B => 
                           mult_28_C92_n536, CI => mult_28_C92_n579, CO => 
                           mult_28_C92_n335, S => mult_28_C92_n336);
   mult_28_C92_U353 : ADFULD1 port map( A => mult_28_C92_n343, B => 
                           mult_28_C92_n564, CI => mult_28_C92_n341, CO => 
                           mult_28_C92_n333, S => mult_28_C92_n334);
   mult_28_C92_U352 : ADFULD1 port map( A => mult_28_C92_n339, B => 
                           mult_28_C92_n336, CI => mult_28_C92_n334, CO => 
                           mult_28_C92_n331, S => mult_28_C92_n332);
   mult_28_C92_U350 : ADFULD1 port map( A => mult_28_C92_n535, B => 
                           mult_28_C92_n549, CI => mult_28_C92_n330, CO => 
                           mult_28_C92_n327, S => mult_28_C92_n328);
   mult_28_C92_U349 : ADFULD1 port map( A => mult_28_C92_n328, B => 
                           mult_28_C92_n335, CI => mult_28_C92_n333, CO => 
                           mult_28_C92_n325, S => mult_28_C92_n326);
   mult_28_C92_U348 : ADFULD1 port map( A => mult_28_C92_n548, B => 
                           mult_28_C92_n329, CI => mult_28_C92_n563, CO => 
                           mult_28_C92_n323, S => mult_28_C92_n324);
   mult_28_C92_U347 : ADFULD1 port map( A => mult_28_C92_n327, B => 
                           mult_28_C92_n534, CI => mult_28_C92_n324, CO => 
                           mult_28_C92_n321, S => mult_28_C92_n322);
   mult_28_C92_U345 : ADFULD1 port map( A => mult_28_C92_n320, B => 
                           mult_28_C92_n533, CI => mult_28_C92_n323, CO => 
                           mult_28_C92_n317, S => mult_28_C92_n318);
   mult_28_C92_U344 : ADFULD1 port map( A => mult_28_C92_n532, B => 
                           mult_28_C92_n319, CI => mult_28_C92_n547, CO => 
                           mult_28_C92_n315, S => mult_28_C92_n316);
   mult_28_C92_U330 : AOI21D1 port map( A1 => mult_28_C92_n1150, A2 => 
                           mult_28_C92_n1152, B => mult_28_C92_n1151, Z => 
                           mult_28_C92_n277);
   mult_28_C92_U324 : OAI21D1 port map( A1 => mult_28_C92_n275, A2 => 
                           mult_28_C92_n277, B => mult_28_C92_n276, Z => 
                           mult_28_C92_n274);
   mult_28_C92_U242 : NOR2D2 port map( A1 => mult_28_C92_net11792, A2 => 
                           mult_28_C92_n463, Z => mult_28_C92_n220);
   mult_28_C92_U215 : NOR2D2 port map( A1 => mult_28_C92_n412, A2 => 
                           mult_28_C92_n425, Z => mult_28_C92_n202);
   mult_28_C92_U163 : NOR2D2 port map( A1 => mult_28_C92_n354, A2 => 
                           mult_28_C92_n363, Z => mult_28_C92_n161);
   mult_28_C92_U156 : OAI21D1 port map( A1 => mult_28_C92_n171, A2 => 
                           mult_28_C92_n161, B => mult_28_C92_n162, Z => 
                           mult_28_C92_n160);
   mult_28_C92_U154 : AOI21D1 port map( A1 => mult_28_C92_n159, A2 => 
                           mult_28_C92_net12273, B => mult_28_C92_n160, Z => 
                           mult_28_C92_n158);
   mult_28_C92_U142 : OAI21D1 port map( A1 => mult_28_C92_n171, A2 => 
                           mult_28_C92_n150, B => mult_28_C92_n151, Z => 
                           mult_28_C92_n149);
   mult_28_C92_U140 : AOI21D1 port map( A1 => mult_28_C92_net12273, A2 => 
                           mult_28_C92_n148, B => mult_28_C92_n149, Z => 
                           mult_28_C92_n147);
   mult_28_C92_U111 : NOR2D2 port map( A1 => mult_28_C92_n326, A2 => 
                           mult_28_C92_n331, Z => mult_28_C92_n125);
   mult_28_C92_U108 : OAI21D1 port map( A1 => mult_28_C92_n133, A2 => 
                           mult_28_C92_n125, B => mult_28_C92_n126, Z => 
                           mult_28_C92_n120);
   mult_28_C92_U80 : OAI21D1 port map( A1 => mult_28_C92_n113, A2 => 
                           mult_28_C92_n103, B => mult_28_C92_n104, Z => 
                           mult_28_C92_n102);
   mult_28_C92_U78 : AOI21D1 port map( A1 => mult_28_C92_n120, A2 => 
                           mult_28_C92_n101, B => mult_28_C92_n102, Z => 
                           mult_28_C92_n100);
   mult_28_C92_U59 : EXOR2D1 port map( A1 => mult_28_C92_n94, A2 => 
                           mult_28_C92_n55, Z => m1_14);
   mult_28_C92_U54 : EXOR2D1 port map( A1 => mult_28_C92_n85, A2 => 
                           mult_28_C92_n54, Z => m1_15);
   add_102_U267 : INVBD2 port map( A => add_102_n105, Z => add_102_n129);
   add_102_U266 : AOI21DL port map( A1 => add_102_n1, A2 => add_102_n44, B => 
                           add_102_n193, Z => add_102_n43);
   add_102_U265 : EXOR2D4 port map( A1 => add_102_n52, A2 => add_102_n6, Z => 
                           y_11_port);
   add_102_U264 : EXOR2D4 port map( A1 => add_102_n27, A2 => add_102_n3, Z => 
                           y_14_port);
   add_102_U263 : EXOR2D4 port map( A1 => add_102_n43, A2 => add_102_n5, Z => 
                           y_12_port);
   add_102_U262 : EXOR2D4 port map( A1 => add_102_n71, A2 => add_102_n9, Z => 
                           y_8_port);
   add_102_U261 : AOI21DL port map( A1 => add_102_n1, A2 => add_102_n21, B => 
                           add_102_n22, Z => add_102_n20);
   add_102_U260 : EXOR2D4 port map( A1 => add_102_n20, A2 => add_102_n2, Z => 
                           y_15_port);
   add_102_U259 : EXOR2D4 port map( A1 => add_102_n36, A2 => add_102_n4, Z => 
                           y_13_port);
   add_102_U258 : EXOR2D4 port map( A1 => add_102_n80, A2 => add_102_n10, Z => 
                           y_7_port);
   add_102_U257 : NOR2D1 port map( A1 => add_102_n55, A2 => add_102_n50, Z => 
                           add_102_n44);
   add_102_U256 : EXOR2D4 port map( A1 => add_102_n102, A2 => add_102_n14, Z =>
                           y_3_port);
   add_102_U255 : NAN2D1 port map( A1 => add_102_n129, A2 => add_102_n106, Z =>
                           add_102_n15);
   add_102_U254 : NAN2DL port map( A1 => add_102_n101, A2 => add_102_n98, Z => 
                           add_102_n14);
   add_102_U253 : NAN2D1 port map( A1 => z2_3_port, A2 => m1_3, Z => 
                           add_102_n101);
   add_102_U252 : EXOR2D4 port map( A1 => add_102_n94, A2 => add_102_n13, Z => 
                           y_4_port);
   add_102_U251 : EXNOR2D2 port map( A1 => add_102_n16, A2 => add_102_n113, Z 
                           => y_1_port);
   add_102_U250 : NAN2D1 port map( A1 => add_102_n188, A2 => add_102_net11859, 
                           Z => add_102_n10);
   add_102_U249 : NAN2DL port map( A1 => add_102_n202, A2 => add_102_n112, Z =>
                           add_102_n16);
   add_102_U248 : NAN2DL port map( A1 => add_102_n53, A2 => add_102_n56, Z => 
                           add_102_n7);
   add_102_U247 : NOR2D1 port map( A1 => add_102_n39, A2 => add_102_n34, Z => 
                           add_102_n32);
   add_102_U246 : OA21M20DL port map( A1 => add_102_n1, A2 => add_102_n28, B =>
                           add_102_n31, Z => add_102_n27);
   add_102_U245 : EXNOR2D1 port map( A1 => add_102_n1, A2 => add_102_n7, Z => 
                           y_10_port);
   add_102_U244 : INVD1 port map( A => add_102_n95, Z => add_102_n94);
   add_102_U243 : AOI21DL port map( A1 => add_102_n1, A2 => add_102_n37, B => 
                           add_102_n38, Z => add_102_n36);
   add_102_U242 : NAN2D1 port map( A1 => m1_5, A2 => z2_5_port, Z => 
                           add_102_n90);
   add_102_U241 : OR2D1 port map( A1 => m1_15, A2 => z2_15_port, Z => 
                           add_102_n201);
   add_102_U240 : NAN2D1 port map( A1 => m1_12, A2 => z2_12_port, Z => 
                           add_102_n42);
   add_102_U239 : NAN2D1 port map( A1 => z2_0_port, A2 => m1_0, Z => 
                           add_102_n115);
   add_102_U238 : NAN2D1 port map( A1 => m1_11, A2 => z2_11_port, Z => 
                           add_102_n51);
   add_102_U237 : NAN2DL port map( A1 => m1_15, A2 => z2_15_port, Z => 
                           add_102_n19);
   add_102_U236 : NAN2D1 port map( A1 => add_102_n201, A2 => add_102_n19, Z => 
                           add_102_n2);
   add_102_U235 : INVDL port map( A => add_102_n45, Z => add_102_n47);
   add_102_U234 : NOR2M1DL port map( A1 => add_102_n44, A2 => add_102_n39, Z =>
                           add_102_n37);
   add_102_U233 : INVDL port map( A => add_102_n34, Z => add_102_n118);
   add_102_U232 : INVDL port map( A => add_102_n39, Z => add_102_n119);
   add_102_U231 : OA21M20D1 port map( A1 => add_102_n98, A2 => add_102_n104, B 
                           => add_102_n101, Z => add_102_n97);
   add_102_U230 : OA21M20D1 port map( A1 => add_102_n187, A2 => add_102_n113, B
                           => add_102_n112, Z => add_102_n108);
   add_102_U229 : INVDL port map( A => add_102_n23, Z => add_102_n117);
   add_102_U228 : INVDL port map( A => add_102_n50, Z => add_102_n120);
   add_102_U227 : NAN2D1 port map( A1 => add_102_n32, A2 => add_102_n44, Z => 
                           add_102_n30);
   add_102_U226 : NAN2D1 port map( A1 => m1_14, A2 => z2_14_port, Z => 
                           add_102_n26);
   add_102_U225 : NAN2D1 port map( A1 => m1_13, A2 => z2_13_port, Z => 
                           add_102_n35);
   add_102_U224 : NOR2DL port map( A1 => add_102_n30, A2 => add_102_n23, Z => 
                           add_102_n21);
   add_102_U223 : NAN2M1DL port map( A1 => add_102_n92, A2 => add_102_n93, Z =>
                           add_102_n13);
   add_102_U222 : INVDL port map( A => add_102_n55, Z => add_102_n53);
   add_102_U221 : NAN2M1DL port map( A1 => add_102_n89, A2 => add_102_n90, Z =>
                           add_102_n12);
   add_102_U220 : INVDL port map( A => add_102_n30, Z => add_102_n28);
   add_102_U219 : OR2DL port map( A1 => m1_0, A2 => z2_0_port, Z => 
                           add_102_n200);
   add_102_U218 : NAN2DL port map( A1 => add_102_n200, A2 => add_102_n115, Z =>
                           add_102_n17);
   add_102_U217 : NAN2D2 port map( A1 => add_102_net11441, A2 => add_102_n59, Z
                           => add_102_n1);
   add_102_U216 : INVDL port map( A => add_102_n17, Z => y_0_port);
   add_102_U215 : NAN2D1 port map( A1 => add_102_n129, A2 => add_102_n98, Z => 
                           add_102_n96);
   add_102_U214 : NAN2D1 port map( A1 => add_102_n81, A2 => add_102_net11615, Z
                           => add_102_net11329);
   add_102_U213 : INVDL port map( A => add_102_n108, Z => add_102_n199);
   add_102_U212 : INVD1 port map( A => add_102_n199, Z => add_102_n196);
   add_102_U211 : INVD2 port map( A => add_102_n15, Z => add_102_n195);
   add_102_U210 : NAN2D2 port map( A1 => add_102_n198, A2 => add_102_n197, Z =>
                           y_2_port);
   add_102_U209 : NAN2D2 port map( A1 => add_102_n196, A2 => add_102_n195, Z =>
                           add_102_n198);
   add_102_U208 : NAN2D1 port map( A1 => add_102_n199, A2 => add_102_n15, Z => 
                           add_102_n197);
   add_102_U207 : AOI21D1 port map( A1 => add_102_n107, A2 => add_102_n190, B 
                           => add_102_n104, Z => add_102_n102);
   add_102_U206 : NAN2D1 port map( A1 => add_102_n117, A2 => add_102_n26, Z => 
                           add_102_n3);
   add_102_U205 : NAN2M1DL port map( A1 => add_102_n194, A2 => m1_1, Z => 
                           add_102_n112);
   add_102_U204 : INVDL port map( A => add_102_net11615, Z => add_102_n82);
   add_102_U203 : INVD2 port map( A => add_102_n106, Z => add_102_n104);
   add_102_U202 : OAI21DL port map( A1 => add_102_n34, A2 => add_102_n42, B => 
                           add_102_n35, Z => add_102_n33);
   add_102_U201 : OAI21DL port map( A1 => add_102_n47, A2 => add_102_n39, B => 
                           add_102_n42, Z => add_102_n38);
   add_102_U200 : NAN2DL port map( A1 => add_102_n119, A2 => add_102_n42, Z => 
                           add_102_n5);
   add_102_U199 : INVDL port map( A => add_102_n47, Z => add_102_n193);
   add_102_U198 : INVDL port map( A => add_102_net12241, Z => add_102_net12242)
                           ;
   add_102_U197 : NAN2DL port map( A1 => z2_7_port, A2 => add_102_net12242, Z 
                           => add_102_net11859);
   add_102_U196 : INVDL port map( A => m1_7, Z => add_102_net12241);
   add_102_U195 : NOR2D1 port map( A1 => add_102_n89, A2 => add_102_n92, Z => 
                           add_102_n87);
   add_102_U194 : EXOR2D4 port map( A1 => add_102_n86, A2 => add_102_net11329, 
                           Z => y_6_port);
   add_102_U193 : NAN2M1DL port map( A1 => add_102_n192, A2 => m1_7, Z => 
                           add_102_n79);
   add_102_U192 : OAI21DL port map( A1 => add_102_n70, A2 => add_102_n62, B => 
                           add_102_n63, Z => add_102_n61);
   add_102_U191 : NAN2D1 port map( A1 => m1_9, A2 => z2_9_port, Z => 
                           add_102_n63);
   add_102_U190 : NAN2D2 port map( A1 => add_102_net11439, A2 => 
                           add_102_net11440, Z => add_102_net11441);
   add_102_U189 : AOI21DL port map( A1 => add_102_net11440, A2 => add_102_n81, 
                           B => add_102_n82, Z => add_102_n80);
   add_102_U188 : INVD2 port map( A => add_102_n86, Z => add_102_net11440);
   add_102_U187 : INVDL port map( A => add_102_n75, Z => add_102_net11486);
   add_102_U186 : INVDL port map( A => add_102_n73, Z => add_102_n75);
   add_102_U185 : INVDL port map( A => add_102_n62, Z => add_102_n122);
   add_102_U184 : EXOR2D4 port map( A1 => add_102_n64, A2 => add_102_n8, Z => 
                           y_9_port);
   add_102_U183 : NAN2D1 port map( A1 => m1_6, A2 => z2_6_port, Z => 
                           add_102_n84);
   add_102_U182 : NAN2DL port map( A1 => z2_6_port, A2 => m1_6, Z => 
                           add_102_net11615);
   add_102_U181 : NOR2D2 port map( A1 => m1_6, A2 => z2_6_port, Z => 
                           add_102_n83);
   add_102_U180 : NAN2D1 port map( A1 => z2_8_port, A2 => m1_8, Z => 
                           add_102_n70);
   add_102_U179 : INVDL port map( A => add_102_n83, Z => add_102_n81);
   add_102_U178 : BUFDL port map( A => add_102_n67, Z => add_102_net12276);
   add_102_U177 : AOI21DL port map( A1 => add_102_net11440, A2 => add_102_n72, 
                           B => add_102_net11486, Z => add_102_n71);
   add_102_U176 : NAN2D2 port map( A1 => add_102_n72, A2 => add_102_n60, Z => 
                           add_102_n58);
   add_102_U175 : NOR2D1 port map( A1 => add_102_n78, A2 => add_102_n83, Z => 
                           add_102_n72);
   add_102_U174 : NAN2DL port map( A1 => add_102_n123, A2 => add_102_n70, Z => 
                           add_102_n9);
   add_102_U173 : INVDL port map( A => add_102_n67, Z => add_102_n123);
   add_102_U172 : AOI21DL port map( A1 => add_102_n65, A2 => add_102_net11440, 
                           B => add_102_n66, Z => add_102_n64);
   add_102_U171 : EXNOR2D2 port map( A1 => add_102_n91, A2 => add_102_n12, Z =>
                           y_5_port);
   add_102_U170 : INVDL port map( A => add_102_n56, Z => add_102_n191);
   add_102_U169 : AOI21M10D1 port map( A1 => add_102_n55, A2 => add_102_n1, B 
                           => add_102_n191, Z => add_102_n52);
   add_102_U168 : NOR2D2 port map( A1 => m1_10, A2 => z2_10_port, Z => 
                           add_102_n55);
   add_102_U167 : INVBD2 port map( A => add_102_n100, Z => add_102_n98);
   add_102_U166 : INVD1 port map( A => add_102_n189, Z => add_102_n190);
   add_102_U165 : INVDL port map( A => add_102_n129, Z => add_102_n189);
   add_102_U164 : INVD1 port map( A => add_102_n108, Z => add_102_n107);
   add_102_U163 : INVD1 port map( A => add_102_n115, Z => add_102_n113);
   add_102_U162 : INVD2 port map( A => add_102_n58, Z => add_102_net11439);
   add_102_U161 : OR2D1 port map( A1 => z2_7_port, A2 => add_102_net12242, Z =>
                           add_102_n188);
   add_102_U160 : INVD1 port map( A => z2_1_port, Z => add_102_n194);
   add_102_U159 : NAN2DL port map( A1 => add_102_n118, A2 => add_102_n35, Z => 
                           add_102_n4);
   add_102_U158 : NAN2DL port map( A1 => add_102_n120, A2 => add_102_n51, Z => 
                           add_102_n6);
   add_102_U157 : NAN2DL port map( A1 => add_102_n122, A2 => add_102_n63, Z => 
                           add_102_n8);
   add_102_U156 : INVD1 port map( A => z2_7_port, Z => add_102_n192);
   add_102_U155 : AND2D1 port map( A1 => add_102_n72, A2 => add_102_n123, Z => 
                           add_102_n65);
   add_102_U154 : NAN2M1DL port map( A1 => m1_1, A2 => add_102_n194, Z => 
                           add_102_n202);
   add_102_U153 : NAN2M1D1 port map( A1 => m1_1, A2 => add_102_n194, Z => 
                           add_102_n187);
   add_102_U152 : OAI21D1 port map( A1 => add_102_n75, A2 => add_102_net12276, 
                           B => add_102_n70, Z => add_102_n66);
   add_102_U151 : NOR2D1 port map( A1 => m1_13, A2 => z2_13_port, Z => 
                           add_102_n34);
   add_102_U77 : NOR2D2 port map( A1 => m1_8, A2 => z2_8_port, Z => add_102_n67
                           );
   add_102_U63 : NOR2D2 port map( A1 => add_102_n67, A2 => add_102_n62, Z => 
                           add_102_n60);
   add_102_U86 : OAI21D1 port map( A1 => add_102_n78, A2 => add_102_n84, B => 
                           add_102_n79, Z => add_102_n73);
   add_102_U67 : NOR2D2 port map( A1 => m1_9, A2 => z2_9_port, Z => add_102_n62
                           );
   add_102_U62 : AOI21D1 port map( A1 => add_102_n60, A2 => add_102_n73, B => 
                           add_102_n61, Z => add_102_n59);
   add_102_U101 : AOI21D1 port map( A1 => add_102_n95, A2 => add_102_n87, B => 
                           add_102_n88, Z => add_102_n86);
   add_102_U103 : OAI21D1 port map( A1 => add_102_n89, A2 => add_102_n93, B => 
                           add_102_n90, Z => add_102_n88);
   add_102_U89 : NOR2D2 port map( A1 => m1_7, A2 => z2_7_port, Z => add_102_n78
                           );
   add_102_U132 : NAN2D2 port map( A1 => m1_2, A2 => z2_2_port, Z => 
                           add_102_n106);
   add_102_U131 : NOR2D2 port map( A1 => m1_2, A2 => z2_2_port, Z => 
                           add_102_n105);
   add_102_U123 : NOR2D2 port map( A1 => m1_3, A2 => z2_3_port, Z => 
                           add_102_n100);
   add_102_U116 : OAI21D1 port map( A1 => add_102_n96, A2 => add_102_n108, B =>
                           add_102_n97, Z => add_102_n95);
   add_102_U113 : NAN2D2 port map( A1 => m1_4, A2 => z2_4_port, Z => 
                           add_102_n93);
   add_102_U112 : NOR2D2 port map( A1 => m1_4, A2 => z2_4_port, Z => 
                           add_102_n92);
   add_102_U109 : OAI21D1 port map( A1 => add_102_n94, A2 => add_102_n92, B => 
                           add_102_n93, Z => add_102_n91);
   add_102_U106 : NOR2D2 port map( A1 => m1_5, A2 => z2_5_port, Z => 
                           add_102_n89);
   add_102_U58 : NAN2D2 port map( A1 => m1_10, A2 => z2_10_port, Z => 
                           add_102_n56);
   add_102_U49 : NOR2D2 port map( A1 => m1_11, A2 => z2_11_port, Z => 
                           add_102_n50);
   add_102_U46 : OAI21D1 port map( A1 => add_102_n50, A2 => add_102_n56, B => 
                           add_102_n51, Z => add_102_n45);
   add_102_U37 : NOR2D2 port map( A1 => m1_12, A2 => z2_12_port, Z => 
                           add_102_n39);
   add_102_U22 : AOI21D1 port map( A1 => add_102_n32, A2 => add_102_n45, B => 
                           add_102_n33, Z => add_102_n31);
   add_102_U15 : NOR2D2 port map( A1 => m1_14, A2 => z2_14_port, Z => 
                           add_102_n23);
   add_102_U10 : OAI21D1 port map( A1 => add_102_n31, A2 => add_102_n23, B => 
                           add_102_n26, Z => add_102_n22);
   add_0_root_add_0_root_add_101_U248 : OAI21DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n75, A2 => 
                           add_0_root_add_0_root_add_101_net12355, B => 
                           add_0_root_add_0_root_add_101_n70, Z => 
                           add_0_root_add_0_root_add_101_n66);
   add_0_root_add_0_root_add_101_U247 : NAN2D1 port map( A1 => m3_7, A2 => 
                           z2_temp_7, Z => add_0_root_add_0_root_add_101_n79);
   add_0_root_add_0_root_add_101_U246 : NAN2DL port map( A1 => m3_5, A2 => 
                           z2_temp_5, Z => add_0_root_add_0_root_add_101_n90);
   add_0_root_add_0_root_add_101_U245 : NOR2D1 port map( A1 => z2_temp_10, A2 
                           => m3_10, Z => add_0_root_add_0_root_add_101_n55);
   add_0_root_add_0_root_add_101_U244 : NAN2DL port map( A1 => m3_13, A2 => 
                           z2_temp_13, Z => add_0_root_add_0_root_add_101_n35);
   add_0_root_add_0_root_add_101_U243 : NAN2D1 port map( A1 => m3_3, A2 => 
                           z2_temp_3, Z => add_0_root_add_0_root_add_101_n97);
   add_0_root_add_0_root_add_101_U242 : NOR2D1 port map( A1 => m3_6, A2 => 
                           z2_temp_6, Z => add_0_root_add_0_root_add_101_n83);
   add_0_root_add_0_root_add_101_U241 : INVD1 port map( A => 
                           add_0_root_add_0_root_add_101_n102, Z => 
                           add_0_root_add_0_root_add_101_n100);
   add_0_root_add_0_root_add_101_U240 : AND2DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n185, A2 => 
                           add_0_root_add_0_root_add_101_n107, Z => 
                           z2_next_0_port);
   add_0_root_add_0_root_add_101_U239 : NAN2DL port map( A1 => m3_2, A2 => 
                           z2_temp_2, Z => add_0_root_add_0_root_add_101_n102);
   add_0_root_add_0_root_add_101_U238 : NAN2DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n197, A2 => 
                           add_0_root_add_0_root_add_101_n201, Z => 
                           add_0_root_add_0_root_add_101_n15);
   add_0_root_add_0_root_add_101_U237 : INVDL port map( A => 
                           add_0_root_add_0_root_add_101_n56, Z => 
                           add_0_root_add_0_root_add_101_n54);
   add_0_root_add_0_root_add_101_U236 : INVDL port map( A => 
                           add_0_root_add_0_root_add_101_n55, Z => 
                           add_0_root_add_0_root_add_101_n53);
   add_0_root_add_0_root_add_101_U235 : NAN2DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n53, A2 => 
                           add_0_root_add_0_root_add_101_n56, Z => 
                           add_0_root_add_0_root_add_101_n7);
   add_0_root_add_0_root_add_101_U234 : NOR2D2 port map( A1 => m3_13, A2 => 
                           z2_temp_13, Z => add_0_root_add_0_root_add_101_n34);
   add_0_root_add_0_root_add_101_U233 : NAN2D1 port map( A1 => m3_11, A2 => 
                           z2_temp_11, Z => add_0_root_add_0_root_add_101_n51);
   add_0_root_add_0_root_add_101_U232 : NOR2D2 port map( A1 => m3_11, A2 => 
                           z2_temp_11, Z => add_0_root_add_0_root_add_101_n199)
                           ;
   add_0_root_add_0_root_add_101_U231 : NAN2D2 port map( A1 => m3_10, A2 => 
                           z2_temp_10, Z => add_0_root_add_0_root_add_101_n56);
   add_0_root_add_0_root_add_101_U230 : NOR2D2 port map( A1 => 
                           add_0_root_add_0_root_add_101_n55, A2 => 
                           add_0_root_add_0_root_add_101_n50, Z => 
                           add_0_root_add_0_root_add_101_n44);
   add_0_root_add_0_root_add_101_U229 : NAN2D1 port map( A1 => m3_6, A2 => 
                           z2_temp_6, Z => add_0_root_add_0_root_add_101_n84);
   add_0_root_add_0_root_add_101_U228 : NAN2D2 port map( A1 => m3_0, A2 => 
                           z2_temp_0, Z => add_0_root_add_0_root_add_101_n107);
   add_0_root_add_0_root_add_101_U227 : EXNOR2DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n15, A2 => 
                           add_0_root_add_0_root_add_101_n103, Z => 
                           z2_next_2_port);
   add_0_root_add_0_root_add_101_U226 : INVDL port map( A => 
                           add_0_root_add_0_root_add_101_n82, Z => 
                           add_0_root_add_0_root_add_101_net11959);
   add_0_root_add_0_root_add_101_U225 : BUFDL port map( A => 
                           add_0_root_add_0_root_add_101_n179, Z => 
                           add_0_root_add_0_root_add_101_n198);
   add_0_root_add_0_root_add_101_U224 : NAN2D1 port map( A1 => m3_12, A2 => 
                           z2_temp_12, Z => add_0_root_add_0_root_add_101_n42);
   add_0_root_add_0_root_add_101_U223 : INVDL port map( A => 
                           add_0_root_add_0_root_add_101_n100, Z => 
                           add_0_root_add_0_root_add_101_n197);
   add_0_root_add_0_root_add_101_U222 : INVDL port map( A => 
                           add_0_root_add_0_root_add_101_n6, Z => 
                           add_0_root_add_0_root_add_101_n194);
   add_0_root_add_0_root_add_101_U221 : NAN2D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n196, A2 => 
                           add_0_root_add_0_root_add_101_n195, Z => 
                           z2_next_11_port);
   add_0_root_add_0_root_add_101_U220 : NAN2DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n194, A2 => 
                           add_0_root_add_0_root_add_101_n52, Z => 
                           add_0_root_add_0_root_add_101_n195);
   add_0_root_add_0_root_add_101_U219 : EXNOR2DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n27, A2 => 
                           add_0_root_add_0_root_add_101_net12169, Z => 
                           z2_next_14_port);
   add_0_root_add_0_root_add_101_U218 : AOI21DL port map( A1 => 
                           add_0_root_add_0_root_add_101_net9993, A2 => 
                           add_0_root_add_0_root_add_101_n28, B => 
                           add_0_root_add_0_root_add_101_n29, Z => 
                           add_0_root_add_0_root_add_101_n27);
   add_0_root_add_0_root_add_101_U217 : INVD1 port map( A => 
                           add_0_root_add_0_root_add_101_net12354, Z => 
                           add_0_root_add_0_root_add_101_net12355);
   add_0_root_add_0_root_add_101_U216 : NAN2M1DL port map( A1 => 
                           add_0_root_add_0_root_add_101_net12355, A2 => 
                           add_0_root_add_0_root_add_101_n70, Z => 
                           add_0_root_add_0_root_add_101_n9);
   add_0_root_add_0_root_add_101_U215 : INVDL port map( A => 
                           add_0_root_add_0_root_add_101_n84, Z => 
                           add_0_root_add_0_root_add_101_n82);
   add_0_root_add_0_root_add_101_U214 : NAN2M1DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n92, A2 => 
                           add_0_root_add_0_root_add_101_n93, Z => 
                           add_0_root_add_0_root_add_101_n13);
   add_0_root_add_0_root_add_101_U213 : OAI21DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n94, A2 => 
                           add_0_root_add_0_root_add_101_n92, B => 
                           add_0_root_add_0_root_add_101_n93, Z => 
                           add_0_root_add_0_root_add_101_n91);
   add_0_root_add_0_root_add_101_U212 : NAN2M1DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n89, A2 => 
                           add_0_root_add_0_root_add_101_n90, Z => 
                           add_0_root_add_0_root_add_101_n12);
   add_0_root_add_0_root_add_101_U211 : BUFDL port map( A => 
                           add_0_root_add_0_root_add_101_n182, Z => 
                           add_0_root_add_0_root_add_101_net12025);
   add_0_root_add_0_root_add_101_U210 : NOR2D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n92, A2 => 
                           add_0_root_add_0_root_add_101_n89, Z => 
                           add_0_root_add_0_root_add_101_n87);
   add_0_root_add_0_root_add_101_U209 : NOR2M1DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n44, A2 => 
                           add_0_root_add_0_root_add_101_n39, Z => 
                           add_0_root_add_0_root_add_101_n37);
   add_0_root_add_0_root_add_101_U208 : INVDL port map( A => 
                           add_0_root_add_0_root_add_101_n83, Z => 
                           add_0_root_add_0_root_add_101_n81);
   add_0_root_add_0_root_add_101_U207 : INVDL port map( A => 
                           add_0_root_add_0_root_add_101_n78, Z => 
                           add_0_root_add_0_root_add_101_n116);
   add_0_root_add_0_root_add_101_U206 : NOR2M1DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n72, A2 => 
                           add_0_root_add_0_root_add_101_net12355, Z => 
                           add_0_root_add_0_root_add_101_n65);
   add_0_root_add_0_root_add_101_U205 : AOI21D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n85, A2 => 
                           add_0_root_add_0_root_add_101_n72, B => 
                           add_0_root_add_0_root_add_101_n184, Z => 
                           add_0_root_add_0_root_add_101_n71);
   add_0_root_add_0_root_add_101_U204 : NOR2D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n78, A2 => 
                           add_0_root_add_0_root_add_101_n83, Z => 
                           add_0_root_add_0_root_add_101_n72);
   add_0_root_add_0_root_add_101_U203 : NAN2DL port map( A1 => z2_temp_9, A2 =>
                           m3_9, Z => add_0_root_add_0_root_add_101_n63);
   add_0_root_add_0_root_add_101_U202 : NAN2D1 port map( A1 => m3_8, A2 => 
                           z2_temp_8, Z => add_0_root_add_0_root_add_101_n70);
   add_0_root_add_0_root_add_101_U201 : NAN2M1DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n62, A2 => 
                           add_0_root_add_0_root_add_101_n63, Z => 
                           add_0_root_add_0_root_add_101_n8);
   add_0_root_add_0_root_add_101_U200 : OAI21D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n70, A2 => 
                           add_0_root_add_0_root_add_101_n62, B => 
                           add_0_root_add_0_root_add_101_n63, Z => 
                           add_0_root_add_0_root_add_101_n61);
   add_0_root_add_0_root_add_101_U199 : INVDL port map( A => 
                           add_0_root_add_0_root_add_101_n67, Z => 
                           add_0_root_add_0_root_add_101_net12354);
   add_0_root_add_0_root_add_101_U198 : NOR2D2 port map( A1 => 
                           add_0_root_add_0_root_add_101_n62, A2 => 
                           add_0_root_add_0_root_add_101_n67, Z => 
                           add_0_root_add_0_root_add_101_n60);
   add_0_root_add_0_root_add_101_U197 : NAN2M1DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n34, A2 => 
                           add_0_root_add_0_root_add_101_n35, Z => 
                           add_0_root_add_0_root_add_101_n4);
   add_0_root_add_0_root_add_101_U196 : NAN2M1DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n39, A2 => 
                           add_0_root_add_0_root_add_101_n42, Z => 
                           add_0_root_add_0_root_add_101_n5);
   add_0_root_add_0_root_add_101_U195 : OAI21M10DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n45, A2 => 
                           add_0_root_add_0_root_add_101_n39, B => 
                           add_0_root_add_0_root_add_101_n42, Z => 
                           add_0_root_add_0_root_add_101_n38);
   add_0_root_add_0_root_add_101_U194 : INVDL port map( A => 
                           add_0_root_add_0_root_add_101_n73, Z => 
                           add_0_root_add_0_root_add_101_n75);
   add_0_root_add_0_root_add_101_U193 : NAN2D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n60, A2 => 
                           add_0_root_add_0_root_add_101_n72, Z => 
                           add_0_root_add_0_root_add_101_n58);
   add_0_root_add_0_root_add_101_U192 : OAI21D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n180, A2 => 
                           add_0_root_add_0_root_add_101_n190, B => 
                           add_0_root_add_0_root_add_101_n59, Z => 
                           add_0_root_add_0_root_add_101_net9993);
   add_0_root_add_0_root_add_101_U191 : INVDL port map( A => 
                           add_0_root_add_0_root_add_101_n30, Z => 
                           add_0_root_add_0_root_add_101_n28);
   add_0_root_add_0_root_add_101_U190 : NAN2D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n44, A2 => 
                           add_0_root_add_0_root_add_101_n32, Z => 
                           add_0_root_add_0_root_add_101_n30);
   add_0_root_add_0_root_add_101_U189 : AND2D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n109, A2 => 
                           add_0_root_add_0_root_add_101_n26, Z => 
                           add_0_root_add_0_root_add_101_net12169);
   add_0_root_add_0_root_add_101_U188 : NAN2DL port map( A1 => m3_14, A2 => 
                           z2_temp_14, Z => add_0_root_add_0_root_add_101_n26);
   add_0_root_add_0_root_add_101_U187 : INVDL port map( A => 
                           add_0_root_add_0_root_add_101_n23, Z => 
                           add_0_root_add_0_root_add_101_n109);
   add_0_root_add_0_root_add_101_U186 : NOR2D1 port map( A1 => m3_14, A2 => 
                           z2_temp_14, Z => add_0_root_add_0_root_add_101_n23);
   add_0_root_add_0_root_add_101_U185 : OAI21D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n42, A2 => 
                           add_0_root_add_0_root_add_101_n34, B => 
                           add_0_root_add_0_root_add_101_n35, Z => 
                           add_0_root_add_0_root_add_101_n33);
   add_0_root_add_0_root_add_101_U184 : INVDL port map( A => 
                           add_0_root_add_0_root_add_101_n31, Z => 
                           add_0_root_add_0_root_add_101_n29);
   add_0_root_add_0_root_add_101_U183 : AOI21D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n60, A2 => 
                           add_0_root_add_0_root_add_101_n73, B => 
                           add_0_root_add_0_root_add_101_n61, Z => 
                           add_0_root_add_0_root_add_101_net11588);
   add_0_root_add_0_root_add_101_U182 : NOR2DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n30, A2 => 
                           add_0_root_add_0_root_add_101_n23, Z => 
                           add_0_root_add_0_root_add_101_n21);
   add_0_root_add_0_root_add_101_U181 : AOI21DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n21, A2 => 
                           add_0_root_add_0_root_add_101_n1, B => 
                           add_0_root_add_0_root_add_101_n22, Z => 
                           add_0_root_add_0_root_add_101_n20);
   add_0_root_add_0_root_add_101_U180 : OR2D1 port map( A1 => m3_15, A2 => 
                           z2_temp_15, Z => add_0_root_add_0_root_add_101_n192)
                           ;
   add_0_root_add_0_root_add_101_U179 : AND2D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n192, A2 => 
                           add_0_root_add_0_root_add_101_n19, Z => 
                           add_0_root_add_0_root_add_101_net11559);
   add_0_root_add_0_root_add_101_U178 : EXNOR2DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n20, A2 => 
                           add_0_root_add_0_root_add_101_net11559, Z => 
                           z2_next_15_port);
   add_0_root_add_0_root_add_101_U177 : BUFDL port map( A => 
                           add_0_root_add_0_root_add_101_n45, Z => 
                           add_0_root_add_0_root_add_101_n191);
   add_0_root_add_0_root_add_101_U176 : NAN2D1 port map( A1 => m3_1, A2 => 
                           z2_temp_1, Z => add_0_root_add_0_root_add_101_n105);
   add_0_root_add_0_root_add_101_U175 : NAN2M1D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n104, A2 => 
                           add_0_root_add_0_root_add_101_n105, Z => 
                           add_0_root_add_0_root_add_101_n16);
   add_0_root_add_0_root_add_101_U174 : AOI21DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n87, A2 => 
                           add_0_root_add_0_root_add_101_n182, B => 
                           add_0_root_add_0_root_add_101_n88, Z => 
                           add_0_root_add_0_root_add_101_n190);
   add_0_root_add_0_root_add_101_U173 : INVD1 port map( A => 
                           add_0_root_add_0_root_add_101_n52, Z => 
                           add_0_root_add_0_root_add_101_n193);
   add_0_root_add_0_root_add_101_U172 : NAN2D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n193, A2 => 
                           add_0_root_add_0_root_add_101_n6, Z => 
                           add_0_root_add_0_root_add_101_n196);
   add_0_root_add_0_root_add_101_U171 : NOR2D2 port map( A1 => m3_1, A2 => 
                           z2_temp_1, Z => add_0_root_add_0_root_add_101_n104);
   add_0_root_add_0_root_add_101_U170 : NAN2M1D1 port map( A1 => m3_2, A2 => 
                           add_0_root_add_0_root_add_101_n188, Z => 
                           add_0_root_add_0_root_add_101_n201);
   add_0_root_add_0_root_add_101_U169 : AND2DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n116, A2 => 
                           add_0_root_add_0_root_add_101_n79, Z => 
                           add_0_root_add_0_root_add_101_n187);
   add_0_root_add_0_root_add_101_U168 : EXNOR2DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n80, A2 => 
                           add_0_root_add_0_root_add_101_n187, Z => 
                           z2_next_7_port);
   add_0_root_add_0_root_add_101_U167 : AOI21DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n85, A2 => 
                           add_0_root_add_0_root_add_101_n81, B => 
                           add_0_root_add_0_root_add_101_n82, Z => 
                           add_0_root_add_0_root_add_101_n80);
   add_0_root_add_0_root_add_101_U166 : NAN2D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n81, A2 => 
                           add_0_root_add_0_root_add_101_net11959, Z => 
                           add_0_root_add_0_root_add_101_n186);
   add_0_root_add_0_root_add_101_U165 : EXNOR2DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n85, A2 => 
                           add_0_root_add_0_root_add_101_n186, Z => 
                           z2_next_6_port);
   add_0_root_add_0_root_add_101_U164 : INVDL port map( A => 
                           add_0_root_add_0_root_add_101_net12025, Z => 
                           add_0_root_add_0_root_add_101_n94);
   add_0_root_add_0_root_add_101_U163 : EXNOR2D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_net12025, A2 => 
                           add_0_root_add_0_root_add_101_n13, Z => 
                           z2_next_4_port);
   add_0_root_add_0_root_add_101_U162 : NAN2M1DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n96, A2 => 
                           add_0_root_add_0_root_add_101_n97, Z => 
                           add_0_root_add_0_root_add_101_n14);
   add_0_root_add_0_root_add_101_U161 : EXOR2D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n198, A2 => 
                           add_0_root_add_0_root_add_101_n14, Z => 
                           z2_next_3_port);
   add_0_root_add_0_root_add_101_U160 : NAN2D1 port map( A1 => m3_15, A2 => 
                           z2_temp_15, Z => add_0_root_add_0_root_add_101_n19);
   add_0_root_add_0_root_add_101_U159 : INVD1 port map( A => z2_temp_2, Z => 
                           add_0_root_add_0_root_add_101_n188);
   add_0_root_add_0_root_add_101_U158 : NAN2M1DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n199, A2 => 
                           add_0_root_add_0_root_add_101_n51, Z => 
                           add_0_root_add_0_root_add_101_n6);
   add_0_root_add_0_root_add_101_U157 : AOI21D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n87, A2 => 
                           add_0_root_add_0_root_add_101_n95, B => 
                           add_0_root_add_0_root_add_101_n88, Z => 
                           add_0_root_add_0_root_add_101_n189);
   add_0_root_add_0_root_add_101_U156 : OR2DL port map( A1 => m3_0, A2 => 
                           z2_temp_0, Z => add_0_root_add_0_root_add_101_n185);
   add_0_root_add_0_root_add_101_U155 : OAI21DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n78, A2 => 
                           add_0_root_add_0_root_add_101_n84, B => 
                           add_0_root_add_0_root_add_101_n79, Z => 
                           add_0_root_add_0_root_add_101_n184);
   add_0_root_add_0_root_add_101_U154 : AO21DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n85, A2 => 
                           add_0_root_add_0_root_add_101_n65, B => 
                           add_0_root_add_0_root_add_101_n66, Z => 
                           add_0_root_add_0_root_add_101_n183);
   add_0_root_add_0_root_add_101_U153 : EXNOR2DL port map( A1 => 
                           add_0_root_add_0_root_add_101_n183, A2 => 
                           add_0_root_add_0_root_add_101_n8, Z => 
                           z2_next_9_port);
   add_0_root_add_0_root_add_101_U152 : AOI21D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_net9993, A2 => 
                           add_0_root_add_0_root_add_101_n53, B => 
                           add_0_root_add_0_root_add_101_n54, Z => 
                           add_0_root_add_0_root_add_101_n52);
   add_0_root_add_0_root_add_101_U151 : EXNOR2DL port map( A1 => 
                           add_0_root_add_0_root_add_101_net9993, A2 => 
                           add_0_root_add_0_root_add_101_n7, Z => 
                           z2_next_10_port);
   add_0_root_add_0_root_add_101_U150 : INVDL port map( A => 
                           add_0_root_add_0_root_add_101_n189, Z => 
                           add_0_root_add_0_root_add_101_n85);
   add_0_root_add_0_root_add_101_U149 : NOR2D2 port map( A1 => 
                           add_0_root_add_0_root_add_101_n39, A2 => 
                           add_0_root_add_0_root_add_101_n34, Z => 
                           add_0_root_add_0_root_add_101_n32);
   add_0_root_add_0_root_add_101_U148 : NAN2D2 port map( A1 => m3_4, A2 => 
                           z2_temp_4, Z => add_0_root_add_0_root_add_101_n93);
   add_0_root_add_0_root_add_101_U147 : OAI21D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n179, A2 => 
                           add_0_root_add_0_root_add_101_n96, B => 
                           add_0_root_add_0_root_add_101_n97, Z => 
                           add_0_root_add_0_root_add_101_n182);
   add_0_root_add_0_root_add_101_U146 : INVBD32 port map( A => z2_temp_11, Z =>
                           add_0_root_add_0_root_add_101_n181);
   add_0_root_add_0_root_add_101_U145 : NOR2M1D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n181, A2 => m3_11, Z 
                           => add_0_root_add_0_root_add_101_n50);
   add_0_root_add_0_root_add_101_U144 : NAN2D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n60, A2 => 
                           add_0_root_add_0_root_add_101_n72, Z => 
                           add_0_root_add_0_root_add_101_n180);
   add_0_root_add_0_root_add_101_U143 : AOI21D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n103, A2 => 
                           add_0_root_add_0_root_add_101_n201, B => 
                           add_0_root_add_0_root_add_101_n100, Z => 
                           add_0_root_add_0_root_add_101_n179);
   add_0_root_add_0_root_add_101_U10 : OAI21D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n31, A2 => 
                           add_0_root_add_0_root_add_101_n23, B => 
                           add_0_root_add_0_root_add_101_n26, Z => 
                           add_0_root_add_0_root_add_101_n22);
   add_0_root_add_0_root_add_101_U60 : OAI21D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n58, A2 => 
                           add_0_root_add_0_root_add_101_n189, B => 
                           add_0_root_add_0_root_add_101_net11588, Z => 
                           add_0_root_add_0_root_add_101_n1);
   add_0_root_add_0_root_add_101_U40 : AOI21D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n1, A2 => 
                           add_0_root_add_0_root_add_101_n44, B => 
                           add_0_root_add_0_root_add_101_n191, Z => 
                           add_0_root_add_0_root_add_101_n43);
   add_0_root_add_0_root_add_101_U30 : AOI21D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n1, A2 => 
                           add_0_root_add_0_root_add_101_n37, B => 
                           add_0_root_add_0_root_add_101_n38, Z => 
                           add_0_root_add_0_root_add_101_n36);
   add_0_root_add_0_root_add_101_U22 : AOI21D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n32, A2 => 
                           add_0_root_add_0_root_add_101_n45, B => 
                           add_0_root_add_0_root_add_101_n33, Z => 
                           add_0_root_add_0_root_add_101_n31);
   add_0_root_add_0_root_add_101_U62 : AOI21D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n60, A2 => 
                           add_0_root_add_0_root_add_101_n73, B => 
                           add_0_root_add_0_root_add_101_n61, Z => 
                           add_0_root_add_0_root_add_101_n59);
   add_0_root_add_0_root_add_101_U77 : NOR2D2 port map( A1 => m3_8, A2 => 
                           z2_temp_8, Z => add_0_root_add_0_root_add_101_n67);
   add_0_root_add_0_root_add_101_U67 : NOR2D2 port map( A1 => m3_9, A2 => 
                           z2_temp_9, Z => add_0_root_add_0_root_add_101_n62);
   add_0_root_add_0_root_add_101_U86 : OAI21D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n78, A2 => 
                           add_0_root_add_0_root_add_101_n84, B => 
                           add_0_root_add_0_root_add_101_n79, Z => 
                           add_0_root_add_0_root_add_101_n73);
   add_0_root_add_0_root_add_101_U103 : OAI21D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n89, A2 => 
                           add_0_root_add_0_root_add_101_n93, B => 
                           add_0_root_add_0_root_add_101_n90, Z => 
                           add_0_root_add_0_root_add_101_n88);
   add_0_root_add_0_root_add_101_U130 : OAI21D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n104, A2 => 
                           add_0_root_add_0_root_add_101_n107, B => 
                           add_0_root_add_0_root_add_101_n105, Z => 
                           add_0_root_add_0_root_add_101_n103);
   add_0_root_add_0_root_add_101_U129 : EXOR2D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n16, A2 => 
                           add_0_root_add_0_root_add_101_n107, Z => 
                           z2_next_1_port);
   add_0_root_add_0_root_add_101_U122 : AOI21D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n103, A2 => 
                           add_0_root_add_0_root_add_101_n201, B => 
                           add_0_root_add_0_root_add_101_n100, Z => 
                           add_0_root_add_0_root_add_101_n98);
   add_0_root_add_0_root_add_101_U119 : NOR2D2 port map( A1 => m3_3, A2 => 
                           z2_temp_3, Z => add_0_root_add_0_root_add_101_n96);
   add_0_root_add_0_root_add_101_U116 : OAI21D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n98, A2 => 
                           add_0_root_add_0_root_add_101_n96, B => 
                           add_0_root_add_0_root_add_101_n97, Z => 
                           add_0_root_add_0_root_add_101_n95);
   add_0_root_add_0_root_add_101_U112 : NOR2D2 port map( A1 => m3_4, A2 => 
                           z2_temp_4, Z => add_0_root_add_0_root_add_101_n92);
   add_0_root_add_0_root_add_101_U106 : NOR2D2 port map( A1 => m3_5, A2 => 
                           z2_temp_5, Z => add_0_root_add_0_root_add_101_n89);
   add_0_root_add_0_root_add_101_U99 : EXNOR2D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n91, A2 => 
                           add_0_root_add_0_root_add_101_n12, Z => 
                           z2_next_5_port);
   add_0_root_add_0_root_add_101_U89 : NOR2D2 port map( A1 => m3_7, A2 => 
                           z2_temp_7, Z => add_0_root_add_0_root_add_101_n78);
   add_0_root_add_0_root_add_101_U69 : EXOR2D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n71, A2 => 
                           add_0_root_add_0_root_add_101_n9, Z => 
                           z2_next_8_port);
   add_0_root_add_0_root_add_101_U46 : OAI21D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n199, A2 => 
                           add_0_root_add_0_root_add_101_n56, B => 
                           add_0_root_add_0_root_add_101_n51, Z => 
                           add_0_root_add_0_root_add_101_n45);
   add_0_root_add_0_root_add_101_U37 : NOR2D2 port map( A1 => m3_12, A2 => 
                           z2_temp_12, Z => add_0_root_add_0_root_add_101_n39);
   add_0_root_add_0_root_add_101_U29 : EXOR2D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n43, A2 => 
                           add_0_root_add_0_root_add_101_n5, Z => 
                           z2_next_12_port);
   add_0_root_add_0_root_add_101_U17 : EXOR2D1 port map( A1 => 
                           add_0_root_add_0_root_add_101_n36, A2 => 
                           add_0_root_add_0_root_add_101_n4, Z => 
                           z2_next_13_port);
   add_99_U246 : AND2D1 port map( A1 => add_99_n184, A2 => add_99_n19, Z => 
                           add_99_n209);
   add_99_U245 : EXNOR2D1 port map( A1 => add_99_n20, A2 => add_99_n209, Z => 
                           z1_next_15_port);
   add_99_U244 : AND2DL port map( A1 => add_99_n110, A2 => add_99_n35, Z => 
                           add_99_n208);
   add_99_U243 : EXNOR2DL port map( A1 => add_99_n36, A2 => add_99_n208, Z => 
                           z1_next_13_port);
   add_99_U242 : AND2DL port map( A1 => add_99_n112, A2 => add_99_n51, Z => 
                           add_99_n207);
   add_99_U241 : EXNOR2DL port map( A1 => add_99_n52, A2 => add_99_n207, Z => 
                           z1_next_11_port);
   add_99_U240 : OAI21D1 port map( A1 => add_99_n58, A2 => add_99_n86, B => 
                           add_99_n59, Z => add_99_n206);
   add_99_U239 : INVDL port map( A => add_99_n73, Z => add_99_n75);
   add_99_U238 : INVDL port map( A => add_99_n45, Z => add_99_n47);
   add_99_U237 : OAI21DL port map( A1 => add_99_n75, A2 => add_99_n194, B => 
                           add_99_n70, Z => add_99_n66);
   add_99_U236 : INVDL port map( A => add_99_n179, Z => add_99_n116);
   add_99_U235 : NOR2D1 port map( A1 => add_99_n78, A2 => add_99_n83, Z => 
                           add_99_n72);
   add_99_U234 : AOI21DL port map( A1 => add_99_n206, A2 => add_99_n37, B => 
                           add_99_n38, Z => add_99_n36);
   add_99_U233 : AOI21DL port map( A1 => add_99_n21, A2 => add_99_n206, B => 
                           add_99_n22, Z => add_99_n20);
   add_99_U232 : OAI21DL port map( A1 => add_99_n62, A2 => add_99_n70, B => 
                           add_99_n63, Z => add_99_n61);
   add_99_U231 : INVDL port map( A => add_99_n31, Z => add_99_n29);
   add_99_U230 : NAN2DL port map( A1 => add_99_n116, A2 => add_99_n79, Z => 
                           add_99_n10);
   add_99_U229 : NAN2D1 port map( A1 => m5_15, A2 => m4_15, Z => add_99_n19);
   add_99_U228 : NAN2D1 port map( A1 => m5_12, A2 => m4_12, Z => add_99_n42);
   add_99_U227 : NOR2D1 port map( A1 => m5_1, A2 => m4_1, Z => add_99_n104);
   add_99_U226 : NOR2M1DL port map( A1 => add_99_n44, A2 => add_99_n192, Z => 
                           add_99_n37);
   add_99_U225 : NAN2D1 port map( A1 => m4_3, A2 => m5_3, Z => add_99_n97);
   add_99_U224 : NOR2D1 port map( A1 => m5_10, A2 => m4_10, Z => add_99_n55);
   add_99_U223 : NOR2DL port map( A1 => add_99_n30, A2 => add_99_n23, Z => 
                           add_99_n21);
   add_99_U222 : OR2D1 port map( A1 => m5_2, A2 => m4_2, Z => add_99_n205);
   add_99_U221 : INVDL port map( A => add_99_n34, Z => add_99_n110);
   add_99_U220 : INVDL port map( A => add_99_n23, Z => add_99_n109);
   add_99_U219 : INVDL port map( A => add_99_n84, Z => add_99_n82);
   add_99_U218 : INVDL port map( A => add_99_n83, Z => add_99_n81);
   add_99_U217 : NAN2DL port map( A1 => add_99_n81, A2 => add_99_n84, Z => 
                           add_99_n11);
   add_99_U216 : NOR2D1 port map( A1 => add_99_n55, A2 => add_99_n50, Z => 
                           add_99_n44);
   add_99_U215 : INVDL port map( A => add_99_n50, Z => add_99_n112);
   add_99_U214 : NOR2D1 port map( A1 => add_99_n92, A2 => add_99_n89, Z => 
                           add_99_n87);
   add_99_U213 : INVDL port map( A => add_99_n30, Z => add_99_n28);
   add_99_U212 : AND2DL port map( A1 => add_99_n183, A2 => add_99_n107, Z => 
                           z1_next_0_port);
   add_99_U211 : NAN2D1 port map( A1 => m5_14, A2 => m4_14, Z => add_99_n26);
   add_99_U210 : NAN2M1DL port map( A1 => add_99_n104, A2 => add_99_n105, Z => 
                           add_99_n16);
   add_99_U209 : NAN2M1DL port map( A1 => add_99_n39, A2 => add_99_n42, Z => 
                           add_99_n5);
   add_99_U208 : NAN2DL port map( A1 => add_99_n102, A2 => add_99_n205, Z => 
                           add_99_n15);
   add_99_U207 : NAN2M1DL port map( A1 => add_99_n190, A2 => add_99_n97, Z => 
                           add_99_n14);
   add_99_U206 : NAN2M1DL port map( A1 => add_99_n92, A2 => add_99_n93, Z => 
                           add_99_n13);
   add_99_U205 : NAN2M1DL port map( A1 => add_99_n89, A2 => add_99_n90, Z => 
                           add_99_n12);
   add_99_U204 : INVDL port map( A => add_99_n55, Z => add_99_n53);
   add_99_U203 : NAN2M1DL port map( A1 => add_99_n62, A2 => add_99_n63, Z => 
                           add_99_n8);
   add_99_U202 : NAN2M1DL port map( A1 => add_99_n194, A2 => add_99_n70, Z => 
                           add_99_n9);
   add_99_U201 : OAI21DL port map( A1 => add_99_n94, A2 => add_99_n92, B => 
                           add_99_n93, Z => add_99_n91);
   add_99_U200 : NAN2D1 port map( A1 => m5_11, A2 => m4_11, Z => add_99_n51);
   add_99_U199 : INVDL port map( A => add_99_n75, Z => add_99_n203);
   add_99_U198 : AOI21D1 port map( A1 => add_99_n85, A2 => add_99_n182, B => 
                           add_99_n203, Z => add_99_n71);
   add_99_U197 : EXNOR2DL port map( A1 => add_99_n15, A2 => add_99_n103, Z => 
                           z1_next_2_port);
   add_99_U196 : NOR2D2 port map( A1 => add_99_n39, A2 => add_99_n34, Z => 
                           add_99_n32);
   add_99_U195 : NAN2DL port map( A1 => m5_10, A2 => m4_10, Z => add_99_n201);
   add_99_U194 : NAN2D1 port map( A1 => add_99_n72, A2 => add_99_n60, Z => 
                           add_99_n58);
   add_99_U193 : NAN2D2 port map( A1 => m5_0, A2 => m4_0, Z => add_99_n107);
   add_99_U192 : INVD1 port map( A => add_99_n202, Z => add_99_n102);
   add_99_U191 : AND2D1 port map( A1 => m5_2, A2 => m4_2, Z => add_99_n202);
   add_99_U190 : INVDL port map( A => add_99_n206, Z => add_99_n200);
   add_99_U189 : NOR2D1 port map( A1 => add_99_n62, A2 => add_99_n67, Z => 
                           add_99_n60);
   add_99_U188 : INVDL port map( A => add_99_n5, Z => add_99_n197);
   add_99_U187 : NAN2D1 port map( A1 => add_99_n199, A2 => add_99_n198, Z => 
                           z1_next_12_port);
   add_99_U186 : OAI21DL port map( A1 => add_99_n47, A2 => add_99_n192, B => 
                           add_99_n42, Z => add_99_n38);
   add_99_U185 : NOR2D1 port map( A1 => m5_8, A2 => m4_8, Z => add_99_n67);
   add_99_U184 : NOR2DL port map( A1 => m4_8, A2 => add_99_n181, Z => 
                           add_99_n195);
   add_99_U183 : NOR2DL port map( A1 => add_99_n181, A2 => m4_8, Z => 
                           add_99_n194);
   add_99_U182 : AND2D1 port map( A1 => add_99_n109, A2 => add_99_n26, Z => 
                           add_99_n193);
   add_99_U181 : EXNOR2DL port map( A1 => add_99_n27, A2 => add_99_n193, Z => 
                           z1_next_14_port);
   add_99_U180 : NAN2D1 port map( A1 => m5_8, A2 => m4_8, Z => add_99_n70);
   add_99_U179 : NOR2D1 port map( A1 => m5_6, A2 => m4_6, Z => add_99_n83);
   add_99_U178 : NAN2D1 port map( A1 => m5_6, A2 => m4_6, Z => add_99_n84);
   add_99_U177 : OAI21D1 port map( A1 => add_99_n31, A2 => add_99_n23, B => 
                           add_99_n26, Z => add_99_n22);
   add_99_U176 : NAN2D1 port map( A1 => m5_1, A2 => m4_1, Z => add_99_n105);
   add_99_U175 : INVD1 port map( A => add_99_n191, Z => add_99_n192);
   add_99_U174 : INVDL port map( A => add_99_n39, Z => add_99_n191);
   add_99_U173 : NAN2D1 port map( A1 => add_99_n44, A2 => add_99_n32, Z => 
                           add_99_n30);
   add_99_U172 : NOR2DL port map( A1 => m4_3, A2 => m5_3, Z => add_99_n190);
   add_99_U171 : BUFDL port map( A => add_99_n45, Z => add_99_n189);
   add_99_U170 : AOI21DL port map( A1 => add_99_n95, A2 => add_99_n87, B => 
                           add_99_n88, Z => add_99_n86);
   add_99_U169 : AOI21DL port map( A1 => add_99_n95, A2 => add_99_n87, B => 
                           add_99_n88, Z => add_99_n188);
   add_99_U168 : NAN2D1 port map( A1 => m4_13, A2 => m5_13, Z => add_99_n35);
   add_99_U167 : NAN2M1DL port map( A1 => add_99_n187, A2 => m5_9, Z => 
                           add_99_n63);
   add_99_U166 : OA21M20DL port map( A1 => add_99_n206, A2 => add_99_n53, B => 
                           add_99_n201, Z => add_99_n52);
   add_99_U165 : OAI21DL port map( A1 => add_99_n98, A2 => add_99_n96, B => 
                           add_99_n97, Z => add_99_n186);
   add_99_U164 : EXOR2DL port map( A1 => add_99_n14, A2 => add_99_n98, Z => 
                           z1_next_3_port);
   add_99_U163 : NAN2D2 port map( A1 => m5_4, A2 => m4_4, Z => add_99_n93);
   add_99_U162 : AOI21DL port map( A1 => add_99_n1, A2 => add_99_n28, B => 
                           add_99_n29, Z => add_99_n27);
   add_99_U161 : NAN2D1 port map( A1 => add_99_n196, A2 => add_99_n5, Z => 
                           add_99_n199);
   add_99_U160 : NAN2DL port map( A1 => add_99_n43, A2 => add_99_n197, Z => 
                           add_99_n198);
   add_99_U159 : INVD1 port map( A => add_99_n43, Z => add_99_n196);
   add_99_U158 : AND2DL port map( A1 => add_99_n53, A2 => add_99_n201, Z => 
                           add_99_n185);
   add_99_U157 : EXNOR2DL port map( A1 => add_99_n200, A2 => add_99_n185, Z => 
                           z1_next_10_port);
   add_99_U156 : INVD1 port map( A => add_99_n186, Z => add_99_n94);
   add_99_U155 : OR2D1 port map( A1 => m5_15, A2 => m4_15, Z => add_99_n184);
   add_99_U154 : INVD1 port map( A => m4_9, Z => add_99_n187);
   add_99_U153 : NAN2D1 port map( A1 => m5_10, A2 => m4_10, Z => add_99_n56);
   add_99_U152 : OR2DL port map( A1 => m5_0, A2 => m4_0, Z => add_99_n183);
   add_99_U151 : OAI21M20DL port map( A1 => add_99_n95, A2 => add_99_n87, B => 
                           add_99_n180, Z => add_99_n85);
   add_99_U150 : NAN2D1 port map( A1 => m5_7, A2 => m4_7, Z => add_99_n79);
   add_99_U149 : BUFDL port map( A => m5_8, Z => add_99_n181);
   add_99_U148 : BUFDL port map( A => add_99_n72, Z => add_99_n182);
   add_99_U147 : NOR2M1DL port map( A1 => add_99_n72, A2 => add_99_n195, Z => 
                           add_99_n65);
   add_99_U146 : EXNOR2DL port map( A1 => add_99_n85, A2 => add_99_n11, Z => 
                           z1_next_6_port);
   add_99_U145 : NAN2D1 port map( A1 => m5_5, A2 => m4_5, Z => add_99_n90);
   add_99_U144 : OA21DL port map( A1 => add_99_n89, A2 => add_99_n93, B => 
                           add_99_n90, Z => add_99_n180);
   add_99_U143 : BUFDL port map( A => add_99_n78, Z => add_99_n179);
   add_99_U130 : OAI21D1 port map( A1 => add_99_n104, A2 => add_99_n107, B => 
                           add_99_n105, Z => add_99_n103);
   add_99_U129 : EXOR2D1 port map( A1 => add_99_n16, A2 => add_99_n107, Z => 
                           z1_next_1_port);
   add_99_U122 : AOI21D1 port map( A1 => add_99_n205, A2 => add_99_n103, B => 
                           add_99_n202, Z => add_99_n98);
   add_99_U119 : NOR2D2 port map( A1 => m5_3, A2 => m4_3, Z => add_99_n96);
   add_99_U116 : OAI21D1 port map( A1 => add_99_n98, A2 => add_99_n96, B => 
                           add_99_n97, Z => add_99_n95);
   add_99_U112 : NOR2D2 port map( A1 => m5_4, A2 => m4_4, Z => add_99_n92);
   add_99_U108 : EXOR2D1 port map( A1 => add_99_n13, A2 => add_99_n94, Z => 
                           z1_next_4_port);
   add_99_U106 : NOR2D2 port map( A1 => m5_5, A2 => m4_5, Z => add_99_n89);
   add_99_U103 : OAI21D1 port map( A1 => add_99_n89, A2 => add_99_n93, B => 
                           add_99_n90, Z => add_99_n88);
   add_99_U99 : EXNOR2D1 port map( A1 => add_99_n91, A2 => add_99_n12, Z => 
                           z1_next_5_port);
   add_99_U92 : AOI21D1 port map( A1 => add_99_n85, A2 => add_99_n81, B => 
                           add_99_n82, Z => add_99_n80);
   add_99_U89 : NOR2D2 port map( A1 => m5_7, A2 => m4_7, Z => add_99_n78);
   add_99_U86 : OAI21D1 port map( A1 => add_99_n78, A2 => add_99_n84, B => 
                           add_99_n79, Z => add_99_n73);
   add_99_U79 : EXOR2D1 port map( A1 => add_99_n80, A2 => add_99_n10, Z => 
                           z1_next_7_port);
   add_99_U70 : AOI21D1 port map( A1 => add_99_n85, A2 => add_99_n65, B => 
                           add_99_n66, Z => add_99_n64);
   add_99_U69 : EXOR2D1 port map( A1 => add_99_n71, A2 => add_99_n9, Z => 
                           z1_next_8_port);
   add_99_U67 : NOR2D2 port map( A1 => m5_9, A2 => m4_9, Z => add_99_n62);
   add_99_U62 : AOI21D1 port map( A1 => add_99_n60, A2 => add_99_n73, B => 
                           add_99_n61, Z => add_99_n59);
   add_99_U60 : OAI21D1 port map( A1 => add_99_n188, A2 => add_99_n58, B => 
                           add_99_n59, Z => add_99_n1);
   add_99_U59 : EXOR2D1 port map( A1 => add_99_n64, A2 => add_99_n8, Z => 
                           z1_next_9_port);
   add_99_U49 : NOR2D2 port map( A1 => m5_11, A2 => m4_11, Z => add_99_n50);
   add_99_U46 : OAI21D1 port map( A1 => add_99_n50, A2 => add_99_n56, B => 
                           add_99_n51, Z => add_99_n45);
   add_99_U40 : AOI21D1 port map( A1 => add_99_n1, A2 => add_99_n44, B => 
                           add_99_n189, Z => add_99_n43);
   add_99_U37 : NOR2D2 port map( A1 => m5_12, A2 => m4_12, Z => add_99_n39);
   add_99_U27 : NOR2D2 port map( A1 => m5_13, A2 => m4_13, Z => add_99_n34);
   add_99_U24 : OAI21D1 port map( A1 => add_99_n34, A2 => add_99_n42, B => 
                           add_99_n35, Z => add_99_n33);
   add_99_U22 : AOI21D1 port map( A1 => add_99_n32, A2 => add_99_n45, B => 
                           add_99_n33, Z => add_99_n31);
   add_99_U15 : NOR2D2 port map( A1 => m5_14, A2 => m4_14, Z => add_99_n23);
   mult_28_C95_U1276 : EXNOR2DL port map( A1 => y_11_port, A2 => 
                           coeff_memory_17_port, Z => mult_28_C95_n772);
   mult_28_C95_U1275 : EXNOR2DL port map( A1 => y_11_port, A2 => 
                           coeff_memory_27_port, Z => mult_28_C95_n687);
   mult_28_C95_U1274 : EXNOR2DL port map( A1 => mult_28_C95_n914, A2 => 
                           coeff_memory_29_port, Z => mult_28_C95_n670);
   mult_28_C95_U1273 : EXNOR2DL port map( A1 => mult_28_C95_n914, A2 => 
                           coeff_memory_31_port, Z => mult_28_C95_n653);
   mult_28_C95_U1272 : EXNOR2D2 port map( A1 => y_13_port, A2 => 
                           coeff_memory_21_port, Z => mult_28_C95_n736);
   mult_28_C95_U1271 : EXNOR2DL port map( A1 => y_13_port, A2 => 
                           coeff_memory_23_port, Z => mult_28_C95_n719);
   mult_28_C95_U1270 : EXNOR2DL port map( A1 => y_13_port, A2 => 
                           coeff_memory_25_port, Z => mult_28_C95_n702);
   mult_28_C95_U1269 : EXNOR2DL port map( A1 => y_13_port, A2 => 
                           coeff_memory_27_port, Z => mult_28_C95_n685);
   mult_28_C95_U1268 : EXNOR2DL port map( A1 => y_13_port, A2 => 
                           coeff_memory_29_port, Z => mult_28_C95_n668);
   mult_28_C95_U1267 : EXNOR2DL port map( A1 => y_13_port, A2 => 
                           coeff_memory_31_port, Z => mult_28_C95_n651);
   mult_28_C95_U1266 : NAN2DL port map( A1 => mult_28_C95_n288, A2 => 
                           mult_28_C95_n201, Z => mult_28_C95_n67);
   mult_28_C95_U1265 : AOI21DL port map( A1 => mult_28_C95_net12285, A2 => 
                           mult_28_C95_n115, B => mult_28_C95_n116, Z => 
                           mult_28_C95_n114);
   mult_28_C95_U1264 : AOI21DL port map( A1 => mult_28_C95_net12285, A2 => 
                           mult_28_C95_n95, B => mult_28_C95_n96, Z => 
                           mult_28_C95_n94);
   mult_28_C95_U1263 : AOI21DL port map( A1 => mult_28_C95_net12285, A2 => 
                           mult_28_C95_n86, B => mult_28_C95_n87, Z => 
                           mult_28_C95_n85);
   mult_28_C95_U1262 : AOI21D1 port map( A1 => mult_28_C95_net12285, A2 => 
                           mult_28_C95_n141, B => mult_28_C95_n142, Z => 
                           mult_28_C95_n140);
   mult_28_C95_U1261 : OAI21DL port map( A1 => mult_28_C95_n52, A2 => 
                           mult_28_C95_n108, B => mult_28_C95_n109, Z => 
                           mult_28_C95_n107);
   mult_28_C95_U1260 : INVDL port map( A => mult_28_C95_net12183, Z => 
                           mult_28_C95_n129);
   mult_28_C95_U1259 : OAI21DL port map( A1 => mult_28_C95_n52, A2 => 
                           mult_28_C95_n117, B => mult_28_C95_n118, Z => 
                           mult_28_C95_n116);
   mult_28_C95_U1258 : EXNOR2DL port map( A1 => y_14_port, A2 => 
                           coeff_memory_25_port, Z => mult_28_C95_n701);
   mult_28_C95_U1257 : EXNOR2DL port map( A1 => y_14_port, A2 => 
                           coeff_memory_27_port, Z => mult_28_C95_n684);
   mult_28_C95_U1256 : EXNOR2DL port map( A1 => y_14_port, A2 => 
                           coeff_memory_29_port, Z => mult_28_C95_n667);
   mult_28_C95_U1255 : EXNOR2DL port map( A1 => y_14_port, A2 => 
                           coeff_memory_31_port, Z => mult_28_C95_n650);
   mult_28_C95_U1254 : NAN2D1 port map( A1 => mult_28_C95_n388, A2 => 
                           mult_28_C95_n401, Z => mult_28_C95_n196);
   mult_28_C95_U1253 : NOR2D1 port map( A1 => mult_28_C95_n354, A2 => 
                           mult_28_C95_n363, Z => mult_28_C95_n172);
   mult_28_C95_U1252 : NAN3D1 port map( A1 => mult_28_C95_n1011, A2 => 
                           mult_28_C95_n1013, A3 => mult_28_C95_n1012, Z => 
                           mult_28_C95_n363);
   mult_28_C95_U1251 : NAN2DL port map( A1 => mult_28_C95_n368, A2 => 
                           mult_28_C95_net12257, Z => mult_28_C95_n1013);
   mult_28_C95_U1250 : NAN2DL port map( A1 => mult_28_C95_n366, A2 => 
                           mult_28_C95_n368, Z => mult_28_C95_n1012);
   mult_28_C95_U1249 : NAN2DL port map( A1 => mult_28_C95_n366, A2 => 
                           mult_28_C95_net12257, Z => mult_28_C95_n1011);
   mult_28_C95_U1248 : EXNOR2DL port map( A1 => n42, A2 => coeff_memory_25_port
                           , Z => mult_28_C95_n705);
   mult_28_C95_U1247 : EXNOR2DL port map( A1 => n42, A2 => coeff_memory_31_port
                           , Z => mult_28_C95_n654);
   mult_28_C95_U1246 : EXNOR2DL port map( A1 => y_15_port, A2 => 
                           coeff_memory_31_port, Z => mult_28_C95_n649);
   mult_28_C95_U1245 : EXNOR2DL port map( A1 => y_15_port, A2 => 
                           coeff_memory_29_port, Z => mult_28_C95_n666);
   mult_28_C95_U1244 : EXNOR2DL port map( A1 => y_15_port, A2 => 
                           coeff_memory_27_port, Z => mult_28_C95_n683);
   mult_28_C95_U1243 : EXNOR2DL port map( A1 => y_15_port, A2 => 
                           coeff_memory_25_port, Z => mult_28_C95_n700);
   mult_28_C95_U1242 : EXNOR2DL port map( A1 => y_15_port, A2 => 
                           coeff_memory_23_port, Z => mult_28_C95_n717);
   mult_28_C95_U1241 : EXNOR2DL port map( A1 => y_15_port, A2 => 
                           coeff_memory_19_port, Z => mult_28_C95_n751);
   mult_28_C95_U1240 : EXNOR2DL port map( A1 => n38, A2 => coeff_memory_21_port
                           , Z => mult_28_C95_n744);
   mult_28_C95_U1239 : EXNOR2DL port map( A1 => n38, A2 => coeff_memory_31_port
                           , Z => mult_28_C95_n659);
   mult_28_C95_U1238 : EXNOR2DL port map( A1 => n38, A2 => coeff_memory_19_port
                           , Z => mult_28_C95_n761);
   mult_28_C95_U1237 : EXNOR2DL port map( A1 => n38, A2 => coeff_memory_17_port
                           , Z => mult_28_C95_n778);
   mult_28_C95_U1236 : OAI21DL port map( A1 => mult_28_C95_net12183, A2 => 
                           mult_28_C95_n97, B => mult_28_C95_n100, Z => 
                           mult_28_C95_n96);
   mult_28_C95_U1235 : OAI21DL port map( A1 => mult_28_C95_n997, A2 => 
                           mult_28_C95_net12183, B => mult_28_C95_n996, Z => 
                           mult_28_C95_n87);
   mult_28_C95_U1234 : INVDL port map( A => mult_28_C95_n913, Z => 
                           mult_28_C95_n285);
   mult_28_C95_U1233 : AOI21DL port map( A1 => mult_28_C95_n202, A2 => 
                           mult_28_C95_net12127, B => mult_28_C95_net12033, Z 
                           => mult_28_C95_n188);
   mult_28_C95_U1232 : EXNOR2DL port map( A1 => n36, A2 => coeff_memory_23_port
                           , Z => mult_28_C95_n731);
   mult_28_C95_U1231 : EXNOR2DL port map( A1 => n36, A2 => coeff_memory_21_port
                           , Z => mult_28_C95_n748);
   mult_28_C95_U1230 : EXNOR2DL port map( A1 => n36, A2 => coeff_memory_19_port
                           , Z => mult_28_C95_n765);
   mult_28_C95_U1229 : EXNOR2DL port map( A1 => n36, A2 => coeff_memory_17_port
                           , Z => mult_28_C95_n782);
   mult_28_C95_U1228 : INVDL port map( A => mult_28_C95_n201, Z => 
                           mult_28_C95_n199);
   mult_28_C95_U1227 : INVD1 port map( A => coeff_memory_17_port, Z => 
                           mult_28_C95_n832);
   mult_28_C95_U1226 : NAN2D1 port map( A1 => mult_28_C95_n808, A2 => 
                           mult_28_C95_n824, Z => mult_28_C95_n6);
   mult_28_C95_U1225 : NAN2D1 port map( A1 => mult_28_C95_n806, A2 => 
                           mult_28_C95_n16, Z => mult_28_C95_n18);
   mult_28_C95_U1224 : EXNOR2D1 port map( A1 => coeff_memory_19_port, A2 => 
                           coeff_memory_20_port, Z => mult_28_C95_n16);
   mult_28_C95_U1223 : NAN2D1 port map( A1 => mult_28_C95_n807, A2 => 
                           mult_28_C95_n9, Z => mult_28_C95_n12);
   mult_28_C95_U1222 : EXNOR2D1 port map( A1 => coeff_memory_17_port, A2 => 
                           coeff_memory_18_port, Z => mult_28_C95_n9);
   mult_28_C95_U1221 : NAN2D1 port map( A1 => mult_28_C95_n805, A2 => 
                           mult_28_C95_n22, Z => mult_28_C95_n24);
   mult_28_C95_U1220 : EXNOR2D1 port map( A1 => coeff_memory_21_port, A2 => 
                           coeff_memory_22_port, Z => mult_28_C95_n22);
   mult_28_C95_U1219 : NAN2D1 port map( A1 => mult_28_C95_n801, A2 => 
                           mult_28_C95_n46, Z => mult_28_C95_n48);
   mult_28_C95_U1218 : EXNOR2D1 port map( A1 => coeff_memory_29_port, A2 => 
                           coeff_memory_30_port, Z => mult_28_C95_n46);
   mult_28_C95_U1217 : INVD1 port map( A => coeff_memory_19_port, Z => 
                           mult_28_C95_n831);
   mult_28_C95_U1216 : ADHALFDL port map( A => mult_28_C95_n631, B => 
                           mult_28_C95_n519, CO => mult_28_C95_n511, S => 
                           mult_28_C95_n512);
   mult_28_C95_U1215 : INVD1 port map( A => coeff_memory_21_port, Z => 
                           mult_28_C95_n830);
   mult_28_C95_U1214 : ADHALFDL port map( A => mult_28_C95_n614, B => 
                           mult_28_C95_n518, CO => mult_28_C95_n507, S => 
                           mult_28_C95_n508);
   mult_28_C95_U1213 : INVD1 port map( A => coeff_memory_23_port, Z => 
                           mult_28_C95_n829);
   mult_28_C95_U1212 : ADHALFDL port map( A => mult_28_C95_n597, B => 
                           mult_28_C95_n517, CO => mult_28_C95_n499, S => 
                           mult_28_C95_n500);
   mult_28_C95_U1211 : INVD1 port map( A => coeff_memory_25_port, Z => 
                           mult_28_C95_n828);
   mult_28_C95_U1210 : EXNOR2DL port map( A1 => n42, A2 => coeff_memory_17_port
                           , Z => mult_28_C95_n773);
   mult_28_C95_U1209 : INVD1 port map( A => coeff_memory_27_port, Z => 
                           mult_28_C95_n827);
   mult_28_C95_U1208 : EXNOR2DL port map( A1 => n38, A2 => coeff_memory_23_port
                           , Z => mult_28_C95_n727);
   mult_28_C95_U1207 : INVD1 port map( A => coeff_memory_29_port, Z => 
                           mult_28_C95_n826);
   mult_28_C95_U1206 : OR2D1 port map( A1 => mult_28_C95_n305, A2 => 
                           mult_28_C95_n1010, Z => mult_28_C95_n1009);
   mult_28_C95_U1205 : AO21D1 port map( A1 => mult_28_C95_n42, A2 => 
                           mult_28_C95_n40, B => mult_28_C95_n666, Z => 
                           mult_28_C95_n532);
   mult_28_C95_U1204 : INVDL port map( A => mult_28_C95_n309, Z => 
                           mult_28_C95_n310);
   mult_28_C95_U1203 : AND2D1 port map( A1 => mult_28_C95_n648, A2 => 
                           mult_28_C95_n520, Z => mult_28_C95_n1008);
   mult_28_C95_U1202 : NOR2DL port map( A1 => mult_28_C95_n646, A2 => 
                           mult_28_C95_n512, Z => mult_28_C95_n265);
   mult_28_C95_U1201 : NAN2DL port map( A1 => mult_28_C95_n646, A2 => 
                           mult_28_C95_n512, Z => mult_28_C95_n266);
   mult_28_C95_U1200 : AO21D1 port map( A1 => mult_28_C95_n36, A2 => 
                           mult_28_C95_n34, B => mult_28_C95_n683, Z => 
                           mult_28_C95_n548);
   mult_28_C95_U1199 : INVDL port map( A => mult_28_C95_n319, Z => 
                           mult_28_C95_n320);
   mult_28_C95_U1198 : NAN2DL port map( A1 => mult_28_C95_n305, A2 => 
                           mult_28_C95_n1010, Z => mult_28_C95_n84);
   mult_28_C95_U1197 : NAN2D1 port map( A1 => mult_28_C95_n1009, A2 => 
                           mult_28_C95_n84, Z => mult_28_C95_n54);
   mult_28_C95_U1196 : AO21D1 port map( A1 => mult_28_C95_n24, A2 => 
                           mult_28_C95_n22, B => mult_28_C95_n717, Z => 
                           mult_28_C95_n582);
   mult_28_C95_U1195 : INVDL port map( A => mult_28_C95_n333, Z => 
                           mult_28_C95_n334);
   mult_28_C95_U1194 : AO21D1 port map( A1 => mult_28_C95_n30, A2 => 
                           mult_28_C95_n28, B => mult_28_C95_n700, Z => 
                           mult_28_C95_n565);
   mult_28_C95_U1193 : AO21D1 port map( A1 => mult_28_C95_n18, A2 => 
                           mult_28_C95_n16, B => mult_28_C95_n734, Z => 
                           mult_28_C95_n599);
   mult_28_C95_U1192 : NAN2DL port map( A1 => mult_28_C95_n307, A2 => 
                           mult_28_C95_n306, Z => mult_28_C95_n93);
   mult_28_C95_U1191 : NOR2D1 port map( A1 => mult_28_C95_n307, A2 => 
                           mult_28_C95_n306, Z => mult_28_C95_n92);
   mult_28_C95_U1190 : NAN2DL port map( A1 => mult_28_C95_n311, A2 => 
                           mult_28_C95_n308, Z => mult_28_C95_n104);
   mult_28_C95_U1189 : NOR2D1 port map( A1 => mult_28_C95_n311, A2 => 
                           mult_28_C95_n308, Z => mult_28_C95_n103);
   mult_28_C95_U1188 : NAN2D1 port map( A1 => mult_28_C95_n312, A2 => 
                           mult_28_C95_n315, Z => mult_28_C95_n113);
   mult_28_C95_U1187 : NOR2D1 port map( A1 => mult_28_C95_n312, A2 => 
                           mult_28_C95_n315, Z => mult_28_C95_n112);
   mult_28_C95_U1186 : AND2D1 port map( A1 => mult_28_C95_n510, A2 => 
                           mult_28_C95_n645, Z => mult_28_C95_n1005);
   mult_28_C95_U1185 : NAN2DL port map( A1 => mult_28_C95_n506, A2 => 
                           mult_28_C95_n509, Z => mult_28_C95_n258);
   mult_28_C95_U1184 : OR2D1 port map( A1 => mult_28_C95_n502, A2 => 
                           mult_28_C95_n505, Z => mult_28_C95_n1002);
   mult_28_C95_U1183 : AND2D1 port map( A1 => mult_28_C95_n490, A2 => 
                           mult_28_C95_n495, Z => mult_28_C95_n1001);
   mult_28_C95_U1182 : NOR2DL port map( A1 => mult_28_C95_n496, A2 => 
                           mult_28_C95_n501, Z => mult_28_C95_n249);
   mult_28_C95_U1181 : NAN2DL port map( A1 => mult_28_C95_n496, A2 => 
                           mult_28_C95_n501, Z => mult_28_C95_n250);
   mult_28_C95_U1180 : OR2D1 port map( A1 => mult_28_C95_n490, A2 => 
                           mult_28_C95_n495, Z => mult_28_C95_n1000);
   mult_28_C95_U1179 : AND2D1 port map( A1 => mult_28_C95_n482, A2 => 
                           mult_28_C95_n489, Z => mult_28_C95_n999);
   mult_28_C95_U1178 : OR2D1 port map( A1 => mult_28_C95_n97, A2 => 
                           mult_28_C95_n92, Z => mult_28_C95_n997);
   mult_28_C95_U1177 : NAN2D1 port map( A1 => mult_28_C95_n316, A2 => 
                           mult_28_C95_n321, Z => mult_28_C95_n118);
   mult_28_C95_U1176 : NOR2D1 port map( A1 => mult_28_C95_n316, A2 => 
                           mult_28_C95_n321, Z => mult_28_C95_n117);
   mult_28_C95_U1175 : OA21DL port map( A1 => mult_28_C95_n100, A2 => 
                           mult_28_C95_n92, B => mult_28_C95_n93, Z => 
                           mult_28_C95_n996);
   mult_28_C95_U1174 : OR2D1 port map( A1 => mult_28_C95_n464, A2 => 
                           mult_28_C95_n473, Z => mult_28_C95_n995);
   mult_28_C95_U1173 : OR2D1 port map( A1 => mult_28_C95_n322, A2 => 
                           mult_28_C95_n327, Z => mult_28_C95_net11083);
   mult_28_C95_U1172 : NAN2D1 port map( A1 => mult_28_C95_n344, A2 => 
                           mult_28_C95_n353, Z => mult_28_C95_n168);
   mult_28_C95_U1171 : AND2DL port map( A1 => mult_28_C95_n442, A2 => 
                           mult_28_C95_n453, Z => mult_28_C95_n994);
   mult_28_C95_U1170 : OR2D1 port map( A1 => mult_28_C95_n454, A2 => 
                           mult_28_C95_n463, Z => mult_28_C95_n993);
   mult_28_C95_U1169 : AND2D1 port map( A1 => mult_28_C95_n454, A2 => 
                           mult_28_C95_n463, Z => mult_28_C95_n992);
   mult_28_C95_U1168 : NAN2D1 port map( A1 => mult_28_C95_n991, A2 => 
                           mult_28_C95_n998, Z => mult_28_C95_n231);
   mult_28_C95_U1167 : OA21M20D1 port map( A1 => mult_28_C95_n124, A2 => 
                           mult_28_C95_n278, B => mult_28_C95_n113, Z => 
                           mult_28_C95_n109);
   mult_28_C95_U1166 : NOR2D1 port map( A1 => mult_28_C95_n402, A2 => 
                           mult_28_C95_n415, Z => mult_28_C95_n200);
   mult_28_C95_U1165 : OR2D1 port map( A1 => mult_28_C95_n442, A2 => 
                           mult_28_C95_n453, Z => mult_28_C95_n990);
   mult_28_C95_U1164 : NOR2DL port map( A1 => mult_28_C95_n53, A2 => 
                           mult_28_C95_n117, Z => mult_28_C95_n115);
   mult_28_C95_U1163 : NAN2DL port map( A1 => mult_28_C95_n101, A2 => 
                           mult_28_C95_n279, Z => mult_28_C95_n97);
   mult_28_C95_U1162 : NAN2D1 port map( A1 => mult_28_C95_n279, A2 => 
                           mult_28_C95_n278, Z => mult_28_C95_n108);
   mult_28_C95_U1161 : NOR2DL port map( A1 => mult_28_C95_n53, A2 => 
                           mult_28_C95_n997, Z => mult_28_C95_n86);
   mult_28_C95_U1160 : INVDL port map( A => mult_28_C95_n172, Z => 
                           mult_28_C95_n284);
   mult_28_C95_U1159 : NOR2DL port map( A1 => mult_28_C95_n53, A2 => 
                           mult_28_C95_n97, Z => mult_28_C95_n95);
   mult_28_C95_U1158 : OA22DL port map( A1 => mult_28_C95_n650, A2 => 
                           mult_28_C95_n48, B1 => mult_28_C95_n649, B2 => 
                           mult_28_C95_n46, Z => mult_28_C95_n1010);
   mult_28_C95_U1157 : OAI22DL port map( A1 => mult_28_C95_n652, A2 => 
                           mult_28_C95_n48, B1 => mult_28_C95_n651, B2 => 
                           mult_28_C95_n46, Z => mult_28_C95_n523);
   mult_28_C95_U1156 : OAI22DL port map( A1 => mult_28_C95_n653, A2 => 
                           mult_28_C95_n48, B1 => mult_28_C95_n652, B2 => 
                           mult_28_C95_n46, Z => mult_28_C95_n524);
   mult_28_C95_U1155 : OAI22DL port map( A1 => mult_28_C95_n670, A2 => 
                           mult_28_C95_n42, B1 => mult_28_C95_n669, B2 => 
                           mult_28_C95_n40, Z => mult_28_C95_n535);
   mult_28_C95_U1154 : OAI22D1 port map( A1 => mult_28_C95_n754, A2 => 
                           mult_28_C95_n12, B1 => mult_28_C95_n753, B2 => 
                           mult_28_C95_n9, Z => mult_28_C95_n619);
   mult_28_C95_U1153 : AND2DL port map( A1 => mult_28_C95_n647, A2 => 
                           mult_28_C95_n632, Z => mult_28_C95_n1007);
   mult_28_C95_U1152 : OR2DL port map( A1 => mult_28_C95_n510, A2 => 
                           mult_28_C95_n645, Z => mult_28_C95_n1004);
   mult_28_C95_U1151 : NOR2D1 port map( A1 => mult_28_C95_n506, A2 => 
                           mult_28_C95_n509, Z => mult_28_C95_n257);
   mult_28_C95_U1150 : AND2DL port map( A1 => mult_28_C95_n502, A2 => 
                           mult_28_C95_n505, Z => mult_28_C95_n1003);
   mult_28_C95_U1149 : EXNOR2D2 port map( A1 => mult_28_C95_net11025, A2 => 
                           mult_28_C95_n366, Z => mult_28_C95_n364);
   mult_28_C95_U1148 : NOR2DL port map( A1 => mult_28_C95_n112, A2 => 
                           mult_28_C95_n103, Z => mult_28_C95_n101);
   mult_28_C95_U1147 : INVDL port map( A => mult_28_C95_n112, Z => 
                           mult_28_C95_n278);
   mult_28_C95_U1146 : NAN2DL port map( A1 => mult_28_C95_n322, A2 => 
                           mult_28_C95_n327, Z => mult_28_C95_n139);
   mult_28_C95_U1145 : NAN2M1DL port map( A1 => mult_28_C95_n92, A2 => 
                           mult_28_C95_n93, Z => mult_28_C95_n55);
   mult_28_C95_U1144 : AND2DL port map( A1 => mult_28_C95_n278, A2 => 
                           mult_28_C95_n113, Z => mult_28_C95_n988);
   mult_28_C95_U1143 : EXNOR2D2 port map( A1 => mult_28_C95_n114, A2 => 
                           mult_28_C95_n988, Z => m3_12);
   mult_28_C95_U1142 : NAN2M1DL port map( A1 => mult_28_C95_n103, A2 => 
                           mult_28_C95_n104, Z => mult_28_C95_n56);
   mult_28_C95_U1141 : INVDL port map( A => mult_28_C95_n118, Z => 
                           mult_28_C95_n124);
   mult_28_C95_U1140 : INVDL port map( A => mult_28_C95_n117, Z => 
                           mult_28_C95_n279);
   mult_28_C95_U1139 : INVDL port map( A => mult_28_C95_n173, Z => 
                           mult_28_C95_n171);
   mult_28_C95_U1138 : AOI21DL port map( A1 => mult_28_C95_n182, A2 => 
                           mult_28_C95_n202, B => mult_28_C95_n183, Z => 
                           mult_28_C95_n987);
   mult_28_C95_U1137 : EXNOR2D1 port map( A1 => mult_28_C95_n987, A2 => 
                           mult_28_C95_net11172, Z => m3_5);
   mult_28_C95_U1136 : NAN2M1DL port map( A1 => mult_28_C95_net12055, A2 => 
                           mult_28_C95_net11746, Z => mult_28_C95_n65);
   mult_28_C95_U1135 : NAN2DL port map( A1 => mult_28_C95_n284, A2 => 
                           mult_28_C95_net12095, Z => mult_28_C95_n63);
   mult_28_C95_U1134 : AND2DL port map( A1 => mult_28_C95_n283, A2 => 
                           mult_28_C95_n168, Z => mult_28_C95_n989);
   mult_28_C95_U1133 : NOR2DL port map( A1 => mult_28_C95_n53, A2 => 
                           mult_28_C95_n108, Z => mult_28_C95_n106);
   mult_28_C95_U1132 : INVDL port map( A => mult_28_C95_n53, Z => 
                           mult_28_C95_n128);
   mult_28_C95_U1131 : EXNOR2DL port map( A1 => y_2_port, A2 => 
                           coeff_memory_29_port, Z => mult_28_C95_n679);
   mult_28_C95_U1130 : EXNOR2DL port map( A1 => y_2_port, A2 => 
                           coeff_memory_25_port, Z => mult_28_C95_n713);
   mult_28_C95_U1129 : EXNOR2D2 port map( A1 => n42, A2 => coeff_memory_21_port
                           , Z => mult_28_C95_n739);
   mult_28_C95_U1128 : NAN2D2 port map( A1 => mult_28_C95_n402, A2 => 
                           mult_28_C95_n415, Z => mult_28_C95_n201);
   mult_28_C95_U1127 : EXNOR2DL port map( A1 => y_14_port, A2 => 
                           coeff_memory_19_port, Z => mult_28_C95_n752);
   mult_28_C95_U1126 : EXNOR2DL port map( A1 => y_14_port, A2 => 
                           coeff_memory_21_port, Z => mult_28_C95_n735);
   mult_28_C95_U1125 : EXNOR2D2 port map( A1 => y_14_port, A2 => 
                           coeff_memory_17_port, Z => mult_28_C95_n769);
   mult_28_C95_U1124 : EXNOR2D2 port map( A1 => y_6_port, A2 => 
                           coeff_memory_29_port, Z => mult_28_C95_n675);
   mult_28_C95_U1123 : EXNOR2DL port map( A1 => y_6_port, A2 => 
                           coeff_memory_21_port, Z => mult_28_C95_n743);
   mult_28_C95_U1122 : EXNOR2DL port map( A1 => y_9_port, A2 => 
                           coeff_memory_27_port, Z => mult_28_C95_n689);
   mult_28_C95_U1121 : EXNOR2DL port map( A1 => coeff_memory_17_port, A2 => 
                           y_9_port, Z => mult_28_C95_n774);
   mult_28_C95_U1120 : EXNOR2D2 port map( A1 => n38, A2 => coeff_memory_25_port
                           , Z => mult_28_C95_n710);
   mult_28_C95_U1119 : ADFULD1 port map( A => mult_28_C95_n619, B => 
                           mult_28_C95_n437, CI => mult_28_C95_n435, CO => 
                           mult_28_C95_n419, S => mult_28_C95_n420);
   mult_28_C95_U1118 : NAN3D2 port map( A1 => mult_28_C95_n984, A2 => 
                           mult_28_C95_n986, A3 => mult_28_C95_n985, Z => 
                           mult_28_C95_n435);
   mult_28_C95_U1117 : NAN2D1 port map( A1 => mult_28_C95_n449, A2 => 
                           mult_28_C95_n590, Z => mult_28_C95_n986);
   mult_28_C95_U1116 : NAN3D1 port map( A1 => mult_28_C95_net11507, A2 => 
                           mult_28_C95_n983, A3 => mult_28_C95_net11509, Z => 
                           mult_28_C95_n401);
   mult_28_C95_U1115 : NAN2DL port map( A1 => mult_28_C95_n417, A2 => 
                           mult_28_C95_n404, Z => mult_28_C95_n983);
   mult_28_C95_U1114 : NAN3D2 port map( A1 => mult_28_C95_n980, A2 => 
                           mult_28_C95_n981, A3 => mult_28_C95_n982, Z => 
                           mult_28_C95_n403);
   mult_28_C95_U1113 : NAN2D1 port map( A1 => mult_28_C95_n410, A2 => 
                           mult_28_C95_n408, Z => mult_28_C95_n982);
   mult_28_C95_U1112 : NAN2D1 port map( A1 => mult_28_C95_n419, A2 => 
                           mult_28_C95_n408, Z => mult_28_C95_n981);
   mult_28_C95_U1111 : NAN2D1 port map( A1 => mult_28_C95_n419, A2 => 
                           mult_28_C95_n410, Z => mult_28_C95_n980);
   mult_28_C95_U1110 : EXOR3D1 port map( A1 => mult_28_C95_n419, A2 => 
                           mult_28_C95_n410, A3 => mult_28_C95_n408, Z => 
                           mult_28_C95_n404);
   mult_28_C95_U1109 : EXNOR2D2 port map( A1 => y_15_port, A2 => 
                           coeff_memory_17_port, Z => mult_28_C95_n768);
   mult_28_C95_U1108 : EXNOR2DL port map( A1 => y_8_port, A2 => 
                           coeff_memory_25_port, Z => mult_28_C95_n978);
   mult_28_C95_U1107 : EXNOR2DL port map( A1 => y_7_port, A2 => 
                           coeff_memory_21_port, Z => mult_28_C95_n742);
   mult_28_C95_U1106 : EXNOR2DL port map( A1 => coeff_memory_23_port, A2 => 
                           y_14_port, Z => mult_28_C95_n718);
   mult_28_C95_U1105 : EXNOR2DL port map( A1 => y_7_port, A2 => 
                           coeff_memory_31_port, Z => mult_28_C95_n657);
   mult_28_C95_U1104 : EXNOR2DL port map( A1 => y_7_port, A2 => 
                           coeff_memory_19_port, Z => mult_28_C95_n759);
   mult_28_C95_U1103 : EXNOR2DL port map( A1 => y_7_port, A2 => 
                           coeff_memory_17_port, Z => mult_28_C95_n776);
   mult_28_C95_U1102 : OAI22D2 port map( A1 => mult_28_C95_n718, A2 => 
                           mult_28_C95_n24, B1 => mult_28_C95_n717, B2 => 
                           mult_28_C95_n22, Z => mult_28_C95_n583);
   mult_28_C95_U1101 : OAI22DL port map( A1 => mult_28_C95_n701, A2 => 
                           mult_28_C95_n30, B1 => mult_28_C95_n700, B2 => 
                           mult_28_C95_n28, Z => mult_28_C95_n566);
   mult_28_C95_U1100 : OAI22D2 port map( A1 => mult_28_C95_n684, A2 => 
                           mult_28_C95_n36, B1 => mult_28_C95_n683, B2 => 
                           mult_28_C95_n34, Z => mult_28_C95_n549);
   mult_28_C95_U1099 : OAI22DL port map( A1 => mult_28_C95_n668, A2 => 
                           mult_28_C95_n42, B1 => mult_28_C95_n667, B2 => 
                           mult_28_C95_n40, Z => mult_28_C95_n533);
   mult_28_C95_U1098 : EXNOR2DL port map( A1 => y_8_port, A2 => 
                           coeff_memory_19_port, Z => mult_28_C95_n758);
   mult_28_C95_U1097 : EXNOR2DL port map( A1 => y_8_port, A2 => 
                           coeff_memory_17_port, Z => mult_28_C95_n775);
   mult_28_C95_U1096 : EXNOR2DL port map( A1 => y_8_port, A2 => 
                           coeff_memory_29_port, Z => mult_28_C95_n673);
   mult_28_C95_U1095 : ADHALFD2 port map( A => mult_28_C95_n546, B => 
                           mult_28_C95_n514, CO => mult_28_C95_n451, S => 
                           mult_28_C95_n452);
   mult_28_C95_U1094 : EXOR2D4 port map( A1 => mult_28_C95_n188, A2 => 
                           mult_28_C95_n65, Z => m3_4);
   mult_28_C95_U1093 : EXNOR2D2 port map( A1 => y_12_port, A2 => 
                           coeff_memory_23_port, Z => mult_28_C95_n720);
   mult_28_C95_U1092 : EXNOR2D2 port map( A1 => n38, A2 => coeff_memory_29_port
                           , Z => mult_28_C95_n676);
   mult_28_C95_U1091 : EXNOR2DL port map( A1 => y_12_port, A2 => 
                           coeff_memory_31_port, Z => mult_28_C95_n652);
   mult_28_C95_U1090 : EXNOR2DL port map( A1 => y_12_port, A2 => 
                           coeff_memory_29_port, Z => mult_28_C95_n669);
   mult_28_C95_U1089 : EXNOR2DL port map( A1 => y_12_port, A2 => 
                           coeff_memory_27_port, Z => mult_28_C95_n686);
   mult_28_C95_U1088 : EXNOR2DL port map( A1 => y_12_port, A2 => 
                           coeff_memory_25_port, Z => mult_28_C95_n703);
   mult_28_C95_U1087 : EXNOR2DL port map( A1 => y_12_port, A2 => 
                           coeff_memory_19_port, Z => mult_28_C95_n754);
   mult_28_C95_U1086 : EXNOR2DL port map( A1 => y_2_port, A2 => 
                           coeff_memory_27_port, Z => mult_28_C95_n696);
   mult_28_C95_U1085 : EXNOR2DL port map( A1 => y_2_port, A2 => 
                           coeff_memory_31_port, Z => mult_28_C95_n662);
   mult_28_C95_U1084 : OAI22D1 port map( A1 => mult_28_C95_n708, A2 => 
                           mult_28_C95_n30, B1 => mult_28_C95_n978, B2 => 
                           mult_28_C95_n28, Z => mult_28_C95_n573);
   mult_28_C95_U1083 : EXOR2D1 port map( A1 => mult_28_C95_n977, A2 => 
                           mult_28_C95_n588, Z => mult_28_C95_n410);
   mult_28_C95_U1082 : EXOR2D1 port map( A1 => mult_28_C95_n573, A2 => 
                           mult_28_C95_n425, Z => mult_28_C95_n977);
   mult_28_C95_U1081 : EXNOR2DL port map( A1 => y_9_port, A2 => 
                           coeff_memory_23_port, Z => mult_28_C95_n723);
   mult_28_C95_U1080 : EXNOR2DL port map( A1 => y_9_port, A2 => 
                           coeff_memory_21_port, Z => mult_28_C95_n740);
   mult_28_C95_U1079 : EXNOR2D2 port map( A1 => mult_28_C95_n160, A2 => 
                           mult_28_C95_net11662, Z => m3_8);
   mult_28_C95_U1078 : EXNOR2D2 port map( A1 => n42, A2 => coeff_memory_27_port
                           , Z => mult_28_C95_n688);
   mult_28_C95_U1077 : NAN3D2 port map( A1 => mult_28_C95_n974, A2 => 
                           mult_28_C95_n975, A3 => mult_28_C95_n976, Z => 
                           mult_28_C95_n365);
   mult_28_C95_U1076 : NAN2DL port map( A1 => mult_28_C95_n381, A2 => 
                           mult_28_C95_n379, Z => mult_28_C95_n976);
   mult_28_C95_U1075 : NAN2DL port map( A1 => mult_28_C95_n370, A2 => 
                           mult_28_C95_n379, Z => mult_28_C95_n975);
   mult_28_C95_U1074 : NAN2DL port map( A1 => mult_28_C95_n370, A2 => 
                           mult_28_C95_n381, Z => mult_28_C95_n974);
   mult_28_C95_U1073 : EXOR2D1 port map( A1 => mult_28_C95_n370, A2 => 
                           mult_28_C95_n381, Z => mult_28_C95_n973);
   mult_28_C95_U1072 : NAN2DL port map( A1 => mult_28_C95_n616, A2 => 
                           mult_28_C95_n393, Z => mult_28_C95_n972);
   mult_28_C95_U1071 : OAI22D1 port map( A1 => mult_28_C95_n769, A2 => 
                           mult_28_C95_n6, B1 => mult_28_C95_n768, B2 => 
                           mult_28_C95_n824, Z => mult_28_C95_n979);
   mult_28_C95_U1070 : INVD1 port map( A => mult_28_C95_n167, Z => 
                           mult_28_C95_n283);
   mult_28_C95_U1069 : NAN2D1 port map( A1 => mult_28_C95_n430, A2 => 
                           mult_28_C95_n441, Z => mult_28_C95_n210);
   mult_28_C95_U1068 : ADFULD1 port map( A => mult_28_C95_n578, B => 
                           mult_28_C95_n472, CI => mult_28_C95_n593, CO => 
                           mult_28_C95_n469, S => mult_28_C95_n470);
   mult_28_C95_U1067 : NAN3D2 port map( A1 => mult_28_C95_n969, A2 => 
                           mult_28_C95_n971, A3 => mult_28_C95_n970, Z => 
                           mult_28_C95_n457);
   mult_28_C95_U1066 : NAN2D1 port map( A1 => mult_28_C95_n607, A2 => 
                           mult_28_C95_n622, Z => mult_28_C95_n971);
   mult_28_C95_U1065 : NAN2D1 port map( A1 => mult_28_C95_n469, A2 => 
                           mult_28_C95_n622, Z => mult_28_C95_n970);
   mult_28_C95_U1064 : NAN2D1 port map( A1 => mult_28_C95_n469, A2 => 
                           mult_28_C95_n607, Z => mult_28_C95_n969);
   mult_28_C95_U1063 : EXOR3D2 port map( A1 => mult_28_C95_n622, A2 => 
                           mult_28_C95_n469, A3 => mult_28_C95_n607, Z => 
                           mult_28_C95_n458);
   mult_28_C95_U1062 : NAN3D1 port map( A1 => mult_28_C95_n966, A2 => 
                           mult_28_C95_n968, A3 => mult_28_C95_n967, Z => 
                           mult_28_C95_n447);
   mult_28_C95_U1061 : NAN2DL port map( A1 => mult_28_C95_n591, A2 => 
                           mult_28_C95_n461, Z => mult_28_C95_n968);
   mult_28_C95_U1060 : NAN2DL port map( A1 => mult_28_C95_n606, A2 => 
                           mult_28_C95_n591, Z => mult_28_C95_n966);
   mult_28_C95_U1059 : EXOR2D1 port map( A1 => mult_28_C95_n965, A2 => 
                           mult_28_C95_n606, Z => mult_28_C95_n448);
   mult_28_C95_U1058 : EXOR2D1 port map( A1 => mult_28_C95_n461, A2 => 
                           mult_28_C95_n591, Z => mult_28_C95_n965);
   mult_28_C95_U1057 : NAN3D1 port map( A1 => mult_28_C95_n962, A2 => 
                           mult_28_C95_n963, A3 => mult_28_C95_n964, Z => 
                           mult_28_C95_n441);
   mult_28_C95_U1056 : NAN2DL port map( A1 => mult_28_C95_n446, A2 => 
                           mult_28_C95_n444, Z => mult_28_C95_n964);
   mult_28_C95_U1055 : NAN2DL port map( A1 => mult_28_C95_n444, A2 => 
                           mult_28_C95_n455, Z => mult_28_C95_n963);
   mult_28_C95_U1054 : NAN2DL port map( A1 => mult_28_C95_n446, A2 => 
                           mult_28_C95_n455, Z => mult_28_C95_n962);
   mult_28_C95_U1053 : NAN3D2 port map( A1 => mult_28_C95_n959, A2 => 
                           mult_28_C95_n960, A3 => mult_28_C95_n961, Z => 
                           mult_28_C95_n443);
   mult_28_C95_U1052 : NAN2D1 port map( A1 => mult_28_C95_n459, A2 => 
                           mult_28_C95_n448, Z => mult_28_C95_n961);
   mult_28_C95_U1051 : NAN2DL port map( A1 => mult_28_C95_n457, A2 => 
                           mult_28_C95_n448, Z => mult_28_C95_n960);
   mult_28_C95_U1050 : NAN2DL port map( A1 => mult_28_C95_n457, A2 => 
                           mult_28_C95_n459, Z => mult_28_C95_n959);
   mult_28_C95_U1049 : EXOR2D1 port map( A1 => mult_28_C95_n958, A2 => 
                           mult_28_C95_n444, Z => mult_28_C95_n442);
   mult_28_C95_U1048 : EXOR3D1 port map( A1 => mult_28_C95_n457, A2 => 
                           mult_28_C95_n459, A3 => mult_28_C95_n448, Z => 
                           mult_28_C95_n444);
   mult_28_C95_U1047 : OAI22DL port map( A1 => mult_28_C95_n773, A2 => 
                           mult_28_C95_n824, B1 => mult_28_C95_n774, B2 => 
                           mult_28_C95_n6, Z => mult_28_C95_n639);
   mult_28_C95_U1046 : NAN3D1 port map( A1 => mult_28_C95_n955, A2 => 
                           mult_28_C95_n957, A3 => mult_28_C95_n956, Z => 
                           mult_28_C95_n475);
   mult_28_C95_U1045 : NAN2DL port map( A1 => mult_28_C95_n485, A2 => 
                           mult_28_C95_n624, Z => mult_28_C95_n957);
   mult_28_C95_U1044 : NAN2DL port map( A1 => mult_28_C95_n639, A2 => 
                           mult_28_C95_n624, Z => mult_28_C95_n956);
   mult_28_C95_U1043 : NAN2DL port map( A1 => mult_28_C95_n639, A2 => 
                           mult_28_C95_n485, Z => mult_28_C95_n955);
   mult_28_C95_U1042 : EXOR2D1 port map( A1 => mult_28_C95_n954, A2 => 
                           mult_28_C95_n639, Z => mult_28_C95_n476);
   mult_28_C95_U1041 : EXOR2D1 port map( A1 => mult_28_C95_n624, A2 => 
                           mult_28_C95_n485, Z => mult_28_C95_n954);
   mult_28_C95_U1040 : NAN3D1 port map( A1 => mult_28_C95_n951, A2 => 
                           mult_28_C95_n953, A3 => mult_28_C95_n952, Z => 
                           mult_28_C95_n473);
   mult_28_C95_U1039 : NAN2DL port map( A1 => mult_28_C95_n478, A2 => 
                           mult_28_C95_n483, Z => mult_28_C95_n953);
   mult_28_C95_U1038 : NAN2DL port map( A1 => mult_28_C95_n476, A2 => 
                           mult_28_C95_n483, Z => mult_28_C95_n952);
   mult_28_C95_U1037 : NAN2DL port map( A1 => mult_28_C95_n476, A2 => 
                           mult_28_C95_n478, Z => mult_28_C95_n951);
   mult_28_C95_U1036 : EXOR2D1 port map( A1 => mult_28_C95_n950, A2 => 
                           mult_28_C95_n476, Z => mult_28_C95_n474);
   mult_28_C95_U1035 : EXOR2D1 port map( A1 => mult_28_C95_n483, A2 => 
                           mult_28_C95_n478, Z => mult_28_C95_n950);
   mult_28_C95_U1034 : AND2DL port map( A1 => mult_28_C95_n279, A2 => 
                           mult_28_C95_n118, Z => mult_28_C95_n949);
   mult_28_C95_U1033 : EXNOR2D2 port map( A1 => mult_28_C95_n127, A2 => 
                           mult_28_C95_n949, Z => m3_11);
   mult_28_C95_U1032 : EXNOR2D2 port map( A1 => y_6_port, A2 => 
                           coeff_memory_25_port, Z => mult_28_C95_n709);
   mult_28_C95_U1031 : NAN2D1 port map( A1 => mult_28_C95_n943, A2 => 
                           mult_28_C95_n429, Z => mult_28_C95_n207);
   mult_28_C95_U1030 : AND2DL port map( A1 => mult_28_C95_net11083, A2 => 
                           mult_28_C95_n139, Z => mult_28_C95_n948);
   mult_28_C95_U1029 : EXNOR2D2 port map( A1 => mult_28_C95_n140, A2 => 
                           mult_28_C95_n948, Z => m3_10);
   mult_28_C95_U1028 : INVD1 port map( A => mult_28_C95_net11745, Z => 
                           mult_28_C95_net11746);
   mult_28_C95_U1027 : EXNOR2D2 port map( A1 => y_12_port, A2 => 
                           coeff_memory_17_port, Z => mult_28_C95_n771);
   mult_28_C95_U1026 : EXNOR2D2 port map( A1 => mult_28_C95_n105, A2 => 
                           mult_28_C95_n947, Z => m3_13);
   mult_28_C95_U1025 : NAN3D1 port map( A1 => mult_28_C95_n944, A2 => 
                           mult_28_C95_n946, A3 => mult_28_C95_n945, Z => 
                           mult_28_C95_n383);
   mult_28_C95_U1024 : NAN2DL port map( A1 => mult_28_C95_n397, A2 => 
                           mult_28_C95_n556, Z => mult_28_C95_n946);
   mult_28_C95_U1023 : NAN2DL port map( A1 => mult_28_C95_n571, A2 => 
                           mult_28_C95_n556, Z => mult_28_C95_n945);
   mult_28_C95_U1022 : NAN2D1 port map( A1 => mult_28_C95_n571, A2 => 
                           mult_28_C95_n397, Z => mult_28_C95_n944);
   mult_28_C95_U1021 : EXOR2D1 port map( A1 => mult_28_C95_n556, A2 => 
                           mult_28_C95_n397, Z => mult_28_C95_net11829);
   mult_28_C95_U1020 : EXNOR2D2 port map( A1 => y_3_port, A2 => 
                           coeff_memory_27_port, Z => mult_28_C95_n695);
   mult_28_C95_U1019 : EXNOR2D2 port map( A1 => y_3_port, A2 => 
                           coeff_memory_25_port, Z => mult_28_C95_n712);
   mult_28_C95_U1018 : EXNOR2D2 port map( A1 => y_3_port, A2 => 
                           coeff_memory_23_port, Z => mult_28_C95_n729);
   mult_28_C95_U1017 : EXNOR2D2 port map( A1 => y_3_port, A2 => 
                           coeff_memory_21_port, Z => mult_28_C95_n746);
   mult_28_C95_U1016 : EXNOR2DL port map( A1 => y_3_port, A2 => 
                           coeff_memory_19_port, Z => mult_28_C95_n763);
   mult_28_C95_U1015 : EXNOR2D2 port map( A1 => y_3_port, A2 => 
                           coeff_memory_31_port, Z => mult_28_C95_n661);
   mult_28_C95_U1014 : OAI21DL port map( A1 => mult_28_C95_n192, A2 => 
                           mult_28_C95_net12055, B => mult_28_C95_net11746, Z 
                           => mult_28_C95_n183);
   mult_28_C95_U1013 : EXNOR2D2 port map( A1 => y_13_port, A2 => 
                           coeff_memory_17_port, Z => mult_28_C95_n770);
   mult_28_C95_U1012 : EXNOR2DL port map( A1 => y_2_port, A2 => 
                           coeff_memory_19_port, Z => mult_28_C95_n764);
   mult_28_C95_U1011 : ADHALFD2 port map( A => mult_28_C95_n563, B => 
                           mult_28_C95_n515, CO => mult_28_C95_n471, S => 
                           mult_28_C95_n472);
   mult_28_C95_U1010 : OAI22DL port map( A1 => mult_28_C95_n697, A2 => 
                           mult_28_C95_n36, B1 => mult_28_C95_n696, B2 => 
                           mult_28_C95_n34, Z => mult_28_C95_n562);
   mult_28_C95_U1009 : EXNOR2D2 port map( A1 => y_11_port, A2 => 
                           coeff_memory_19_port, Z => mult_28_C95_n755);
   mult_28_C95_U1008 : EXNOR2DL port map( A1 => y_8_port, A2 => 
                           coeff_memory_21_port, Z => mult_28_C95_n741);
   mult_28_C95_U1007 : EXNOR2DL port map( A1 => y_8_port, A2 => 
                           coeff_memory_31_port, Z => mult_28_C95_n656);
   mult_28_C95_U1006 : AOI21DL port map( A1 => mult_28_C95_net12285, A2 => 
                           mult_28_C95_n106, B => mult_28_C95_n107, Z => 
                           mult_28_C95_n105);
   mult_28_C95_U1005 : INVDL port map( A => mult_28_C95_n192, Z => 
                           mult_28_C95_net12033);
   mult_28_C95_U1004 : OAI22D2 port map( A1 => mult_28_C95_n657, A2 => 
                           mult_28_C95_n48, B1 => mult_28_C95_n656, B2 => 
                           mult_28_C95_n46, Z => mult_28_C95_n526);
   mult_28_C95_U1003 : INVD2 port map( A => mult_28_C95_n351, Z => 
                           mult_28_C95_n352);
   mult_28_C95_U1002 : EXNOR2DL port map( A1 => y_8_port, A2 => 
                           coeff_memory_27_port, Z => mult_28_C95_n690);
   mult_28_C95_U1001 : INVD1 port map( A => mult_28_C95_net12054, Z => 
                           mult_28_C95_net12055);
   mult_28_C95_U1000 : INVDL port map( A => mult_28_C95_n373, Z => 
                           mult_28_C95_n374);
   mult_28_C95_U999 : EXNOR2D2 port map( A1 => y_13_port, A2 => 
                           coeff_memory_19_port, Z => mult_28_C95_n753);
   mult_28_C95_U998 : EXOR3DL port map( A1 => mult_28_C95_n431, A2 => 
                           mult_28_C95_n420, A3 => mult_28_C95_n912, Z => 
                           mult_28_C95_n943);
   mult_28_C95_U997 : NAN3D2 port map( A1 => mult_28_C95_n940, A2 => 
                           mult_28_C95_n941, A3 => mult_28_C95_n942, Z => 
                           mult_28_C95_n433);
   mult_28_C95_U996 : NAN2D1 port map( A1 => mult_28_C95_n635, A2 => 
                           mult_28_C95_n438, Z => mult_28_C95_n942);
   mult_28_C95_U995 : NAN2D1 port map( A1 => mult_28_C95_n620, A2 => 
                           mult_28_C95_n438, Z => mult_28_C95_n941);
   mult_28_C95_U994 : NAN2D1 port map( A1 => mult_28_C95_n620, A2 => 
                           mult_28_C95_n635, Z => mult_28_C95_n940);
   mult_28_C95_U993 : NAN3D1 port map( A1 => mult_28_C95_n939, A2 => 
                           mult_28_C95_net12078, A3 => mult_28_C95_net12079, Z 
                           => mult_28_C95_n437);
   mult_28_C95_U992 : NAN2DL port map( A1 => mult_28_C95_n575, A2 => 
                           mult_28_C95_n560, Z => mult_28_C95_n939);
   mult_28_C95_U991 : EXOR2D1 port map( A1 => mult_28_C95_n938, A2 => 
                           mult_28_C95_n438, Z => mult_28_C95_n434);
   mult_28_C95_U990 : EXOR2D1 port map( A1 => mult_28_C95_n620, A2 => 
                           mult_28_C95_n635, Z => mult_28_C95_n938);
   mult_28_C95_U989 : INVDL port map( A => mult_28_C95_n171, Z => 
                           mult_28_C95_net12095);
   mult_28_C95_U988 : EXNOR2D2 port map( A1 => y_7_port, A2 => 
                           coeff_memory_23_port, Z => mult_28_C95_n725);
   mult_28_C95_U987 : EXNOR2D2 port map( A1 => y_7_port, A2 => 
                           coeff_memory_27_port, Z => mult_28_C95_n691);
   mult_28_C95_U986 : EXNOR2D1 port map( A1 => coeff_memory_19_port, A2 => 
                           y_9_port, Z => mult_28_C95_n757);
   mult_28_C95_U985 : OAI22D1 port map( A1 => mult_28_C95_n742, A2 => 
                           mult_28_C95_n18, B1 => mult_28_C95_n741, B2 => 
                           mult_28_C95_n16, Z => mult_28_C95_n607);
   mult_28_C95_U984 : ADHALFD2 port map( A => mult_28_C95_n513, B => 
                           mult_28_C95_n530, CO => mult_28_C95_n427, S => 
                           mult_28_C95_n428);
   mult_28_C95_U983 : NAN3D1 port map( A1 => mult_28_C95_n935, A2 => 
                           mult_28_C95_n937, A3 => mult_28_C95_n936, Z => 
                           mult_28_C95_n425);
   mult_28_C95_U982 : NAN2DL port map( A1 => mult_28_C95_n544, A2 => 
                           mult_28_C95_n428, Z => mult_28_C95_n937);
   mult_28_C95_U981 : NAN2DL port map( A1 => mult_28_C95_n559, A2 => 
                           mult_28_C95_n428, Z => mult_28_C95_n936);
   mult_28_C95_U980 : NAN2DL port map( A1 => mult_28_C95_n559, A2 => 
                           mult_28_C95_n544, Z => mult_28_C95_n935);
   mult_28_C95_U979 : EXOR2D1 port map( A1 => mult_28_C95_n544, A2 => 
                           mult_28_C95_n428, Z => mult_28_C95_n934);
   mult_28_C95_U978 : OAI22DL port map( A1 => mult_28_C95_n738, A2 => 
                           mult_28_C95_n18, B1 => mult_28_C95_n737, B2 => 
                           mult_28_C95_n16, Z => mult_28_C95_n603);
   mult_28_C95_U977 : NAN3D1 port map( A1 => mult_28_C95_n933, A2 => 
                           mult_28_C95_net12126, A3 => mult_28_C95_net12125, Z 
                           => mult_28_C95_n407);
   mult_28_C95_U976 : NAN2DL port map( A1 => mult_28_C95_n618, A2 => 
                           mult_28_C95_n603, Z => mult_28_C95_n933);
   mult_28_C95_U975 : INVD1 port map( A => mult_28_C95_net11693, Z => 
                           mult_28_C95_net12151);
   mult_28_C95_U974 : NAN2D2 port map( A1 => mult_28_C95_net12153, A2 => 
                           mult_28_C95_n932, Z => mult_28_C95_n388);
   mult_28_C95_U973 : NAN2D1 port map( A1 => mult_28_C95_net12151, A2 => 
                           mult_28_C95_net12152, Z => mult_28_C95_n932);
   mult_28_C95_U972 : EXNOR2DL port map( A1 => y_2_port, A2 => 
                           coeff_memory_23_port, Z => mult_28_C95_n730);
   mult_28_C95_U971 : OAI22DL port map( A1 => mult_28_C95_n728, A2 => 
                           mult_28_C95_n24, B1 => mult_28_C95_n727, B2 => 
                           mult_28_C95_n22, Z => mult_28_C95_n593);
   mult_28_C95_U970 : EXNOR2D2 port map( A1 => n42, A2 => coeff_memory_23_port,
                           Z => mult_28_C95_n722);
   mult_28_C95_U969 : EXNOR2DL port map( A1 => y_6_port, A2 => 
                           coeff_memory_31_port, Z => mult_28_C95_n658);
   mult_28_C95_U968 : INVDL port map( A => mult_28_C95_net12249, Z => 
                           mult_28_C95_net12250);
   mult_28_C95_U967 : INVDL port map( A => y_9_port, Z => mult_28_C95_net12249)
                           ;
   mult_28_C95_U966 : NAN2DL port map( A1 => mult_28_C95_n606, A2 => 
                           mult_28_C95_n461, Z => mult_28_C95_n967);
   mult_28_C95_U965 : EXOR3D1 port map( A1 => mult_28_C95_n590, A2 => 
                           mult_28_C95_n449, A3 => mult_28_C95_n605, Z => 
                           mult_28_C95_n436);
   mult_28_C95_U964 : OAI22D1 port map( A1 => mult_28_C95_n656, A2 => 
                           mult_28_C95_n48, B1 => mult_28_C95_n655, B2 => 
                           mult_28_C95_n46, Z => mult_28_C95_n333);
   mult_28_C95_U963 : INVDL port map( A => mult_28_C95_n915, Z => 
                           mult_28_C95_net12257);
   mult_28_C95_U962 : EXNOR2DL port map( A1 => y_6_port, A2 => 
                           coeff_memory_17_port, Z => mult_28_C95_n777);
   mult_28_C95_U961 : EXNOR2D2 port map( A1 => mult_28_C95_net12250, A2 => 
                           coeff_memory_29_port, Z => mult_28_C95_n672);
   mult_28_C95_U960 : EXNOR2D2 port map( A1 => y_11_port, A2 => 
                           coeff_memory_25_port, Z => mult_28_C95_n704);
   mult_28_C95_U959 : EXNOR2D1 port map( A1 => coeff_memory_23_port, A2 => 
                           coeff_memory_24_port, Z => mult_28_C95_n28);
   mult_28_C95_U958 : NAN2D1 port map( A1 => mult_28_C95_n804, A2 => 
                           mult_28_C95_n28, Z => mult_28_C95_n30);
   mult_28_C95_U957 : OAI21D1 port map( A1 => mult_28_C95_n211, A2 => 
                           mult_28_C95_n209, B => mult_28_C95_n931, Z => 
                           mult_28_C95_n208);
   mult_28_C95_U956 : BUFDL port map( A => mult_28_C95_n210, Z => 
                           mult_28_C95_n931);
   mult_28_C95_U955 : INVD1 port map( A => mult_28_C95_n212, Z => 
                           mult_28_C95_n211);
   mult_28_C95_U954 : AND2D1 port map( A1 => mult_28_C95_n285, A2 => 
                           mult_28_C95_n180, Z => mult_28_C95_net11172);
   mult_28_C95_U953 : INVDL port map( A => mult_28_C95_n187, Z => 
                           mult_28_C95_net11745);
   mult_28_C95_U952 : INVDL port map( A => mult_28_C95_n901, Z => 
                           mult_28_C95_n192);
   mult_28_C95_U951 : NOR2D1 port map( A1 => mult_28_C95_n206, A2 => 
                           mult_28_C95_n209, Z => mult_28_C95_n204);
   mult_28_C95_U950 : OAI21D1 port map( A1 => mult_28_C95_n206, A2 => 
                           mult_28_C95_n210, B => mult_28_C95_n207, Z => 
                           mult_28_C95_n205);
   mult_28_C95_U949 : EXOR2D1 port map( A1 => mult_28_C95_net11829, A2 => 
                           mult_28_C95_n571, Z => mult_28_C95_n384);
   mult_28_C95_U948 : AOI21M10DL port map( A1 => mult_28_C95_n900, A2 => 
                           mult_28_C95_n51, B => mult_28_C95_n171, Z => 
                           mult_28_C95_n169);
   mult_28_C95_U947 : NAN2D1 port map( A1 => mult_28_C95_n161, A2 => 
                           mult_28_C95_n132, Z => mult_28_C95_n53);
   mult_28_C95_U946 : NAN3D1 port map( A1 => mult_28_C95_net11585, A2 => 
                           mult_28_C95_net11587, A3 => mult_28_C95_net11586, Z 
                           => mult_28_C95_n387);
   mult_28_C95_U945 : EXNOR2D1 port map( A1 => coeff_memory_27_port, A2 => 
                           coeff_memory_28_port, Z => mult_28_C95_n40);
   mult_28_C95_U944 : NAN2D1 port map( A1 => mult_28_C95_n802, A2 => 
                           mult_28_C95_n40, Z => mult_28_C95_n42);
   mult_28_C95_U943 : EXNOR2D2 port map( A1 => y_3_port, A2 => 
                           coeff_memory_29_port, Z => mult_28_C95_n678);
   mult_28_C95_U942 : EXNOR2D1 port map( A1 => coeff_memory_25_port, A2 => 
                           coeff_memory_26_port, Z => mult_28_C95_n34);
   mult_28_C95_U941 : EXNOR2D2 port map( A1 => y_6_port, A2 => 
                           coeff_memory_27_port, Z => mult_28_C95_n692);
   mult_28_C95_U940 : NAN2D1 port map( A1 => mult_28_C95_n803, A2 => 
                           mult_28_C95_n34, Z => mult_28_C95_n36);
   mult_28_C95_U939 : NAN2DL port map( A1 => mult_28_C95_n588, A2 => 
                           mult_28_C95_n425, Z => mult_28_C95_n928);
   mult_28_C95_U938 : NAN2DL port map( A1 => mult_28_C95_n425, A2 => 
                           mult_28_C95_n573, Z => mult_28_C95_n930);
   mult_28_C95_U937 : NAN2DL port map( A1 => mult_28_C95_n588, A2 => 
                           mult_28_C95_n573, Z => mult_28_C95_n929);
   mult_28_C95_U936 : NAN3D1 port map( A1 => mult_28_C95_n928, A2 => 
                           mult_28_C95_n930, A3 => mult_28_C95_n929, Z => 
                           mult_28_C95_n409);
   mult_28_C95_U935 : EXNOR2D1 port map( A1 => y_8_port, A2 => 
                           coeff_memory_25_port, Z => mult_28_C95_n707);
   mult_28_C95_U934 : EXOR3D2 port map( A1 => mult_28_C95_n412, A2 => 
                           mult_28_C95_n618, A3 => mult_28_C95_n603, Z => 
                           mult_28_C95_n408);
   mult_28_C95_U933 : NAN2DL port map( A1 => mult_28_C95_n618, A2 => 
                           mult_28_C95_n412, Z => mult_28_C95_net12125);
   mult_28_C95_U932 : NAN2DL port map( A1 => mult_28_C95_n603, A2 => 
                           mult_28_C95_n412, Z => mult_28_C95_net12126);
   mult_28_C95_U931 : NAN2D1 port map( A1 => mult_28_C95_n395, A2 => 
                           mult_28_C95_n616, Z => mult_28_C95_net11666);
   mult_28_C95_U930 : NAN2DL port map( A1 => mult_28_C95_n395, A2 => 
                           mult_28_C95_n393, Z => mult_28_C95_net11667);
   mult_28_C95_U929 : EXOR3D1 port map( A1 => mult_28_C95_n395, A2 => 
                           mult_28_C95_n616, A3 => mult_28_C95_n393, Z => 
                           mult_28_C95_n380);
   mult_28_C95_U928 : NAN2DL port map( A1 => mult_28_C95_n403, A2 => 
                           mult_28_C95_n392, Z => mult_28_C95_net11587);
   mult_28_C95_U927 : EXNOR2D1 port map( A1 => mult_28_C95_n392, A2 => 
                           mult_28_C95_n403, Z => mult_28_C95_net11693);
   mult_28_C95_U926 : EXOR3D2 port map( A1 => mult_28_C95_n575, A2 => 
                           mult_28_C95_n560, A3 => mult_28_C95_n440, Z => 
                           mult_28_C95_n438);
   mult_28_C95_U925 : NAN2DL port map( A1 => mult_28_C95_n575, A2 => 
                           mult_28_C95_n440, Z => mult_28_C95_net12078);
   mult_28_C95_U924 : NAN2DL port map( A1 => mult_28_C95_n560, A2 => 
                           mult_28_C95_n440, Z => mult_28_C95_net12079);
   mult_28_C95_U923 : AO21D2 port map( A1 => mult_28_C95_n6, A2 => 
                           mult_28_C95_n824, B => mult_28_C95_n768, Z => 
                           mult_28_C95_n633);
   mult_28_C95_U922 : NAN2DL port map( A1 => mult_28_C95_n604, A2 => 
                           mult_28_C95_n426, Z => mult_28_C95_n925);
   mult_28_C95_U921 : NAN2D1 port map( A1 => mult_28_C95_n634, A2 => 
                           mult_28_C95_n426, Z => mult_28_C95_n927);
   mult_28_C95_U920 : INVD1 port map( A => coeff_memory_16_port, Z => 
                           mult_28_C95_n824);
   mult_28_C95_U919 : NAN2D1 port map( A1 => mult_28_C95_n634, A2 => 
                           mult_28_C95_n905, Z => mult_28_C95_n926);
   mult_28_C95_U918 : NAN3D2 port map( A1 => mult_28_C95_n925, A2 => 
                           mult_28_C95_n927, A3 => mult_28_C95_n926, Z => 
                           mult_28_C95_n421);
   mult_28_C95_U917 : EXOR2D2 port map( A1 => mult_28_C95_n417, A2 => 
                           mult_28_C95_n406, Z => mult_28_C95_net11503);
   mult_28_C95_U916 : NAN2DL port map( A1 => mult_28_C95_n417, A2 => 
                           mult_28_C95_n406, Z => mult_28_C95_net11507);
   mult_28_C95_U915 : NAN2DL port map( A1 => mult_28_C95_n406, A2 => 
                           mult_28_C95_n404, Z => mult_28_C95_net11509);
   mult_28_C95_U914 : NAN2D1 port map( A1 => mult_28_C95_n390, A2 => 
                           mult_28_C95_n392, Z => mult_28_C95_net11586);
   mult_28_C95_U913 : NAN2DL port map( A1 => mult_28_C95_n390, A2 => 
                           mult_28_C95_n403, Z => mult_28_C95_net11585);
   mult_28_C95_U912 : NAN2D1 port map( A1 => mult_28_C95_net11693, A2 => 
                           mult_28_C95_n390, Z => mult_28_C95_net12153);
   mult_28_C95_U911 : INVDL port map( A => mult_28_C95_n390, Z => 
                           mult_28_C95_net12152);
   mult_28_C95_U910 : ADFULD2 port map( A => mult_28_C95_n394, B => 
                           mult_28_C95_n407, CI => mult_28_C95_n405, CO => 
                           mult_28_C95_n389, S => mult_28_C95_n390);
   mult_28_C95_U909 : EXOR3DL port map( A1 => mult_28_C95_n389, A2 => 
                           mult_28_C95_n380, A3 => mult_28_C95_n902, Z => 
                           mult_28_C95_net12019);
   mult_28_C95_U908 : NAN2D1 port map( A1 => mult_28_C95_net12019, A2 => 
                           mult_28_C95_n387, Z => mult_28_C95_n187);
   mult_28_C95_U907 : NAN2D1 port map( A1 => mult_28_C95_n375, A2 => 
                           mult_28_C95_n364, Z => mult_28_C95_n180);
   mult_28_C95_U906 : NOR2D1 port map( A1 => mult_28_C95_n172, A2 => 
                           mult_28_C95_n167, Z => mult_28_C95_n161);
   mult_28_C95_U905 : AOI21DL port map( A1 => mult_28_C95_n132, A2 => 
                           mult_28_C95_n162, B => mult_28_C95_n903, Z => 
                           mult_28_C95_n52);
   mult_28_C95_U904 : AOI21DL port map( A1 => mult_28_C95_n132, A2 => 
                           mult_28_C95_n162, B => mult_28_C95_n903, Z => 
                           mult_28_C95_net12183);
   mult_28_C95_U903 : AND2DL port map( A1 => mult_28_C95_n282, A2 => 
                           mult_28_C95_n155, Z => mult_28_C95_net11662);
   mult_28_C95_U902 : NAN2D1 port map( A1 => mult_28_C95_n336, A2 => 
                           mult_28_C95_n343, Z => mult_28_C95_n155);
   mult_28_C95_U901 : NOR2D1 port map( A1 => mult_28_C95_n134, A2 => 
                           mult_28_C95_n154, Z => mult_28_C95_n132);
   mult_28_C95_U900 : INVD1 port map( A => mult_28_C95_n154, Z => 
                           mult_28_C95_n282);
   mult_28_C95_U899 : NOR2D1 port map( A1 => mult_28_C95_n336, A2 => 
                           mult_28_C95_n343, Z => mult_28_C95_n154);
   mult_28_C95_U898 : INVD1 port map( A => mult_28_C95_n150, Z => 
                           mult_28_C95_n148);
   mult_28_C95_U897 : NAN2DL port map( A1 => mult_28_C95_n328, A2 => 
                           mult_28_C95_n335, Z => mult_28_C95_n150);
   mult_28_C95_U896 : AOI21M10DL port map( A1 => mult_28_C95_n155, A2 => 
                           mult_28_C95_net11096, B => mult_28_C95_n148, Z => 
                           mult_28_C95_n144);
   mult_28_C95_U895 : NAN2D1 port map( A1 => mult_28_C95_net11096, A2 => 
                           mult_28_C95_net11083, Z => mult_28_C95_n134);
   mult_28_C95_U894 : NAN2DL port map( A1 => mult_28_C95_n282, A2 => 
                           mult_28_C95_net11096, Z => mult_28_C95_n143);
   mult_28_C95_U893 : OR2D1 port map( A1 => mult_28_C95_n328, A2 => 
                           mult_28_C95_n335, Z => mult_28_C95_net11096);
   mult_28_C95_U892 : INVBD2 port map( A => mult_28_C95_net10037, Z => 
                           mult_28_C95_net12285);
   mult_28_C95_U891 : INVD2 port map( A => mult_28_C95_n51, Z => 
                           mult_28_C95_net10037);
   mult_28_C95_U890 : EXNOR2DL port map( A1 => mult_28_C95_net11621, A2 => 
                           mult_28_C95_n63, Z => m3_6);
   mult_28_C95_U889 : NOR2DL port map( A1 => mult_28_C95_n163, A2 => 
                           mult_28_C95_n143, Z => mult_28_C95_n141);
   mult_28_C95_U888 : INVDL port map( A => mult_28_C95_n161, Z => 
                           mult_28_C95_n163);
   mult_28_C95_U887 : AND2DL port map( A1 => mult_28_C95_net11096, A2 => 
                           mult_28_C95_n150, Z => mult_28_C95_net11675);
   mult_28_C95_U886 : EXNOR2D2 port map( A1 => mult_28_C95_n151, A2 => 
                           mult_28_C95_net11675, Z => m3_9);
   mult_28_C95_U885 : INVDL port map( A => mult_28_C95_n200, Z => 
                           mult_28_C95_n288);
   mult_28_C95_U884 : OAI21D1 port map( A1 => mult_28_C95_n195, A2 => 
                           mult_28_C95_n201, B => mult_28_C95_n196, Z => 
                           mult_28_C95_net12065);
   mult_28_C95_U883 : INVDL port map( A => mult_28_C95_n195, Z => 
                           mult_28_C95_n287);
   mult_28_C95_U882 : OAI21D1 port map( A1 => mult_28_C95_n187, A2 => 
                           mult_28_C95_n179, B => mult_28_C95_n180, Z => 
                           mult_28_C95_n178);
   mult_28_C95_U881 : INVDL port map( A => mult_28_C95_n184, Z => 
                           mult_28_C95_net12054);
   mult_28_C95_U880 : NOR2M1DL port map( A1 => mult_28_C95_n189, A2 => 
                           mult_28_C95_net12055, Z => mult_28_C95_n182);
   mult_28_C95_U879 : BUFDL port map( A => mult_28_C95_n189, Z => 
                           mult_28_C95_net12127);
   mult_28_C95_U878 : NOR2D1 port map( A1 => mult_28_C95_n195, A2 => 
                           mult_28_C95_n200, Z => mult_28_C95_n189);
   mult_28_C95_U877 : NOR2D2 port map( A1 => mult_28_C95_n184, A2 => 
                           mult_28_C95_n179, Z => mult_28_C95_n177);
   mult_28_C95_U876 : OAI21D1 port map( A1 => mult_28_C95_n175, A2 => 
                           mult_28_C95_n203, B => mult_28_C95_n176, Z => 
                           mult_28_C95_n51);
   mult_28_C95_U875 : NAN2D1 port map( A1 => mult_28_C95_n177, A2 => 
                           mult_28_C95_n189, Z => mult_28_C95_n175);
   mult_28_C95_U874 : EXNOR2D2 port map( A1 => n38, A2 => coeff_memory_27_port,
                           Z => mult_28_C95_n693);
   mult_28_C95_U873 : EXOR3D1 port map( A1 => mult_28_C95_n389, A2 => 
                           mult_28_C95_n380, A3 => mult_28_C95_n902, Z => 
                           mult_28_C95_n376);
   mult_28_C95_U872 : INVDL port map( A => mult_28_C95_n173, Z => 
                           mult_28_C95_n924);
   mult_28_C95_U871 : OA21M20D1 port map( A1 => mult_28_C95_n283, A2 => 
                           mult_28_C95_n924, B => mult_28_C95_n168, Z => 
                           mult_28_C95_n164);
   mult_28_C95_U870 : INVDL port map( A => mult_28_C95_n473, Z => 
                           mult_28_C95_n923);
   mult_28_C95_U869 : AOI21M20DL port map( A1 => mult_28_C95_n336, A2 => 
                           mult_28_C95_n343, B => mult_28_C95_n163, Z => 
                           mult_28_C95_n152);
   mult_28_C95_U868 : NAN2D1 port map( A1 => mult_28_C95_n605, A2 => 
                           mult_28_C95_n590, Z => mult_28_C95_n985);
   mult_28_C95_U867 : NAN2M1D1 port map( A1 => mult_28_C95_n209, A2 => 
                           mult_28_C95_n931, Z => mult_28_C95_n69);
   mult_28_C95_U866 : EXNOR2D2 port map( A1 => n36, A2 => coeff_memory_25_port,
                           Z => mult_28_C95_n714);
   mult_28_C95_U865 : ADHALFD1 port map( A => mult_28_C95_n580, B => 
                           mult_28_C95_n516, CO => mult_28_C95_n487, S => 
                           mult_28_C95_n488);
   mult_28_C95_U864 : NAN2D1 port map( A1 => mult_28_C95_n990, A2 => 
                           mult_28_C95_n993, Z => mult_28_C95_n213);
   mult_28_C95_U863 : AOI21DL port map( A1 => mult_28_C95_n288, A2 => 
                           mult_28_C95_n202, B => mult_28_C95_n199, Z => 
                           mult_28_C95_n197);
   mult_28_C95_U862 : INVBD2 port map( A => mult_28_C95_net10037, Z => 
                           mult_28_C95_net11621);
   mult_28_C95_U861 : INVD2 port map( A => n36, Z => mult_28_C95_n919);
   mult_28_C95_U860 : NAN2D2 port map( A1 => mult_28_C95_n921, A2 => 
                           mult_28_C95_n922, Z => mult_28_C95_n663);
   mult_28_C95_U859 : NAN2D2 port map( A1 => mult_28_C95_n919, A2 => 
                           mult_28_C95_n920, Z => mult_28_C95_n922);
   mult_28_C95_U858 : NAN2D1 port map( A1 => n36, A2 => coeff_memory_31_port, Z
                           => mult_28_C95_n921);
   mult_28_C95_U857 : INVDL port map( A => mult_28_C95_n368, Z => 
                           mult_28_C95_n916);
   mult_28_C95_U856 : NAN2D1 port map( A1 => mult_28_C95_n917, A2 => 
                           mult_28_C95_n918, Z => mult_28_C95_net11025);
   mult_28_C95_U855 : NAN2D1 port map( A1 => mult_28_C95_n915, A2 => 
                           mult_28_C95_n916, Z => mult_28_C95_n918);
   mult_28_C95_U854 : NAN2DL port map( A1 => mult_28_C95_n377, A2 => 
                           mult_28_C95_n368, Z => mult_28_C95_n917);
   mult_28_C95_U853 : ADFULD2 port map( A => mult_28_C95_n574, B => 
                           mult_28_C95_n439, CI => mult_28_C95_n589, CO => 
                           mult_28_C95_n423, S => mult_28_C95_n424);
   mult_28_C95_U852 : ADFULD2 port map( A => mult_28_C95_n380, B => 
                           mult_28_C95_n389, CI => mult_28_C95_n378, CO => 
                           mult_28_C95_n375, S => mult_28_C95_n_1033);
   mult_28_C95_U851 : EXNOR2DL port map( A1 => y_2_port, A2 => 
                           coeff_memory_21_port, Z => mult_28_C95_n747);
   mult_28_C95_U850 : EXNOR2D2 port map( A1 => mult_28_C95_n169, A2 => 
                           mult_28_C95_n989, Z => m3_7);
   mult_28_C95_U849 : EXNOR2D2 port map( A1 => mult_28_C95_n208, A2 => 
                           mult_28_C95_n68, Z => m3_1);
   mult_28_C95_U848 : EXNOR2DL port map( A1 => y_6_port, A2 => 
                           coeff_memory_19_port, Z => mult_28_C95_n760);
   mult_28_C95_U847 : BUFDL port map( A => y_11_port, Z => mult_28_C95_n914);
   mult_28_C95_U846 : OAI22D1 port map( A1 => mult_28_C95_n769, A2 => 
                           mult_28_C95_n6, B1 => mult_28_C95_n768, B2 => 
                           mult_28_C95_n824, Z => mult_28_C95_n634);
   mult_28_C95_U845 : EXNOR2DL port map( A1 => y_2_port, A2 => 
                           coeff_memory_17_port, Z => mult_28_C95_n781);
   mult_28_C95_U844 : EXOR3D2 port map( A1 => mult_28_C95_n979, A2 => 
                           mult_28_C95_n905, A3 => mult_28_C95_n426, Z => 
                           mult_28_C95_n422);
   mult_28_C95_U843 : NAN2D1 port map( A1 => mult_28_C95_n605, A2 => 
                           mult_28_C95_n449, Z => mult_28_C95_n984);
   mult_28_C95_U842 : NAN3D1 port map( A1 => mult_28_C95_net11666, A2 => 
                           mult_28_C95_net11667, A3 => mult_28_C95_n972, Z => 
                           mult_28_C95_n379);
   mult_28_C95_U841 : NOR2DL port map( A1 => mult_28_C95_n364, A2 => 
                           mult_28_C95_n375, Z => mult_28_C95_n913);
   mult_28_C95_U840 : AOI22M10D1 port map( B1 => mult_28_C95_n995, B2 => 
                           mult_28_C95_n230, A1 => mult_28_C95_n923, A2 => 
                           mult_28_C95_n464, Z => mult_28_C95_n225);
   mult_28_C95_U839 : EXNOR2DL port map( A1 => y_3_port, A2 => 
                           coeff_memory_17_port, Z => mult_28_C95_n780);
   mult_28_C95_U838 : EXNOR2D2 port map( A1 => n42, A2 => coeff_memory_19_port,
                           Z => mult_28_C95_n756);
   mult_28_C95_U837 : OR2D2 port map( A1 => mult_28_C95_n474, A2 => 
                           mult_28_C95_n481, Z => mult_28_C95_n991);
   mult_28_C95_U836 : NAN2M1D1 port map( A1 => mult_28_C95_n206, A2 => 
                           mult_28_C95_n207, Z => mult_28_C95_n68);
   mult_28_C95_U835 : EXOR3DL port map( A1 => mult_28_C95_n424, A2 => 
                           mult_28_C95_n433, A3 => mult_28_C95_n422, Z => 
                           mult_28_C95_n912);
   mult_28_C95_U834 : EXOR2D2 port map( A1 => mult_28_C95_n455, A2 => 
                           mult_28_C95_n446, Z => mult_28_C95_n958);
   mult_28_C95_U833 : AND2DL port map( A1 => mult_28_C95_n474, A2 => 
                           mult_28_C95_n481, Z => mult_28_C95_n911);
   mult_28_C95_U832 : AOI21D1 port map( A1 => mult_28_C95_n991, A2 => 
                           mult_28_C95_n999, B => mult_28_C95_n911, Z => 
                           mult_28_C95_n232);
   mult_28_C95_U831 : OR2DL port map( A1 => mult_28_C95_n482, A2 => 
                           mult_28_C95_n489, Z => mult_28_C95_n998);
   mult_28_C95_U830 : EXNOR2D1 port map( A1 => y_11_port, A2 => 
                           coeff_memory_23_port, Z => mult_28_C95_n721);
   mult_28_C95_U829 : AND2DL port map( A1 => mult_28_C95_n287, A2 => 
                           mult_28_C95_n196, Z => mult_28_C95_n910);
   mult_28_C95_U828 : EXNOR2D2 port map( A1 => mult_28_C95_n197, A2 => 
                           mult_28_C95_n910, Z => m3_3);
   mult_28_C95_U827 : INVD1 port map( A => coeff_memory_31_port, Z => 
                           mult_28_C95_n920);
   mult_28_C95_U826 : INVD1 port map( A => mult_28_C95_n377, Z => 
                           mult_28_C95_n915);
   mult_28_C95_U825 : INVD1 port map( A => mult_28_C95_n56, Z => 
                           mult_28_C95_n947);
   mult_28_C95_U824 : EXOR2D1 port map( A1 => mult_28_C95_n934, A2 => 
                           mult_28_C95_n559, Z => mult_28_C95_n426);
   mult_28_C95_U823 : OAI22DL port map( A1 => mult_28_C95_n741, A2 => 
                           mult_28_C95_n18, B1 => mult_28_C95_n740, B2 => 
                           mult_28_C95_n16, Z => mult_28_C95_n606);
   mult_28_C95_U822 : OAI22DL port map( A1 => mult_28_C95_n688, A2 => 
                           mult_28_C95_n36, B1 => mult_28_C95_n687, B2 => 
                           mult_28_C95_n34, Z => mult_28_C95_n553);
   mult_28_C95_U821 : OAI22D2 port map( A1 => mult_28_C95_n752, A2 => 
                           mult_28_C95_n12, B1 => mult_28_C95_n751, B2 => 
                           mult_28_C95_n9, Z => mult_28_C95_n617);
   mult_28_C95_U820 : NAN2DL port map( A1 => mult_28_C95_n409, A2 => 
                           mult_28_C95_n617, Z => mult_28_C95_n909);
   mult_28_C95_U819 : NAN2D1 port map( A1 => mult_28_C95_n396, A2 => 
                           mult_28_C95_n617, Z => mult_28_C95_n908);
   mult_28_C95_U818 : NAN2D1 port map( A1 => mult_28_C95_n396, A2 => 
                           mult_28_C95_n409, Z => mult_28_C95_n907);
   mult_28_C95_U817 : EXOR2D1 port map( A1 => mult_28_C95_n906, A2 => 
                           mult_28_C95_n396, Z => mult_28_C95_n392);
   mult_28_C95_U816 : EXOR2D1 port map( A1 => mult_28_C95_n617, A2 => 
                           mult_28_C95_n409, Z => mult_28_C95_n906);
   mult_28_C95_U815 : OAI22D4 port map( A1 => mult_28_C95_n662, A2 => 
                           mult_28_C95_n48, B1 => mult_28_C95_n661, B2 => 
                           mult_28_C95_n46, Z => mult_28_C95_n399);
   mult_28_C95_U814 : INVD4 port map( A => mult_28_C95_n399, Z => 
                           mult_28_C95_n400);
   mult_28_C95_U813 : EXNOR2D1 port map( A1 => y_12_port, A2 => 
                           coeff_memory_21_port, Z => mult_28_C95_n737);
   mult_28_C95_U812 : NAN2D2 port map( A1 => mult_28_C95_n354, A2 => 
                           mult_28_C95_n363, Z => mult_28_C95_n173);
   mult_28_C95_U811 : EXNOR2D2 port map( A1 => y_11_port, A2 => 
                           coeff_memory_21_port, Z => mult_28_C95_n738);
   mult_28_C95_U810 : OAI22DL port map( A1 => mult_28_C95_n739, A2 => 
                           mult_28_C95_n18, B1 => mult_28_C95_n738, B2 => 
                           mult_28_C95_n16, Z => mult_28_C95_n604);
   mult_28_C95_U809 : OAI22D1 port map( A1 => mult_28_C95_n739, A2 => 
                           mult_28_C95_n18, B1 => mult_28_C95_n738, B2 => 
                           mult_28_C95_n16, Z => mult_28_C95_n905);
   mult_28_C95_U808 : EXNOR2DL port map( A1 => y_4_port, A2 => 
                           coeff_memory_19_port, Z => mult_28_C95_n762);
   mult_28_C95_U807 : EXNOR2DL port map( A1 => y_4_port, A2 => 
                           coeff_memory_17_port, Z => mult_28_C95_n779);
   mult_28_C95_U806 : EXNOR2DL port map( A1 => y_4_port, A2 => 
                           coeff_memory_31_port, Z => mult_28_C95_n660);
   mult_28_C95_U805 : EXNOR2D2 port map( A1 => y_7_port, A2 => 
                           coeff_memory_25_port, Z => mult_28_C95_n708);
   mult_28_C95_U804 : EXNOR2D1 port map( A1 => y_15_port, A2 => 
                           coeff_memory_21_port, Z => mult_28_C95_n734);
   mult_28_C95_U803 : OAI22D1 port map( A1 => mult_28_C95_n726, A2 => 
                           mult_28_C95_n24, B1 => mult_28_C95_n725, B2 => 
                           mult_28_C95_n22, Z => mult_28_C95_n591);
   mult_28_C95_U802 : OAI22D1 port map( A1 => mult_28_C95_n16, A2 => 
                           mult_28_C95_n734, B1 => mult_28_C95_n18, B2 => 
                           mult_28_C95_n735, Z => mult_28_C95_n600);
   mult_28_C95_U801 : EXNOR2D2 port map( A1 => y_8_port, A2 => 
                           coeff_memory_23_port, Z => mult_28_C95_n724);
   mult_28_C95_U800 : EXNOR2D2 port map( A1 => n36, A2 => coeff_memory_27_port,
                           Z => mult_28_C95_n697);
   mult_28_C95_U799 : NAN3D2 port map( A1 => mult_28_C95_n907, A2 => 
                           mult_28_C95_n909, A3 => mult_28_C95_n908, Z => 
                           mult_28_C95_n391);
   mult_28_C95_U798 : EXNOR2D2 port map( A1 => y_7_port, A2 => 
                           coeff_memory_29_port, Z => mult_28_C95_n674);
   mult_28_C95_U797 : INVDL port map( A => mult_28_C95_n203, Z => 
                           mult_28_C95_n202);
   mult_28_C95_U796 : EXNOR2D2 port map( A1 => y_9_port, A2 => 
                           coeff_memory_31_port, Z => mult_28_C95_n655);
   mult_28_C95_U795 : OAI21DL port map( A1 => mult_28_C95_n164, A2 => 
                           mult_28_C95_n154, B => mult_28_C95_n155, Z => 
                           mult_28_C95_n153);
   mult_28_C95_U794 : BUFDL port map( A => mult_28_C95_n162, Z => 
                           mult_28_C95_n904);
   mult_28_C95_U793 : OA21M20DL port map( A1 => mult_28_C95_net11083, A2 => 
                           mult_28_C95_n148, B => mult_28_C95_n139, Z => 
                           mult_28_C95_n135);
   mult_28_C95_U792 : OAI21DL port map( A1 => mult_28_C95_n134, A2 => 
                           mult_28_C95_n155, B => mult_28_C95_n135, Z => 
                           mult_28_C95_n903);
   mult_28_C95_U791 : EXNOR2D2 port map( A1 => y_9_port, A2 => 
                           coeff_memory_25_port, Z => mult_28_C95_n706);
   mult_28_C95_U790 : EXNOR2D2 port map( A1 => y_6_port, A2 => 
                           coeff_memory_23_port, Z => mult_28_C95_n726);
   mult_28_C95_U789 : EXOR3D1 port map( A1 => mult_28_C95_n382, A2 => 
                           mult_28_C95_n384, A3 => mult_28_C95_n391, Z => 
                           mult_28_C95_n902);
   mult_28_C95_U788 : OAI21DL port map( A1 => mult_28_C95_n195, A2 => 
                           mult_28_C95_n201, B => mult_28_C95_n196, Z => 
                           mult_28_C95_n901);
   mult_28_C95_U787 : INVDL port map( A => mult_28_C95_n284, Z => 
                           mult_28_C95_n900);
   mult_28_C95_U786 : EXOR2D2 port map( A1 => mult_28_C95_n973, A2 => 
                           mult_28_C95_n379, Z => mult_28_C95_n366);
   mult_28_C95_U785 : AOI21M10D1 port map( A1 => mult_28_C95_n163, A2 => 
                           mult_28_C95_net11621, B => mult_28_C95_n904, Z => 
                           mult_28_C95_n160);
   mult_28_C95_U784 : EXNOR2D1 port map( A1 => n42, A2 => coeff_memory_29_port,
                           Z => mult_28_C95_n671);
   mult_28_C95_U783 : OR2DL port map( A1 => mult_28_C95_n647, A2 => 
                           mult_28_C95_n632, Z => mult_28_C95_n1006);
   mult_28_C95_U782 : ADFULDL port map( A => mult_28_C95_n511, B => 
                           mult_28_C95_n615, CI => mult_28_C95_n630, CO => 
                           mult_28_C95_n509, S => mult_28_C95_n510);
   mult_28_C95_U781 : OR2D1 port map( A1 => mult_28_C95_n529, A2 => 
                           mult_28_C95_n427, Z => mult_28_C95_n413);
   mult_28_C95_U780 : EXNOR2D1 port map( A1 => mult_28_C95_n529, A2 => 
                           mult_28_C95_n427, Z => mult_28_C95_n414);
   mult_28_C95_U779 : OAI22DL port map( A1 => mult_28_C95_n781, A2 => 
                           mult_28_C95_n6, B1 => mult_28_C95_n780, B2 => 
                           mult_28_C95_n824, Z => mult_28_C95_n646);
   mult_28_C95_U778 : OAI22DL port map( A1 => mult_28_C95_n747, A2 => 
                           mult_28_C95_n18, B1 => mult_28_C95_n746, B2 => 
                           mult_28_C95_n16, Z => mult_28_C95_n612);
   mult_28_C95_U777 : OAI22DL port map( A1 => mult_28_C95_n748, A2 => 
                           mult_28_C95_n18, B1 => mult_28_C95_n747, B2 => 
                           mult_28_C95_n16, Z => mult_28_C95_n613);
   mult_28_C95_U776 : OAI22DL port map( A1 => mult_28_C95_n730, A2 => 
                           mult_28_C95_n24, B1 => mult_28_C95_n729, B2 => 
                           mult_28_C95_n22, Z => mult_28_C95_n595);
   mult_28_C95_U775 : OAI22DL port map( A1 => mult_28_C95_n731, A2 => 
                           mult_28_C95_n24, B1 => mult_28_C95_n730, B2 => 
                           mult_28_C95_n22, Z => mult_28_C95_n596);
   mult_28_C95_U774 : OAI22DL port map( A1 => mult_28_C95_n764, A2 => 
                           mult_28_C95_n12, B1 => mult_28_C95_n763, B2 => 
                           mult_28_C95_n9, Z => mult_28_C95_n629);
   mult_28_C95_U773 : OAI22DL port map( A1 => mult_28_C95_n765, A2 => 
                           mult_28_C95_n12, B1 => mult_28_C95_n764, B2 => 
                           mult_28_C95_n9, Z => mult_28_C95_n630);
   mult_28_C95_U772 : OAI22DL port map( A1 => mult_28_C95_n663, A2 => 
                           mult_28_C95_n48, B1 => mult_28_C95_n662, B2 => 
                           mult_28_C95_n46, Z => mult_28_C95_n529);
   mult_28_C95_U771 : OAI22DL port map( A1 => mult_28_C95_n713, A2 => 
                           mult_28_C95_n30, B1 => mult_28_C95_n712, B2 => 
                           mult_28_C95_n28, Z => mult_28_C95_n578);
   mult_28_C95_U770 : OAI22DL port map( A1 => mult_28_C95_n714, A2 => 
                           mult_28_C95_n30, B1 => mult_28_C95_n713, B2 => 
                           mult_28_C95_n28, Z => mult_28_C95_n579);
   mult_28_C95_U769 : EXNOR2D2 port map( A1 => n36, A2 => coeff_memory_29_port,
                           Z => mult_28_C95_n680);
   mult_28_C95_U768 : OAI22D1 port map( A1 => mult_28_C95_n680, A2 => 
                           mult_28_C95_n42, B1 => mult_28_C95_n679, B2 => 
                           mult_28_C95_n40, Z => mult_28_C95_n545);
   mult_28_C95_U767 : EXOR2D1 port map( A1 => mult_28_C95_net11503, A2 => 
                           mult_28_C95_n404, Z => mult_28_C95_n402);
   mult_28_C95_U551 : OAI22D1 port map( A1 => mult_28_C95_n707, A2 => 
                           mult_28_C95_n30, B1 => mult_28_C95_n706, B2 => 
                           mult_28_C95_n28, Z => mult_28_C95_n572);
   mult_28_C95_U178 : AOI21D1 port map( A1 => mult_28_C95_n177, A2 => 
                           mult_28_C95_net12065, B => mult_28_C95_n178, Z => 
                           mult_28_C95_n176);
   mult_28_C95_U144 : AOI21D1 port map( A1 => mult_28_C95_net11621, A2 => 
                           mult_28_C95_n152, B => mult_28_C95_n153, Z => 
                           mult_28_C95_n151);
   mult_28_C95_U132 : OAI21D1 port map( A1 => mult_28_C95_n164, A2 => 
                           mult_28_C95_n143, B => mult_28_C95_n144, Z => 
                           mult_28_C95_n142);
   mult_28_C95_U162 : OAI21D1 port map( A1 => mult_28_C95_n167, A2 => 
                           mult_28_C95_n173, B => mult_28_C95_n168, Z => 
                           mult_28_C95_n162);
   mult_28_C95_U193 : NOR2D2 port map( A1 => mult_28_C95_n376, A2 => 
                           mult_28_C95_n387, Z => mult_28_C95_n184);
   mult_28_C95_U183 : NOR2D2 port map( A1 => mult_28_C95_n364, A2 => 
                           mult_28_C95_n375, Z => mult_28_C95_n179);
   mult_28_C95_U384 : ADFULD1 port map( A => mult_28_C95_n423, B => 
                           mult_28_C95_n633, CI => mult_28_C95_n421, CO => 
                           mult_28_C95_n405, S => mult_28_C95_n406);
   mult_28_C95_U391 : ADFULD1 port map( A => mult_28_C95_n433, B => 
                           mult_28_C95_n424, CI => mult_28_C95_n422, CO => 
                           mult_28_C95_n417, S => mult_28_C95_n418);
   mult_28_C95_U586 : OAI22D1 port map( A1 => mult_28_C95_n24, A2 => 
                           mult_28_C95_n724, B1 => mult_28_C95_n723, B2 => 
                           mult_28_C95_n22, Z => mult_28_C95_n589);
   mult_28_C95_U402 : ADFULD1 port map( A => mult_28_C95_n451, B => 
                           mult_28_C95_n531, CI => mult_28_C95_n545, CO => 
                           mult_28_C95_n439, S => mult_28_C95_n440);
   mult_28_C95_U370 : ADFULD1 port map( A => mult_28_C95_n382, B => 
                           mult_28_C95_n384, CI => mult_28_C95_n391, CO => 
                           mult_28_C95_n377, S => mult_28_C95_n378);
   mult_28_C95_U379 : ADFULD1 port map( A => mult_28_C95_n572, B => 
                           mult_28_C95_n557, CI => mult_28_C95_n411, CO => 
                           mult_28_C95_n395, S => mult_28_C95_n396);
   mult_28_C95_U387 : ADFULD1 port map( A => mult_28_C95_n414, B => 
                           mult_28_C95_n543, CI => mult_28_C95_n558, CO => 
                           mult_28_C95_n411, S => mult_28_C95_n412);
   mult_28_C95_U519 : OAI22D1 port map( A1 => mult_28_C95_n693, A2 => 
                           mult_28_C95_n36, B1 => mult_28_C95_n692, B2 => 
                           mult_28_C95_n34, Z => mult_28_C95_n558);
   mult_28_C95_U486 : OAI22D1 port map( A1 => mult_28_C95_n678, A2 => 
                           mult_28_C95_n42, B1 => mult_28_C95_n677, B2 => 
                           mult_28_C95_n40, Z => mult_28_C95_n543);
   mult_28_C95_U518 : OAI22D1 port map( A1 => mult_28_C95_n692, A2 => 
                           mult_28_C95_n36, B1 => mult_28_C95_n691, B2 => 
                           mult_28_C95_n34, Z => mult_28_C95_n557);
   mult_28_C95_U520 : OAI22D1 port map( A1 => mult_28_C95_n694, A2 => 
                           mult_28_C95_n36, B1 => mult_28_C95_n693, B2 => 
                           mult_28_C95_n34, Z => mult_28_C95_n559);
   mult_28_C95_U748 : EXOR2D1 port map( A1 => coeff_memory_27_port, A2 => 
                           coeff_memory_26_port, Z => mult_28_C95_n803);
   mult_28_C95_U487 : OAI22D1 port map( A1 => mult_28_C95_n679, A2 => 
                           mult_28_C95_n42, B1 => mult_28_C95_n678, B2 => 
                           mult_28_C95_n40, Z => mult_28_C95_n544);
   mult_28_C95_U745 : EXOR2D1 port map( A1 => coeff_memory_29_port, A2 => 
                           coeff_memory_28_port, Z => mult_28_C95_n802);
   mult_28_C95_U502 : EXNOR2D1 port map( A1 => y_4_port, A2 => 
                           coeff_memory_29_port, Z => mult_28_C95_n677);
   mult_28_C95_U485 : OAI22D1 port map( A1 => mult_28_C95_n677, A2 => 
                           mult_28_C95_n42, B1 => mult_28_C95_n676, B2 => 
                           mult_28_C95_n40, Z => mult_28_C95_n542);
   mult_28_C95_U217 : AOI21D1 port map( A1 => mult_28_C95_n204, A2 => 
                           mult_28_C95_n212, B => mult_28_C95_n205, Z => 
                           mult_28_C95_n203);
   mult_28_C95_U751 : EXOR2D1 port map( A1 => coeff_memory_25_port, A2 => 
                           coeff_memory_24_port, Z => mult_28_C95_n804);
   mult_28_C95_U763 : EXOR2D1 port map( A1 => coeff_memory_17_port, A2 => 
                           coeff_memory_16_port, Z => mult_28_C95_n808);
   mult_28_C95_U760 : EXOR2D1 port map( A1 => coeff_memory_19_port, A2 => 
                           coeff_memory_18_port, Z => mult_28_C95_n807);
   mult_28_C95_U757 : EXOR2D1 port map( A1 => coeff_memory_21_port, A2 => 
                           coeff_memory_20_port, Z => mult_28_C95_n806);
   mult_28_C95_U754 : EXOR2D1 port map( A1 => coeff_memory_23_port, A2 => 
                           coeff_memory_22_port, Z => mult_28_C95_n805);
   mult_28_C95_U742 : EXOR2D1 port map( A1 => coeff_memory_31_port, A2 => 
                           coeff_memory_30_port, Z => mult_28_C95_n801);
   mult_28_C95_U717 : NAN2M1D1 port map( A1 => n39, A2 => coeff_memory_17_port,
                           Z => mult_28_C95_n784);
   mult_28_C95_U716 : EXNOR2D1 port map( A1 => n39, A2 => coeff_memory_17_port,
                           Z => mult_28_C95_n783);
   mult_28_C95_U699 : OAI22D1 port map( A1 => mult_28_C95_n783, A2 => 
                           mult_28_C95_n6, B1 => mult_28_C95_n782, B2 => 
                           mult_28_C95_n824, Z => mult_28_C95_n648);
   mult_28_C95_U698 : OAI22D1 port map( A1 => mult_28_C95_n782, A2 => 
                           mult_28_C95_n6, B1 => mult_28_C95_n781, B2 => 
                           mult_28_C95_n824, Z => mult_28_C95_n647);
   mult_28_C95_U696 : OAI22D1 port map( A1 => mult_28_C95_n780, A2 => 
                           mult_28_C95_n6, B1 => mult_28_C95_n779, B2 => 
                           mult_28_C95_n824, Z => mult_28_C95_n645);
   mult_28_C95_U695 : OAI22D1 port map( A1 => mult_28_C95_n779, A2 => 
                           mult_28_C95_n6, B1 => mult_28_C95_n778, B2 => 
                           mult_28_C95_n824, Z => mult_28_C95_n644);
   mult_28_C95_U694 : OAI22D1 port map( A1 => mult_28_C95_n778, A2 => 
                           mult_28_C95_n6, B1 => mult_28_C95_n777, B2 => 
                           mult_28_C95_n824, Z => mult_28_C95_n643);
   mult_28_C95_U693 : OAI22D1 port map( A1 => mult_28_C95_n777, A2 => 
                           mult_28_C95_n6, B1 => mult_28_C95_n776, B2 => 
                           mult_28_C95_n824, Z => mult_28_C95_n642);
   mult_28_C95_U692 : OAI22D1 port map( A1 => mult_28_C95_n776, A2 => 
                           mult_28_C95_n6, B1 => mult_28_C95_n775, B2 => 
                           mult_28_C95_n824, Z => mult_28_C95_n641);
   mult_28_C95_U691 : OAI22D1 port map( A1 => mult_28_C95_n775, A2 => 
                           mult_28_C95_n6, B1 => mult_28_C95_n774, B2 => 
                           mult_28_C95_n824, Z => mult_28_C95_n640);
   mult_28_C95_U689 : OAI22D1 port map( A1 => mult_28_C95_n773, A2 => 
                           mult_28_C95_n6, B1 => mult_28_C95_n772, B2 => 
                           mult_28_C95_n824, Z => mult_28_C95_n638);
   mult_28_C95_U688 : OAI22D1 port map( A1 => mult_28_C95_n772, A2 => 
                           mult_28_C95_n6, B1 => mult_28_C95_n771, B2 => 
                           mult_28_C95_n824, Z => mult_28_C95_n637);
   mult_28_C95_U687 : OAI22D1 port map( A1 => mult_28_C95_n771, A2 => 
                           mult_28_C95_n6, B1 => mult_28_C95_n770, B2 => 
                           mult_28_C95_n824, Z => mult_28_C95_n636);
   mult_28_C95_U686 : OAI22D1 port map( A1 => mult_28_C95_n770, A2 => 
                           mult_28_C95_n6, B1 => mult_28_C95_n769, B2 => 
                           mult_28_C95_n824, Z => mult_28_C95_n635);
   mult_28_C95_U683 : OAI22D1 port map( A1 => mult_28_C95_n6, A2 => 
                           mult_28_C95_n832, B1 => mult_28_C95_n784, B2 => 
                           mult_28_C95_n824, Z => mult_28_C95_n520);
   mult_28_C95_U682 : NAN2M1D1 port map( A1 => n39, A2 => coeff_memory_19_port,
                           Z => mult_28_C95_n767);
   mult_28_C95_U681 : EXNOR2D1 port map( A1 => n39, A2 => coeff_memory_19_port,
                           Z => mult_28_C95_n766);
   mult_28_C95_U665 : NOR2M1D1 port map( A1 => n39, A2 => mult_28_C95_n9, Z => 
                           mult_28_C95_n632);
   mult_28_C95_U664 : OAI22D1 port map( A1 => mult_28_C95_n766, A2 => 
                           mult_28_C95_n12, B1 => mult_28_C95_n765, B2 => 
                           mult_28_C95_n9, Z => mult_28_C95_n631);
   mult_28_C95_U661 : OAI22D1 port map( A1 => mult_28_C95_n763, A2 => 
                           mult_28_C95_n12, B1 => mult_28_C95_n762, B2 => 
                           mult_28_C95_n9, Z => mult_28_C95_n628);
   mult_28_C95_U660 : OAI22D1 port map( A1 => mult_28_C95_n762, A2 => 
                           mult_28_C95_n12, B1 => mult_28_C95_n761, B2 => 
                           mult_28_C95_n9, Z => mult_28_C95_n627);
   mult_28_C95_U659 : OAI22D1 port map( A1 => mult_28_C95_n761, A2 => 
                           mult_28_C95_n12, B1 => mult_28_C95_n760, B2 => 
                           mult_28_C95_n9, Z => mult_28_C95_n626);
   mult_28_C95_U658 : OAI22D1 port map( A1 => mult_28_C95_n760, A2 => 
                           mult_28_C95_n12, B1 => mult_28_C95_n759, B2 => 
                           mult_28_C95_n9, Z => mult_28_C95_n625);
   mult_28_C95_U657 : OAI22D1 port map( A1 => mult_28_C95_n759, A2 => 
                           mult_28_C95_n12, B1 => mult_28_C95_n758, B2 => 
                           mult_28_C95_n9, Z => mult_28_C95_n624);
   mult_28_C95_U656 : OAI22D1 port map( A1 => mult_28_C95_n758, A2 => 
                           mult_28_C95_n12, B1 => mult_28_C95_n757, B2 => 
                           mult_28_C95_n9, Z => mult_28_C95_n623);
   mult_28_C95_U655 : OAI22D1 port map( A1 => mult_28_C95_n756, A2 => 
                           mult_28_C95_n9, B1 => mult_28_C95_n757, B2 => 
                           mult_28_C95_n12, Z => mult_28_C95_n622);
   mult_28_C95_U654 : OAI22D1 port map( A1 => mult_28_C95_n756, A2 => 
                           mult_28_C95_n12, B1 => mult_28_C95_n755, B2 => 
                           mult_28_C95_n9, Z => mult_28_C95_n621);
   mult_28_C95_U653 : OAI22D1 port map( A1 => mult_28_C95_n755, A2 => 
                           mult_28_C95_n12, B1 => mult_28_C95_n754, B2 => 
                           mult_28_C95_n9, Z => mult_28_C95_n620);
   mult_28_C95_U651 : OAI22D1 port map( A1 => mult_28_C95_n753, A2 => 
                           mult_28_C95_n12, B1 => mult_28_C95_n752, B2 => 
                           mult_28_C95_n9, Z => mult_28_C95_n618);
   mult_28_C95_U649 : AO21D2 port map( A1 => mult_28_C95_n12, A2 => 
                           mult_28_C95_n9, B => mult_28_C95_n751, Z => 
                           mult_28_C95_n616);
   mult_28_C95_U648 : OAI22D1 port map( A1 => mult_28_C95_n12, A2 => 
                           mult_28_C95_n831, B1 => mult_28_C95_n767, B2 => 
                           mult_28_C95_n9, Z => mult_28_C95_n519);
   mult_28_C95_U647 : NAN2M1D1 port map( A1 => n39, A2 => coeff_memory_21_port,
                           Z => mult_28_C95_n750);
   mult_28_C95_U646 : EXNOR2D1 port map( A1 => n39, A2 => coeff_memory_21_port,
                           Z => mult_28_C95_n749);
   mult_28_C95_U642 : EXNOR2D1 port map( A1 => y_4_port, A2 => 
                           coeff_memory_21_port, Z => mult_28_C95_n745);
   mult_28_C95_U630 : NOR2M1D1 port map( A1 => n39, A2 => mult_28_C95_n16, Z =>
                           mult_28_C95_n615);
   mult_28_C95_U629 : OAI22D1 port map( A1 => mult_28_C95_n749, A2 => 
                           mult_28_C95_n18, B1 => mult_28_C95_n748, B2 => 
                           mult_28_C95_n16, Z => mult_28_C95_n614);
   mult_28_C95_U626 : OAI22D1 port map( A1 => mult_28_C95_n746, A2 => 
                           mult_28_C95_n18, B1 => mult_28_C95_n745, B2 => 
                           mult_28_C95_n16, Z => mult_28_C95_n611);
   mult_28_C95_U625 : OAI22D1 port map( A1 => mult_28_C95_n745, A2 => 
                           mult_28_C95_n18, B1 => mult_28_C95_n744, B2 => 
                           mult_28_C95_n16, Z => mult_28_C95_n610);
   mult_28_C95_U624 : OAI22D1 port map( A1 => mult_28_C95_n744, A2 => 
                           mult_28_C95_n18, B1 => mult_28_C95_n743, B2 => 
                           mult_28_C95_n16, Z => mult_28_C95_n609);
   mult_28_C95_U623 : OAI22D1 port map( A1 => mult_28_C95_n743, A2 => 
                           mult_28_C95_n18, B1 => mult_28_C95_n742, B2 => 
                           mult_28_C95_n16, Z => mult_28_C95_n608);
   mult_28_C95_U620 : OAI22D1 port map( A1 => mult_28_C95_n739, A2 => 
                           mult_28_C95_n16, B1 => mult_28_C95_n740, B2 => 
                           mult_28_C95_n18, Z => mult_28_C95_n605);
   mult_28_C95_U617 : OAI22D1 port map( A1 => mult_28_C95_n737, A2 => 
                           mult_28_C95_n18, B1 => mult_28_C95_n736, B2 => 
                           mult_28_C95_n16, Z => mult_28_C95_n602);
   mult_28_C95_U616 : OAI22D1 port map( A1 => mult_28_C95_n736, A2 => 
                           mult_28_C95_n18, B1 => mult_28_C95_n735, B2 => 
                           mult_28_C95_n16, Z => mult_28_C95_n601);
   mult_28_C95_U613 : OAI22D1 port map( A1 => mult_28_C95_n18, A2 => 
                           mult_28_C95_n830, B1 => mult_28_C95_n750, B2 => 
                           mult_28_C95_n16, Z => mult_28_C95_n518);
   mult_28_C95_U612 : NAN2M1D1 port map( A1 => n39, A2 => coeff_memory_23_port,
                           Z => mult_28_C95_n733);
   mult_28_C95_U611 : EXNOR2D1 port map( A1 => n39, A2 => coeff_memory_23_port,
                           Z => mult_28_C95_n732);
   mult_28_C95_U607 : EXNOR2D1 port map( A1 => y_4_port, A2 => 
                           coeff_memory_23_port, Z => mult_28_C95_n728);
   mult_28_C95_U595 : NOR2M1D1 port map( A1 => n39, A2 => mult_28_C95_n22, Z =>
                           mult_28_C95_n598);
   mult_28_C95_U594 : OAI22D1 port map( A1 => mult_28_C95_n732, A2 => 
                           mult_28_C95_n24, B1 => mult_28_C95_n731, B2 => 
                           mult_28_C95_n22, Z => mult_28_C95_n597);
   mult_28_C95_U591 : OAI22D1 port map( A1 => mult_28_C95_n729, A2 => 
                           mult_28_C95_n24, B1 => mult_28_C95_n728, B2 => 
                           mult_28_C95_n22, Z => mult_28_C95_n594);
   mult_28_C95_U589 : OAI22D1 port map( A1 => mult_28_C95_n727, A2 => 
                           mult_28_C95_n24, B1 => mult_28_C95_n726, B2 => 
                           mult_28_C95_n22, Z => mult_28_C95_n592);
   mult_28_C95_U587 : OAI22D1 port map( A1 => mult_28_C95_n725, A2 => 
                           mult_28_C95_n24, B1 => mult_28_C95_n724, B2 => 
                           mult_28_C95_n22, Z => mult_28_C95_n590);
   mult_28_C95_U585 : OAI22D1 port map( A1 => mult_28_C95_n722, A2 => 
                           mult_28_C95_n22, B1 => mult_28_C95_n723, B2 => 
                           mult_28_C95_n24, Z => mult_28_C95_n588);
   mult_28_C95_U584 : OAI22D1 port map( A1 => mult_28_C95_n722, A2 => 
                           mult_28_C95_n24, B1 => mult_28_C95_n721, B2 => 
                           mult_28_C95_n22, Z => mult_28_C95_n587);
   mult_28_C95_U583 : OAI22D1 port map( A1 => mult_28_C95_n721, A2 => 
                           mult_28_C95_n24, B1 => mult_28_C95_n720, B2 => 
                           mult_28_C95_n22, Z => mult_28_C95_n586);
   mult_28_C95_U582 : OAI22D1 port map( A1 => mult_28_C95_n720, A2 => 
                           mult_28_C95_n24, B1 => mult_28_C95_n719, B2 => 
                           mult_28_C95_n22, Z => mult_28_C95_n585);
   mult_28_C95_U581 : OAI22D1 port map( A1 => mult_28_C95_n719, A2 => 
                           mult_28_C95_n24, B1 => mult_28_C95_n718, B2 => 
                           mult_28_C95_n22, Z => mult_28_C95_n584);
   mult_28_C95_U578 : OAI22D1 port map( A1 => mult_28_C95_n24, A2 => 
                           mult_28_C95_n829, B1 => mult_28_C95_n733, B2 => 
                           mult_28_C95_n22, Z => mult_28_C95_n517);
   mult_28_C95_U577 : NAN2M1D1 port map( A1 => n39, A2 => coeff_memory_25_port,
                           Z => mult_28_C95_n716);
   mult_28_C95_U576 : EXNOR2D1 port map( A1 => n39, A2 => coeff_memory_25_port,
                           Z => mult_28_C95_n715);
   mult_28_C95_U572 : EXNOR2D1 port map( A1 => y_4_port, A2 => 
                           coeff_memory_25_port, Z => mult_28_C95_n711);
   mult_28_C95_U560 : NOR2M1D1 port map( A1 => n39, A2 => mult_28_C95_n28, Z =>
                           mult_28_C95_n581);
   mult_28_C95_U559 : OAI22D1 port map( A1 => mult_28_C95_n715, A2 => 
                           mult_28_C95_n30, B1 => mult_28_C95_n714, B2 => 
                           mult_28_C95_n28, Z => mult_28_C95_n580);
   mult_28_C95_U556 : OAI22D1 port map( A1 => mult_28_C95_n712, A2 => 
                           mult_28_C95_n30, B1 => mult_28_C95_n711, B2 => 
                           mult_28_C95_n28, Z => mult_28_C95_n577);
   mult_28_C95_U555 : OAI22D1 port map( A1 => mult_28_C95_n711, A2 => 
                           mult_28_C95_n30, B1 => mult_28_C95_n710, B2 => 
                           mult_28_C95_n28, Z => mult_28_C95_n576);
   mult_28_C95_U554 : OAI22D1 port map( A1 => mult_28_C95_n710, A2 => 
                           mult_28_C95_n30, B1 => mult_28_C95_n709, B2 => 
                           mult_28_C95_n28, Z => mult_28_C95_n575);
   mult_28_C95_U553 : OAI22D1 port map( A1 => mult_28_C95_n709, A2 => 
                           mult_28_C95_n30, B1 => mult_28_C95_n708, B2 => 
                           mult_28_C95_n28, Z => mult_28_C95_n574);
   mult_28_C95_U550 : OAI22D1 port map( A1 => mult_28_C95_n705, A2 => 
                           mult_28_C95_n28, B1 => mult_28_C95_n706, B2 => 
                           mult_28_C95_n30, Z => mult_28_C95_n571);
   mult_28_C95_U549 : OAI22D1 port map( A1 => mult_28_C95_n30, A2 => 
                           mult_28_C95_n705, B1 => mult_28_C95_n704, B2 => 
                           mult_28_C95_n28, Z => mult_28_C95_n570);
   mult_28_C95_U548 : OAI22D1 port map( A1 => mult_28_C95_n704, A2 => 
                           mult_28_C95_n30, B1 => mult_28_C95_n703, B2 => 
                           mult_28_C95_n28, Z => mult_28_C95_n569);
   mult_28_C95_U547 : OAI22D1 port map( A1 => mult_28_C95_n703, A2 => 
                           mult_28_C95_n30, B1 => mult_28_C95_n702, B2 => 
                           mult_28_C95_n28, Z => mult_28_C95_n568);
   mult_28_C95_U546 : OAI22D1 port map( A1 => mult_28_C95_n702, A2 => 
                           mult_28_C95_n30, B1 => mult_28_C95_n701, B2 => 
                           mult_28_C95_n28, Z => mult_28_C95_n567);
   mult_28_C95_U543 : OAI22D1 port map( A1 => mult_28_C95_n30, A2 => 
                           mult_28_C95_n828, B1 => mult_28_C95_n716, B2 => 
                           mult_28_C95_n28, Z => mult_28_C95_n516);
   mult_28_C95_U542 : NAN2M1D1 port map( A1 => n39, A2 => coeff_memory_27_port,
                           Z => mult_28_C95_n699);
   mult_28_C95_U541 : EXNOR2D1 port map( A1 => n39, A2 => coeff_memory_27_port,
                           Z => mult_28_C95_n698);
   mult_28_C95_U537 : EXNOR2D1 port map( A1 => y_4_port, A2 => 
                           coeff_memory_27_port, Z => mult_28_C95_n694);
   mult_28_C95_U525 : NOR2M1D1 port map( A1 => n39, A2 => mult_28_C95_n34, Z =>
                           mult_28_C95_n564);
   mult_28_C95_U524 : OAI22D1 port map( A1 => mult_28_C95_n698, A2 => 
                           mult_28_C95_n36, B1 => mult_28_C95_n697, B2 => 
                           mult_28_C95_n34, Z => mult_28_C95_n563);
   mult_28_C95_U522 : OAI22D1 port map( A1 => mult_28_C95_n696, A2 => 
                           mult_28_C95_n36, B1 => mult_28_C95_n695, B2 => 
                           mult_28_C95_n34, Z => mult_28_C95_n561);
   mult_28_C95_U521 : OAI22D1 port map( A1 => mult_28_C95_n695, A2 => 
                           mult_28_C95_n36, B1 => mult_28_C95_n694, B2 => 
                           mult_28_C95_n34, Z => mult_28_C95_n560);
   mult_28_C95_U517 : OAI22D1 port map( A1 => mult_28_C95_n691, A2 => 
                           mult_28_C95_n36, B1 => mult_28_C95_n690, B2 => 
                           mult_28_C95_n34, Z => mult_28_C95_n556);
   mult_28_C95_U516 : OAI22D1 port map( A1 => mult_28_C95_n690, A2 => 
                           mult_28_C95_n36, B1 => mult_28_C95_n689, B2 => 
                           mult_28_C95_n34, Z => mult_28_C95_n555);
   mult_28_C95_U515 : OAI22D1 port map( A1 => mult_28_C95_n688, A2 => 
                           mult_28_C95_n34, B1 => mult_28_C95_n689, B2 => 
                           mult_28_C95_n36, Z => mult_28_C95_n554);
   mult_28_C95_U513 : OAI22D1 port map( A1 => mult_28_C95_n687, A2 => 
                           mult_28_C95_n36, B1 => mult_28_C95_n686, B2 => 
                           mult_28_C95_n34, Z => mult_28_C95_n552);
   mult_28_C95_U512 : OAI22D1 port map( A1 => mult_28_C95_n686, A2 => 
                           mult_28_C95_n36, B1 => mult_28_C95_n685, B2 => 
                           mult_28_C95_n34, Z => mult_28_C95_n551);
   mult_28_C95_U511 : OAI22D1 port map( A1 => mult_28_C95_n685, A2 => 
                           mult_28_C95_n36, B1 => mult_28_C95_n684, B2 => 
                           mult_28_C95_n34, Z => mult_28_C95_n550);
   mult_28_C95_U508 : OAI22D1 port map( A1 => mult_28_C95_n36, A2 => 
                           mult_28_C95_n827, B1 => mult_28_C95_n699, B2 => 
                           mult_28_C95_n34, Z => mult_28_C95_n515);
   mult_28_C95_U507 : NAN2M1D1 port map( A1 => n39, A2 => coeff_memory_29_port,
                           Z => mult_28_C95_n682);
   mult_28_C95_U506 : EXNOR2D1 port map( A1 => n39, A2 => coeff_memory_29_port,
                           Z => mult_28_C95_n681);
   mult_28_C95_U490 : NOR2M1D1 port map( A1 => n39, A2 => mult_28_C95_n40, Z =>
                           mult_28_C95_n547);
   mult_28_C95_U489 : OAI22D1 port map( A1 => mult_28_C95_n681, A2 => 
                           mult_28_C95_n42, B1 => mult_28_C95_n680, B2 => 
                           mult_28_C95_n40, Z => mult_28_C95_n546);
   mult_28_C95_U484 : OAI22D1 port map( A1 => mult_28_C95_n676, A2 => 
                           mult_28_C95_n42, B1 => mult_28_C95_n675, B2 => 
                           mult_28_C95_n40, Z => mult_28_C95_n541);
   mult_28_C95_U483 : OAI22D1 port map( A1 => mult_28_C95_n675, A2 => 
                           mult_28_C95_n42, B1 => mult_28_C95_n674, B2 => 
                           mult_28_C95_n40, Z => mult_28_C95_n540);
   mult_28_C95_U482 : OAI22D1 port map( A1 => mult_28_C95_n674, A2 => 
                           mult_28_C95_n42, B1 => mult_28_C95_n673, B2 => 
                           mult_28_C95_n40, Z => mult_28_C95_n539);
   mult_28_C95_U481 : OAI22D1 port map( A1 => mult_28_C95_n673, A2 => 
                           mult_28_C95_n42, B1 => mult_28_C95_n672, B2 => 
                           mult_28_C95_n40, Z => mult_28_C95_n538);
   mult_28_C95_U480 : OAI22D1 port map( A1 => mult_28_C95_n671, A2 => 
                           mult_28_C95_n40, B1 => mult_28_C95_n672, B2 => 
                           mult_28_C95_n42, Z => mult_28_C95_n537);
   mult_28_C95_U479 : OAI22D1 port map( A1 => mult_28_C95_n42, A2 => 
                           mult_28_C95_n671, B1 => mult_28_C95_n670, B2 => 
                           mult_28_C95_n40, Z => mult_28_C95_n536);
   mult_28_C95_U477 : OAI22D1 port map( A1 => mult_28_C95_n669, A2 => 
                           mult_28_C95_n42, B1 => mult_28_C95_n668, B2 => 
                           mult_28_C95_n40, Z => mult_28_C95_n534);
   mult_28_C95_U475 : OAI22D1 port map( A1 => mult_28_C95_n667, A2 => 
                           mult_28_C95_n42, B1 => mult_28_C95_n666, B2 => 
                           mult_28_C95_n40, Z => mult_28_C95_n309);
   mult_28_C95_U473 : OAI22D1 port map( A1 => mult_28_C95_n42, A2 => 
                           mult_28_C95_n826, B1 => mult_28_C95_n682, B2 => 
                           mult_28_C95_n40, Z => mult_28_C95_n514);
   mult_28_C95_U472 : NAN2M1D1 port map( A1 => n39, A2 => coeff_memory_31_port,
                           Z => mult_28_C95_n665);
   mult_28_C95_U471 : EXNOR2D1 port map( A1 => n39, A2 => coeff_memory_31_port,
                           Z => mult_28_C95_n664);
   mult_28_C95_U455 : NOR2M1D1 port map( A1 => n39, A2 => mult_28_C95_n46, Z =>
                           mult_28_C95_n531);
   mult_28_C95_U454 : OAI22D1 port map( A1 => mult_28_C95_n664, A2 => 
                           mult_28_C95_n48, B1 => mult_28_C95_n663, B2 => 
                           mult_28_C95_n46, Z => mult_28_C95_n530);
   mult_28_C95_U451 : OAI22D1 port map( A1 => mult_28_C95_n661, A2 => 
                           mult_28_C95_n48, B1 => mult_28_C95_n660, B2 => 
                           mult_28_C95_n46, Z => mult_28_C95_n528);
   mult_28_C95_U450 : OAI22D1 port map( A1 => mult_28_C95_n660, A2 => 
                           mult_28_C95_n48, B1 => mult_28_C95_n659, B2 => 
                           mult_28_C95_n46, Z => mult_28_C95_n373);
   mult_28_C95_U449 : OAI22D1 port map( A1 => mult_28_C95_n659, A2 => 
                           mult_28_C95_n48, B1 => mult_28_C95_n658, B2 => 
                           mult_28_C95_n46, Z => mult_28_C95_n527);
   mult_28_C95_U448 : OAI22D1 port map( A1 => mult_28_C95_n658, A2 => 
                           mult_28_C95_n48, B1 => mult_28_C95_n657, B2 => 
                           mult_28_C95_n46, Z => mult_28_C95_n351);
   mult_28_C95_U445 : OAI22D1 port map( A1 => mult_28_C95_n654, A2 => 
                           mult_28_C95_n46, B1 => mult_28_C95_n655, B2 => 
                           mult_28_C95_n48, Z => mult_28_C95_n525);
   mult_28_C95_U444 : OAI22D1 port map( A1 => mult_28_C95_n654, A2 => 
                           mult_28_C95_n48, B1 => mult_28_C95_n653, B2 => 
                           mult_28_C95_n46, Z => mult_28_C95_n319);
   mult_28_C95_U441 : OAI22D1 port map( A1 => mult_28_C95_n651, A2 => 
                           mult_28_C95_n48, B1 => mult_28_C95_n650, B2 => 
                           mult_28_C95_n46, Z => mult_28_C95_n522);
   mult_28_C95_U439 : OAI22D1 port map( A1 => mult_28_C95_n48, A2 => 
                           mult_28_C95_n920, B1 => mult_28_C95_n665, B2 => 
                           mult_28_C95_n46, Z => mult_28_C95_n513);
   mult_28_C95_U435 : ADFULD1 port map( A => mult_28_C95_n629, B => 
                           mult_28_C95_n508, CI => mult_28_C95_n644, CO => 
                           mult_28_C95_n505, S => mult_28_C95_n506);
   mult_28_C95_U434 : ADFULD1 port map( A => mult_28_C95_n507, B => 
                           mult_28_C95_n598, CI => mult_28_C95_n613, CO => 
                           mult_28_C95_n503, S => mult_28_C95_n504);
   mult_28_C95_U433 : ADFULD1 port map( A => mult_28_C95_n643, B => 
                           mult_28_C95_n628, CI => mult_28_C95_n504, CO => 
                           mult_28_C95_n501, S => mult_28_C95_n502);
   mult_28_C95_U431 : ADFULD1 port map( A => mult_28_C95_n612, B => 
                           mult_28_C95_n500, CI => mult_28_C95_n627, CO => 
                           mult_28_C95_n497, S => mult_28_C95_n498);
   mult_28_C95_U430 : ADFULD1 port map( A => mult_28_C95_n642, B => 
                           mult_28_C95_n503, CI => mult_28_C95_n498, CO => 
                           mult_28_C95_n495, S => mult_28_C95_n496);
   mult_28_C95_U429 : ADFULD1 port map( A => mult_28_C95_n499, B => 
                           mult_28_C95_n581, CI => mult_28_C95_n596, CO => 
                           mult_28_C95_n493, S => mult_28_C95_n494);
   mult_28_C95_U428 : ADFULD1 port map( A => mult_28_C95_n626, B => 
                           mult_28_C95_n611, CI => mult_28_C95_n494, CO => 
                           mult_28_C95_n491, S => mult_28_C95_n492);
   mult_28_C95_U427 : ADFULD1 port map( A => mult_28_C95_n641, B => 
                           mult_28_C95_n497, CI => mult_28_C95_n492, CO => 
                           mult_28_C95_n489, S => mult_28_C95_n490);
   mult_28_C95_U425 : ADFULD1 port map( A => mult_28_C95_n595, B => 
                           mult_28_C95_n488, CI => mult_28_C95_n610, CO => 
                           mult_28_C95_n485, S => mult_28_C95_n486);
   mult_28_C95_U424 : ADFULD1 port map( A => mult_28_C95_n625, B => 
                           mult_28_C95_n493, CI => mult_28_C95_n640, CO => 
                           mult_28_C95_n483, S => mult_28_C95_n484);
   mult_28_C95_U423 : ADFULD1 port map( A => mult_28_C95_n491, B => 
                           mult_28_C95_n486, CI => mult_28_C95_n484, CO => 
                           mult_28_C95_n481, S => mult_28_C95_n482);
   mult_28_C95_U422 : ADFULD1 port map( A => mult_28_C95_n487, B => 
                           mult_28_C95_n564, CI => mult_28_C95_n579, CO => 
                           mult_28_C95_n479, S => mult_28_C95_n480);
   mult_28_C95_U421 : ADFULD1 port map( A => mult_28_C95_n609, B => 
                           mult_28_C95_n594, CI => mult_28_C95_n480, CO => 
                           mult_28_C95_n477, S => mult_28_C95_n478);
   mult_28_C95_U416 : ADFULD1 port map( A => mult_28_C95_n608, B => 
                           mult_28_C95_n479, CI => mult_28_C95_n623, CO => 
                           mult_28_C95_n467, S => mult_28_C95_n468);
   mult_28_C95_U415 : ADFULD1 port map( A => mult_28_C95_n470, B => 
                           mult_28_C95_n638, CI => mult_28_C95_n477, CO => 
                           mult_28_C95_n465, S => mult_28_C95_n466);
   mult_28_C95_U414 : ADFULD1 port map( A => mult_28_C95_n468, B => 
                           mult_28_C95_n475, CI => mult_28_C95_n466, CO => 
                           mult_28_C95_n463, S => mult_28_C95_n464);
   mult_28_C95_U413 : ADFULD1 port map( A => mult_28_C95_n471, B => 
                           mult_28_C95_n547, CI => mult_28_C95_n562, CO => 
                           mult_28_C95_n461, S => mult_28_C95_n462);
   mult_28_C95_U412 : ADFULD1 port map( A => mult_28_C95_n592, B => 
                           mult_28_C95_n577, CI => mult_28_C95_n462, CO => 
                           mult_28_C95_n459, S => mult_28_C95_n460);
   mult_28_C95_U410 : ADFULD1 port map( A => mult_28_C95_n460, B => 
                           mult_28_C95_n637, CI => mult_28_C95_n467, CO => 
                           mult_28_C95_n455, S => mult_28_C95_n456);
   mult_28_C95_U409 : ADFULD1 port map( A => mult_28_C95_n458, B => 
                           mult_28_C95_n465, CI => mult_28_C95_n456, CO => 
                           mult_28_C95_n453, S => mult_28_C95_n454);
   mult_28_C95_U407 : ADFULD1 port map( A => mult_28_C95_n561, B => 
                           mult_28_C95_n452, CI => mult_28_C95_n576, CO => 
                           mult_28_C95_n449, S => mult_28_C95_n450);
   mult_28_C95_U405 : ADFULD1 port map( A => mult_28_C95_n450, B => 
                           mult_28_C95_n621, CI => mult_28_C95_n636, CO => 
                           mult_28_C95_n445, S => mult_28_C95_n446);
   mult_28_C95_U398 : ADFULD1 port map( A => mult_28_C95_n447, B => 
                           mult_28_C95_n445, CI => mult_28_C95_n436, CO => 
                           mult_28_C95_n431, S => mult_28_C95_n432);
   mult_28_C95_U397 : ADFULD1 port map( A => mult_28_C95_n443, B => 
                           mult_28_C95_n434, CI => mult_28_C95_n432, CO => 
                           mult_28_C95_n429, S => mult_28_C95_n430);
   mult_28_C95_U390 : ADFULD1 port map( A => mult_28_C95_n431, B => 
                           mult_28_C95_n420, CI => mult_28_C95_n418, CO => 
                           mult_28_C95_n415, S => mult_28_C95_n416);
   mult_28_C95_U380 : ADFULD1 port map( A => mult_28_C95_n400, B => 
                           mult_28_C95_n413, CI => mult_28_C95_n542, CO => 
                           mult_28_C95_n397, S => mult_28_C95_n398);
   mult_28_C95_U378 : ADFULD1 port map( A => mult_28_C95_n398, B => 
                           mult_28_C95_n587, CI => mult_28_C95_n602, CO => 
                           mult_28_C95_n393, S => mult_28_C95_n394);
   mult_28_C95_U374 : ADFULD1 port map( A => mult_28_C95_n528, B => 
                           mult_28_C95_n399, CI => mult_28_C95_n541, CO => 
                           mult_28_C95_n385, S => mult_28_C95_n386);
   mult_28_C95_U372 : ADFULD1 port map( A => mult_28_C95_n386, B => 
                           mult_28_C95_n586, CI => mult_28_C95_n601, CO => 
                           mult_28_C95_n381, S => mult_28_C95_n382);
   mult_28_C95_U367 : ADFULD1 port map( A => mult_28_C95_n540, B => 
                           mult_28_C95_n374, CI => mult_28_C95_n555, CO => 
                           mult_28_C95_n371, S => mult_28_C95_n372);
   mult_28_C95_U366 : ADFULD1 port map( A => mult_28_C95_n570, B => 
                           mult_28_C95_n385, CI => mult_28_C95_n600, CO => 
                           mult_28_C95_n369, S => mult_28_C95_n370);
   mult_28_C95_U365 : ADFULD1 port map( A => mult_28_C95_n383, B => 
                           mult_28_C95_n585, CI => mult_28_C95_n372, CO => 
                           mult_28_C95_n367, S => mult_28_C95_n368);
   mult_28_C95_U362 : ADFULD1 port map( A => mult_28_C95_n527, B => 
                           mult_28_C95_n373, CI => mult_28_C95_n554, CO => 
                           mult_28_C95_n361, S => mult_28_C95_n362);
   mult_28_C95_U361 : ADFULD1 port map( A => mult_28_C95_n569, B => 
                           mult_28_C95_n539, CI => mult_28_C95_n584, CO => 
                           mult_28_C95_n359, S => mult_28_C95_n360);
   mult_28_C95_U360 : ADFULD1 port map( A => mult_28_C95_n371, B => 
                           mult_28_C95_n599, CI => mult_28_C95_n362, CO => 
                           mult_28_C95_n357, S => mult_28_C95_n358);
   mult_28_C95_U359 : ADFULD1 port map( A => mult_28_C95_n360, B => 
                           mult_28_C95_n369, CI => mult_28_C95_n367, CO => 
                           mult_28_C95_n355, S => mult_28_C95_n356);
   mult_28_C95_U358 : ADFULD1 port map( A => mult_28_C95_n365, B => 
                           mult_28_C95_n358, CI => mult_28_C95_n356, CO => 
                           mult_28_C95_n353, S => mult_28_C95_n354);
   mult_28_C95_U356 : ADFULD1 port map( A => mult_28_C95_n352, B => 
                           mult_28_C95_n538, CI => mult_28_C95_n553, CO => 
                           mult_28_C95_n349, S => mult_28_C95_n350);
   mult_28_C95_U355 : ADFULD1 port map( A => mult_28_C95_n568, B => 
                           mult_28_C95_n583, CI => mult_28_C95_n361, CO => 
                           mult_28_C95_n347, S => mult_28_C95_n348);
   mult_28_C95_U354 : ADFULD1 port map( A => mult_28_C95_n350, B => 
                           mult_28_C95_n359, CI => mult_28_C95_n357, CO => 
                           mult_28_C95_n345, S => mult_28_C95_n346);
   mult_28_C95_U353 : ADFULD1 port map( A => mult_28_C95_n355, B => 
                           mult_28_C95_n348, CI => mult_28_C95_n346, CO => 
                           mult_28_C95_n343, S => mult_28_C95_n344);
   mult_28_C95_U352 : ADFULD1 port map( A => mult_28_C95_n537, B => 
                           mult_28_C95_n351, CI => mult_28_C95_n526, CO => 
                           mult_28_C95_n341, S => mult_28_C95_n342);
   mult_28_C95_U351 : ADFULD1 port map( A => mult_28_C95_n567, B => 
                           mult_28_C95_n552, CI => mult_28_C95_n582, CO => 
                           mult_28_C95_n339, S => mult_28_C95_n340);
   mult_28_C95_U350 : ADFULD1 port map( A => mult_28_C95_n342, B => 
                           mult_28_C95_n349, CI => mult_28_C95_n347, CO => 
                           mult_28_C95_n337, S => mult_28_C95_n338);
   mult_28_C95_U349 : ADFULD1 port map( A => mult_28_C95_n345, B => 
                           mult_28_C95_n340, CI => mult_28_C95_n338, CO => 
                           mult_28_C95_n335, S => mult_28_C95_n336);
   mult_28_C95_U347 : ADFULD1 port map( A => mult_28_C95_n536, B => 
                           mult_28_C95_n334, CI => mult_28_C95_n551, CO => 
                           mult_28_C95_n331, S => mult_28_C95_n332);
   mult_28_C95_U346 : ADFULD1 port map( A => mult_28_C95_n341, B => 
                           mult_28_C95_n566, CI => mult_28_C95_n339, CO => 
                           mult_28_C95_n329, S => mult_28_C95_n330);
   mult_28_C95_U345 : ADFULD1 port map( A => mult_28_C95_n337, B => 
                           mult_28_C95_n332, CI => mult_28_C95_n330, CO => 
                           mult_28_C95_n327, S => mult_28_C95_n328);
   mult_28_C95_U344 : ADFULD1 port map( A => mult_28_C95_n333, B => 
                           mult_28_C95_n525, CI => mult_28_C95_n550, CO => 
                           mult_28_C95_n325, S => mult_28_C95_n326);
   mult_28_C95_U343 : ADFULD1 port map( A => mult_28_C95_n565, B => 
                           mult_28_C95_n535, CI => mult_28_C95_n331, CO => 
                           mult_28_C95_n323, S => mult_28_C95_n324);
   mult_28_C95_U342 : ADFULD1 port map( A => mult_28_C95_n329, B => 
                           mult_28_C95_n326, CI => mult_28_C95_n324, CO => 
                           mult_28_C95_n321, S => mult_28_C95_n322);
   mult_28_C95_U340 : ADFULD1 port map( A => mult_28_C95_n534, B => 
                           mult_28_C95_n549, CI => mult_28_C95_n320, CO => 
                           mult_28_C95_n317, S => mult_28_C95_n318);
   mult_28_C95_U339 : ADFULD1 port map( A => mult_28_C95_n318, B => 
                           mult_28_C95_n325, CI => mult_28_C95_n323, CO => 
                           mult_28_C95_n315, S => mult_28_C95_n316);
   mult_28_C95_U338 : ADFULD1 port map( A => mult_28_C95_n524, B => 
                           mult_28_C95_n319, CI => mult_28_C95_n548, CO => 
                           mult_28_C95_n313, S => mult_28_C95_n314);
   mult_28_C95_U337 : ADFULD1 port map( A => mult_28_C95_n317, B => 
                           mult_28_C95_n533, CI => mult_28_C95_n314, CO => 
                           mult_28_C95_n311, S => mult_28_C95_n312);
   mult_28_C95_U335 : ADFULD1 port map( A => mult_28_C95_n310, B => 
                           mult_28_C95_n523, CI => mult_28_C95_n313, CO => 
                           mult_28_C95_n307, S => mult_28_C95_n308);
   mult_28_C95_U334 : ADFULD1 port map( A => mult_28_C95_n522, B => 
                           mult_28_C95_n309, CI => mult_28_C95_n532, CO => 
                           mult_28_C95_n305, S => mult_28_C95_n306);
   mult_28_C95_U320 : AOI21D1 port map( A1 => mult_28_C95_n1006, A2 => 
                           mult_28_C95_n1008, B => mult_28_C95_n1007, Z => 
                           mult_28_C95_n267);
   mult_28_C95_U314 : OAI21D1 port map( A1 => mult_28_C95_n267, A2 => 
                           mult_28_C95_n265, B => mult_28_C95_n266, Z => 
                           mult_28_C95_n264);
   mult_28_C95_U306 : AOI21D1 port map( A1 => mult_28_C95_n1004, A2 => 
                           mult_28_C95_n264, B => mult_28_C95_n1005, Z => 
                           mult_28_C95_n259);
   mult_28_C95_U300 : OAI21D1 port map( A1 => mult_28_C95_n257, A2 => 
                           mult_28_C95_n259, B => mult_28_C95_n258, Z => 
                           mult_28_C95_n256);
   mult_28_C95_U292 : AOI21D1 port map( A1 => mult_28_C95_n256, A2 => 
                           mult_28_C95_n1002, B => mult_28_C95_n1003, Z => 
                           mult_28_C95_n251);
   mult_28_C95_U286 : OAI21D1 port map( A1 => mult_28_C95_n249, A2 => 
                           mult_28_C95_n251, B => mult_28_C95_n250, Z => 
                           mult_28_C95_n248);
   mult_28_C95_U278 : AOI21D1 port map( A1 => mult_28_C95_n248, A2 => 
                           mult_28_C95_n1000, B => mult_28_C95_n1001, Z => 
                           mult_28_C95_n243);
   mult_28_C95_U259 : OAI21D1 port map( A1 => mult_28_C95_n231, A2 => 
                           mult_28_C95_n243, B => mult_28_C95_n232, Z => 
                           mult_28_C95_n230);
   mult_28_C95_U234 : AOI21D1 port map( A1 => mult_28_C95_n990, A2 => 
                           mult_28_C95_n992, B => mult_28_C95_n994, Z => 
                           mult_28_C95_n214);
   mult_28_C95_U232 : OAI21D1 port map( A1 => mult_28_C95_n225, A2 => 
                           mult_28_C95_n213, B => mult_28_C95_n214, Z => 
                           mult_28_C95_n212);
   mult_28_C95_U228 : NOR2D2 port map( A1 => mult_28_C95_n430, A2 => 
                           mult_28_C95_n441, Z => mult_28_C95_n209);
   mult_28_C95_U224 : EXOR2D1 port map( A1 => mult_28_C95_n211, A2 => 
                           mult_28_C95_n69, Z => m3_0);
   mult_28_C95_U222 : NOR2D2 port map( A1 => mult_28_C95_n416, A2 => 
                           mult_28_C95_n429, Z => mult_28_C95_n206);
   mult_28_C95_U207 : EXNOR2D1 port map( A1 => mult_28_C95_n202, A2 => 
                           mult_28_C95_n67, Z => m3_2);
   mult_28_C95_U205 : NOR2D2 port map( A1 => mult_28_C95_n388, A2 => 
                           mult_28_C95_n401, Z => mult_28_C95_n195);
   mult_28_C95_U165 : NOR2D2 port map( A1 => mult_28_C95_n344, A2 => 
                           mult_28_C95_n353, Z => mult_28_C95_n167);
   mult_28_C95_U114 : AOI21D1 port map( A1 => mult_28_C95_net12285, A2 => 
                           mult_28_C95_n128, B => mult_28_C95_n129, Z => 
                           mult_28_C95_n127);
   mult_28_C95_U80 : OAI21D1 port map( A1 => mult_28_C95_n113, A2 => 
                           mult_28_C95_n103, B => mult_28_C95_n104, Z => 
                           mult_28_C95_n102);
   mult_28_C95_U78 : AOI21D1 port map( A1 => mult_28_C95_n101, A2 => 
                           mult_28_C95_n124, B => mult_28_C95_n102, Z => 
                           mult_28_C95_n100);
   mult_28_C95_U59 : EXOR2D1 port map( A1 => mult_28_C95_n94, A2 => 
                           mult_28_C95_n55, Z => m3_14);
   mult_28_C95_U54 : EXOR2D1 port map( A1 => mult_28_C95_n85, A2 => 
                           mult_28_C95_n54, Z => m3_15);
   mult_28_C96_U1329 : EXNOR2DL port map( A1 => y_11_port, A2 => 
                           coeff_memory_1_port, Z => mult_28_C96_n772);
   mult_28_C96_U1328 : EXNOR2DL port map( A1 => y_11_port, A2 => 
                           coeff_memory_11_port, Z => mult_28_C96_n687);
   mult_28_C96_U1327 : EXNOR2DL port map( A1 => y_11_port, A2 => 
                           coeff_memory_13_port, Z => mult_28_C96_n670);
   mult_28_C96_U1326 : EXNOR2DL port map( A1 => y_11_port, A2 => 
                           coeff_memory_15_port, Z => mult_28_C96_n653);
   mult_28_C96_U1325 : AOI21DL port map( A1 => mult_28_C96_n202, A2 => 
                           mult_28_C96_n968, B => mult_28_C96_n1057, Z => 
                           mult_28_C96_n188);
   mult_28_C96_U1324 : EXNOR2DL port map( A1 => y_13_port, A2 => 
                           coeff_memory_7_port, Z => mult_28_C96_n719);
   mult_28_C96_U1323 : EXNOR2DL port map( A1 => y_13_port, A2 => 
                           coeff_memory_9_port, Z => mult_28_C96_n702);
   mult_28_C96_U1322 : EXNOR2DL port map( A1 => y_13_port, A2 => 
                           coeff_memory_11_port, Z => mult_28_C96_n685);
   mult_28_C96_U1321 : EXNOR2DL port map( A1 => y_13_port, A2 => 
                           coeff_memory_13_port, Z => mult_28_C96_n668);
   mult_28_C96_U1320 : EXNOR2DL port map( A1 => y_13_port, A2 => 
                           coeff_memory_15_port, Z => mult_28_C96_n651);
   mult_28_C96_U1319 : NAN2D1 port map( A1 => mult_28_C96_n909, A2 => 
                           mult_28_C96_n401, Z => mult_28_C96_n196);
   mult_28_C96_U1318 : AOI21DL port map( A1 => mult_28_C96_n1020, A2 => 
                           mult_28_C96_n152, B => mult_28_C96_n153, Z => 
                           mult_28_C96_n151);
   mult_28_C96_U1317 : AOI21DL port map( A1 => mult_28_C96_n128, A2 => 
                           mult_28_C96_n1020, B => mult_28_C96_n129, Z => 
                           mult_28_C96_n127);
   mult_28_C96_U1316 : NAN2D1 port map( A1 => mult_28_C96_n1065, A2 => 
                           mult_28_C96_n375, Z => mult_28_C96_n180);
   mult_28_C96_U1315 : NAN2DL port map( A1 => mult_28_C96_n378, A2 => 
                           mult_28_C96_n380, Z => mult_28_C96_n1094);
   mult_28_C96_U1314 : NAN2DL port map( A1 => mult_28_C96_n389, A2 => 
                           mult_28_C96_n378, Z => mult_28_C96_n1093);
   mult_28_C96_U1313 : INVDL port map( A => mult_28_C96_n1066, Z => 
                           mult_28_C96_n199);
   mult_28_C96_U1312 : EXNOR2DL port map( A1 => mult_28_C96_n1059, A2 => 
                           coeff_memory_11_port, Z => mult_28_C96_n684);
   mult_28_C96_U1311 : EXNOR2DL port map( A1 => coeff_memory_13_port, A2 => 
                           mult_28_C96_n1059, Z => mult_28_C96_n667);
   mult_28_C96_U1310 : EXNOR2DL port map( A1 => mult_28_C96_n1059, A2 => 
                           coeff_memory_15_port, Z => mult_28_C96_n650);
   mult_28_C96_U1309 : EXNOR2DL port map( A1 => n42, A2 => coeff_memory_13_port
                           , Z => mult_28_C96_n671);
   mult_28_C96_U1308 : EXNOR2DL port map( A1 => n42, A2 => coeff_memory_15_port
                           , Z => mult_28_C96_n654);
   mult_28_C96_U1307 : OAI22M10D1 port map( A1 => coeff_memory_0_port, A2 => 
                           mult_28_C96_n769, B1 => mult_28_C96_n770, B2 => 
                           mult_28_C96_n6, Z => mult_28_C96_n635);
   mult_28_C96_U1306 : EXNOR2DL port map( A1 => y_15_port, A2 => 
                           coeff_memory_15_port, Z => mult_28_C96_n649);
   mult_28_C96_U1305 : OAI21DL port map( A1 => mult_28_C96_n934, A2 => 
                           mult_28_C96_n97, B => mult_28_C96_n100, Z => 
                           mult_28_C96_n96);
   mult_28_C96_U1304 : OAI21DL port map( A1 => mult_28_C96_n52, A2 => 
                           mult_28_C96_n1081, B => mult_28_C96_n1080, Z => 
                           mult_28_C96_n87);
   mult_28_C96_U1303 : EXNOR2DL port map( A1 => n33, A2 => coeff_memory_15_port
                           , Z => mult_28_C96_n659);
   mult_28_C96_U1302 : EXNOR2DL port map( A1 => n33, A2 => coeff_memory_3_port,
                           Z => mult_28_C96_n761);
   mult_28_C96_U1301 : EXNOR2DL port map( A1 => n33, A2 => coeff_memory_1_port,
                           Z => mult_28_C96_n778);
   mult_28_C96_U1300 : OAI22D1 port map( A1 => mult_28_C96_n771, A2 => 
                           mult_28_C96_n6, B1 => mult_28_C96_n770, B2 => 
                           mult_28_C96_n824, Z => mult_28_C96_n636);
   mult_28_C96_U1299 : INVDL port map( A => mult_28_C96_n954, Z => 
                           mult_28_C96_n192);
   mult_28_C96_U1298 : INVD1 port map( A => mult_28_C96_n212, Z => 
                           mult_28_C96_n211);
   mult_28_C96_U1297 : OAI21DL port map( A1 => mult_28_C96_n192, A2 => 
                           mult_28_C96_n914, B => mult_28_C96_n187, Z => 
                           mult_28_C96_n183);
   mult_28_C96_U1296 : EXNOR2DL port map( A1 => n34, A2 => coeff_memory_9_port,
                           Z => mult_28_C96_n714);
   mult_28_C96_U1295 : EXNOR2DL port map( A1 => n34, A2 => coeff_memory_7_port,
                           Z => mult_28_C96_n731);
   mult_28_C96_U1294 : EXNOR2DL port map( A1 => n34, A2 => coeff_memory_5_port,
                           Z => mult_28_C96_n748);
   mult_28_C96_U1293 : EXNOR2DL port map( A1 => n34, A2 => coeff_memory_3_port,
                           Z => mult_28_C96_n765);
   mult_28_C96_U1292 : EXNOR2DL port map( A1 => n34, A2 => coeff_memory_1_port,
                           Z => mult_28_C96_n782);
   mult_28_C96_U1291 : INVD1 port map( A => coeff_memory_1_port, Z => 
                           mult_28_C96_n832);
   mult_28_C96_U1290 : INVD1 port map( A => coeff_memory_0_port, Z => 
                           mult_28_C96_n824);
   mult_28_C96_U1289 : NAN2D1 port map( A1 => mult_28_C96_n808, A2 => 
                           mult_28_C96_n824, Z => mult_28_C96_n6);
   mult_28_C96_U1288 : NAN2D1 port map( A1 => mult_28_C96_n806, A2 => 
                           mult_28_C96_n16, Z => mult_28_C96_n18);
   mult_28_C96_U1287 : EXNOR2D1 port map( A1 => coeff_memory_3_port, A2 => 
                           coeff_memory_4_port, Z => mult_28_C96_n16);
   mult_28_C96_U1286 : NAN2D1 port map( A1 => mult_28_C96_n807, A2 => 
                           mult_28_C96_n9, Z => mult_28_C96_n12);
   mult_28_C96_U1285 : EXNOR2D1 port map( A1 => coeff_memory_1_port, A2 => 
                           coeff_memory_2_port, Z => mult_28_C96_n9);
   mult_28_C96_U1284 : NAN2D1 port map( A1 => mult_28_C96_n805, A2 => 
                           mult_28_C96_n22, Z => mult_28_C96_n24);
   mult_28_C96_U1283 : EXNOR2D1 port map( A1 => coeff_memory_5_port, A2 => 
                           coeff_memory_6_port, Z => mult_28_C96_n22);
   mult_28_C96_U1282 : NAN2D1 port map( A1 => mult_28_C96_n804, A2 => 
                           mult_28_C96_n28, Z => mult_28_C96_n30);
   mult_28_C96_U1281 : EXNOR2D1 port map( A1 => coeff_memory_7_port, A2 => 
                           coeff_memory_8_port, Z => mult_28_C96_n28);
   mult_28_C96_U1280 : NAN2D1 port map( A1 => mult_28_C96_n803, A2 => 
                           mult_28_C96_n34, Z => mult_28_C96_n36);
   mult_28_C96_U1279 : EXNOR2D1 port map( A1 => coeff_memory_9_port, A2 => 
                           coeff_memory_10_port, Z => mult_28_C96_n34);
   mult_28_C96_U1278 : NAN2D1 port map( A1 => mult_28_C96_n802, A2 => 
                           mult_28_C96_n40, Z => mult_28_C96_n42);
   mult_28_C96_U1277 : EXNOR2D1 port map( A1 => coeff_memory_11_port, A2 => 
                           coeff_memory_12_port, Z => mult_28_C96_n40);
   mult_28_C96_U1276 : NAN2D1 port map( A1 => mult_28_C96_n801, A2 => 
                           mult_28_C96_n46, Z => mult_28_C96_n48);
   mult_28_C96_U1275 : EXNOR2D1 port map( A1 => coeff_memory_13_port, A2 => 
                           coeff_memory_14_port, Z => mult_28_C96_n46);
   mult_28_C96_U1274 : INVD1 port map( A => coeff_memory_3_port, Z => 
                           mult_28_C96_n831);
   mult_28_C96_U1273 : ADHALFDL port map( A => mult_28_C96_n631, B => 
                           mult_28_C96_n519, CO => mult_28_C96_n511, S => 
                           mult_28_C96_n512);
   mult_28_C96_U1272 : INVD1 port map( A => coeff_memory_5_port, Z => 
                           mult_28_C96_n830);
   mult_28_C96_U1271 : INVD1 port map( A => coeff_memory_7_port, Z => 
                           mult_28_C96_n829);
   mult_28_C96_U1270 : INVD1 port map( A => coeff_memory_9_port, Z => 
                           mult_28_C96_n828);
   mult_28_C96_U1269 : INVD1 port map( A => coeff_memory_11_port, Z => 
                           mult_28_C96_n827);
   mult_28_C96_U1268 : INVD1 port map( A => coeff_memory_15_port, Z => 
                           mult_28_C96_n825);
   mult_28_C96_U1267 : INVD1 port map( A => coeff_memory_13_port, Z => 
                           mult_28_C96_n826);
   mult_28_C96_U1266 : OR2D1 port map( A1 => mult_28_C96_n305, A2 => 
                           mult_28_C96_n1092, Z => mult_28_C96_n1091);
   mult_28_C96_U1265 : AO21D1 port map( A1 => mult_28_C96_n42, A2 => 
                           mult_28_C96_n40, B => mult_28_C96_n666, Z => 
                           mult_28_C96_n532);
   mult_28_C96_U1264 : INVD2 port map( A => mult_28_C96_n309, Z => 
                           mult_28_C96_n310);
   mult_28_C96_U1263 : AND2D1 port map( A1 => mult_28_C96_n648, A2 => 
                           mult_28_C96_n520, Z => mult_28_C96_n1090);
   mult_28_C96_U1262 : NOR2DL port map( A1 => mult_28_C96_n646, A2 => 
                           mult_28_C96_n512, Z => mult_28_C96_n265);
   mult_28_C96_U1261 : NAN2DL port map( A1 => mult_28_C96_n646, A2 => 
                           mult_28_C96_n512, Z => mult_28_C96_n266);
   mult_28_C96_U1260 : AO21D1 port map( A1 => mult_28_C96_n36, A2 => 
                           mult_28_C96_n34, B => mult_28_C96_n683, Z => 
                           mult_28_C96_n548);
   mult_28_C96_U1259 : NAN2DL port map( A1 => mult_28_C96_n305, A2 => 
                           mult_28_C96_n1092, Z => mult_28_C96_n84);
   mult_28_C96_U1258 : NAN2D1 port map( A1 => mult_28_C96_n1091, A2 => 
                           mult_28_C96_n84, Z => mult_28_C96_n54);
   mult_28_C96_U1257 : INVD2 port map( A => mult_28_C96_n333, Z => 
                           mult_28_C96_n334);
   mult_28_C96_U1256 : INVD2 port map( A => mult_28_C96_n351, Z => 
                           mult_28_C96_n352);
   mult_28_C96_U1255 : INVD2 port map( A => mult_28_C96_n373, Z => 
                           mult_28_C96_n374);
   mult_28_C96_U1254 : AO21D1 port map( A1 => mult_28_C96_n18, A2 => 
                           mult_28_C96_n16, B => mult_28_C96_n734, Z => 
                           mult_28_C96_n599);
   mult_28_C96_U1253 : AO21D1 port map( A1 => mult_28_C96_n6, A2 => 
                           mult_28_C96_n824, B => mult_28_C96_n768, Z => 
                           mult_28_C96_n633);
   mult_28_C96_U1252 : NAN2DL port map( A1 => mult_28_C96_n307, A2 => 
                           mult_28_C96_n306, Z => mult_28_C96_n93);
   mult_28_C96_U1251 : NAN2DL port map( A1 => mult_28_C96_n311, A2 => 
                           mult_28_C96_n308, Z => mult_28_C96_n104);
   mult_28_C96_U1250 : NAN2D1 port map( A1 => mult_28_C96_n312, A2 => 
                           mult_28_C96_n315, Z => mult_28_C96_n113);
   mult_28_C96_U1249 : AND2D1 port map( A1 => mult_28_C96_n647, A2 => 
                           mult_28_C96_n632, Z => mult_28_C96_n1089);
   mult_28_C96_U1248 : OR2D1 port map( A1 => mult_28_C96_n647, A2 => 
                           mult_28_C96_n632, Z => mult_28_C96_n1088);
   mult_28_C96_U1247 : AND2D1 port map( A1 => mult_28_C96_n510, A2 => 
                           mult_28_C96_n645, Z => mult_28_C96_n1087);
   mult_28_C96_U1246 : NAN2DL port map( A1 => mult_28_C96_n506, A2 => 
                           mult_28_C96_n509, Z => mult_28_C96_n258);
   mult_28_C96_U1245 : OR2D1 port map( A1 => mult_28_C96_n502, A2 => 
                           mult_28_C96_n505, Z => mult_28_C96_n1084);
   mult_28_C96_U1244 : NOR2DL port map( A1 => mult_28_C96_n496, A2 => 
                           mult_28_C96_n501, Z => mult_28_C96_n249);
   mult_28_C96_U1243 : NAN2DL port map( A1 => mult_28_C96_n496, A2 => 
                           mult_28_C96_n501, Z => mult_28_C96_n250);
   mult_28_C96_U1242 : AND2D1 port map( A1 => mult_28_C96_n490, A2 => 
                           mult_28_C96_n495, Z => mult_28_C96_n1083);
   mult_28_C96_U1241 : NAN2D1 port map( A1 => mult_28_C96_n430, A2 => 
                           mult_28_C96_n441, Z => mult_28_C96_n210);
   mult_28_C96_U1240 : EXNOR2D1 port map( A1 => mult_28_C96_n380, A2 => 
                           mult_28_C96_n389, Z => mult_28_C96_n1082);
   mult_28_C96_U1239 : NOR2D1 port map( A1 => mult_28_C96_n112, A2 => 
                           mult_28_C96_n103, Z => mult_28_C96_n101);
   mult_28_C96_U1238 : OR2D1 port map( A1 => mult_28_C96_n97, A2 => 
                           mult_28_C96_n92, Z => mult_28_C96_n1081);
   mult_28_C96_U1237 : NAN2D1 port map( A1 => mult_28_C96_n316, A2 => 
                           mult_28_C96_n321, Z => mult_28_C96_n118);
   mult_28_C96_U1236 : OA21DL port map( A1 => mult_28_C96_n100, A2 => 
                           mult_28_C96_n92, B => mult_28_C96_n93, Z => 
                           mult_28_C96_n1080);
   mult_28_C96_U1235 : AND2D1 port map( A1 => mult_28_C96_n464, A2 => 
                           mult_28_C96_n473, Z => mult_28_C96_n1079);
   mult_28_C96_U1234 : NAN2D1 port map( A1 => mult_28_C96_n336, A2 => 
                           mult_28_C96_n343, Z => mult_28_C96_n155);
   mult_28_C96_U1233 : NAN2D1 port map( A1 => mult_28_C96_n344, A2 => 
                           mult_28_C96_n353, Z => mult_28_C96_n168);
   mult_28_C96_U1232 : NAN2D1 port map( A1 => mult_28_C96_n328, A2 => 
                           mult_28_C96_n335, Z => mult_28_C96_n150);
   mult_28_C96_U1231 : INVD2 port map( A => mult_28_C96_n149, Z => 
                           mult_28_C96_n281);
   mult_28_C96_U1230 : OA21M20D1 port map( A1 => mult_28_C96_n960, A2 => 
                           mult_28_C96_n278, B => mult_28_C96_n113, Z => 
                           mult_28_C96_n109);
   mult_28_C96_U1229 : NOR2D1 port map( A1 => mult_28_C96_n53, A2 => 
                           mult_28_C96_n117, Z => mult_28_C96_n115);
   mult_28_C96_U1228 : NAN2D1 port map( A1 => mult_28_C96_n279, A2 => 
                           mult_28_C96_n278, Z => mult_28_C96_n108);
   mult_28_C96_U1227 : NOR2DL port map( A1 => mult_28_C96_n53, A2 => 
                           mult_28_C96_n1081, Z => mult_28_C96_n86);
   mult_28_C96_U1226 : INVDL port map( A => mult_28_C96_n154, Z => 
                           mult_28_C96_n282);
   mult_28_C96_U1225 : NAN2D1 port map( A1 => mult_28_C96_n282, A2 => 
                           mult_28_C96_n281, Z => mult_28_C96_n143);
   mult_28_C96_U1224 : NOR2M1DL port map( A1 => mult_28_C96_n912, A2 => 
                           mult_28_C96_n914, Z => mult_28_C96_n182);
   mult_28_C96_U1223 : INVDL port map( A => mult_28_C96_n200, Z => 
                           mult_28_C96_n288);
   mult_28_C96_U1222 : NAN2DL port map( A1 => mult_28_C96_n284, A2 => 
                           mult_28_C96_n173, Z => mult_28_C96_n63);
   mult_28_C96_U1221 : NOR2D1 port map( A1 => mult_28_C96_n163, A2 => 
                           mult_28_C96_n143, Z => mult_28_C96_n141);
   mult_28_C96_U1220 : AND2DL port map( A1 => mult_28_C96_n285, A2 => 
                           mult_28_C96_n180, Z => mult_28_C96_n1076);
   mult_28_C96_U1219 : AND2D1 port map( A1 => mult_28_C96_n279, A2 => 
                           mult_28_C96_n118, Z => mult_28_C96_n1075);
   mult_28_C96_U1218 : OA21M20D1 port map( A1 => mult_28_C96_n148, A2 => 
                           mult_28_C96_n1078, B => mult_28_C96_n139, Z => 
                           mult_28_C96_n135);
   mult_28_C96_U1217 : NOR2D1 port map( A1 => mult_28_C96_n200, A2 => 
                           mult_28_C96_n913, Z => mult_28_C96_n189);
   mult_28_C96_U1216 : INVDL port map( A => mult_28_C96_n184, Z => 
                           mult_28_C96_n286);
   mult_28_C96_U1215 : NOR2DL port map( A1 => mult_28_C96_n53, A2 => 
                           mult_28_C96_n97, Z => mult_28_C96_n95);
   mult_28_C96_U1214 : OA22DL port map( A1 => mult_28_C96_n650, A2 => 
                           mult_28_C96_n48, B1 => mult_28_C96_n649, B2 => 
                           mult_28_C96_n46, Z => mult_28_C96_n1092);
   mult_28_C96_U1213 : OAI22DL port map( A1 => mult_28_C96_n652, A2 => 
                           mult_28_C96_n48, B1 => mult_28_C96_n651, B2 => 
                           mult_28_C96_n46, Z => mult_28_C96_n523);
   mult_28_C96_U1212 : OAI22DL port map( A1 => mult_28_C96_n653, A2 => 
                           mult_28_C96_n48, B1 => mult_28_C96_n652, B2 => 
                           mult_28_C96_n46, Z => mult_28_C96_n524);
   mult_28_C96_U1211 : OAI22DL port map( A1 => mult_28_C96_n684, A2 => 
                           mult_28_C96_n36, B1 => mult_28_C96_n683, B2 => 
                           mult_28_C96_n34, Z => mult_28_C96_n549);
   mult_28_C96_U1210 : OAI22DL port map( A1 => mult_28_C96_n688, A2 => 
                           mult_28_C96_n36, B1 => mult_28_C96_n687, B2 => 
                           mult_28_C96_n34, Z => mult_28_C96_n553);
   mult_28_C96_U1209 : AND2DL port map( A1 => mult_28_C96_n502, A2 => 
                           mult_28_C96_n505, Z => mult_28_C96_n1085);
   mult_28_C96_U1208 : OR2D1 port map( A1 => mult_28_C96_n490, A2 => 
                           mult_28_C96_n495, Z => mult_28_C96_n1071);
   mult_28_C96_U1207 : NAN2DL port map( A1 => mult_28_C96_n416, A2 => 
                           mult_28_C96_n429, Z => mult_28_C96_n207);
   mult_28_C96_U1206 : INVD1 port map( A => mult_28_C96_n112, Z => 
                           mult_28_C96_n278);
   mult_28_C96_U1205 : NAN2DL port map( A1 => mult_28_C96_n322, A2 => 
                           mult_28_C96_n327, Z => mult_28_C96_n139);
   mult_28_C96_U1204 : NAN2DL port map( A1 => mult_28_C96_n276, A2 => 
                           mult_28_C96_n93, Z => mult_28_C96_n1070);
   mult_28_C96_U1203 : AOI21DL port map( A1 => mult_28_C96_n1019, A2 => 
                           mult_28_C96_n95, B => mult_28_C96_n96, Z => 
                           mult_28_C96_n1069);
   mult_28_C96_U1202 : EXOR2D1 port map( A1 => mult_28_C96_n1069, A2 => 
                           mult_28_C96_n1070, Z => m5_14);
   mult_28_C96_U1201 : OAI21D1 port map( A1 => mult_28_C96_n1068, A2 => 
                           mult_28_C96_n243, B => mult_28_C96_n232, Z => 
                           mult_28_C96_n230);
   mult_28_C96_U1200 : NAN2M1DL port map( A1 => mult_28_C96_n206, A2 => 
                           mult_28_C96_n207, Z => mult_28_C96_n68);
   mult_28_C96_U1199 : NAN2M1DL port map( A1 => mult_28_C96_n103, A2 => 
                           mult_28_C96_n104, Z => mult_28_C96_n56);
   mult_28_C96_U1198 : NAN2DL port map( A1 => mult_28_C96_n278, A2 => 
                           mult_28_C96_n113, Z => mult_28_C96_n57);
   mult_28_C96_U1197 : INVD2 port map( A => mult_28_C96_n117, Z => 
                           mult_28_C96_n279);
   mult_28_C96_U1196 : NAN2D2 port map( A1 => mult_28_C96_n281, A2 => 
                           mult_28_C96_n1078, Z => mult_28_C96_n134);
   mult_28_C96_U1195 : INVDL port map( A => mult_28_C96_n1028, Z => 
                           mult_28_C96_n284);
   mult_28_C96_U1194 : AOI21M10DL port map( A1 => mult_28_C96_n155, A2 => 
                           mult_28_C96_n281, B => mult_28_C96_n148, Z => 
                           mult_28_C96_n144);
   mult_28_C96_U1193 : NAN2M1DL port map( A1 => mult_28_C96_n913, A2 => 
                           mult_28_C96_n196, Z => mult_28_C96_n66);
   mult_28_C96_U1192 : AOI21DL port map( A1 => mult_28_C96_n182, A2 => 
                           mult_28_C96_n202, B => mult_28_C96_n183, Z => 
                           mult_28_C96_n1067);
   mult_28_C96_U1191 : EXNOR2D1 port map( A1 => mult_28_C96_n1067, A2 => 
                           mult_28_C96_n1076, Z => m5_5);
   mult_28_C96_U1190 : EXNOR2D2 port map( A1 => mult_28_C96_n160, A2 => 
                           mult_28_C96_n1074, Z => m5_8);
   mult_28_C96_U1189 : AND2DL port map( A1 => mult_28_C96_n282, A2 => 
                           mult_28_C96_n155, Z => mult_28_C96_n1074);
   mult_28_C96_U1188 : EXNOR2D2 port map( A1 => mult_28_C96_n151, A2 => 
                           mult_28_C96_n1073, Z => m5_9);
   mult_28_C96_U1187 : AND2DL port map( A1 => mult_28_C96_n281, A2 => 
                           mult_28_C96_n150, Z => mult_28_C96_n1073);
   mult_28_C96_U1186 : INVDL port map( A => mult_28_C96_n319, Z => 
                           mult_28_C96_n320);
   mult_28_C96_U1185 : OR2D1 port map( A1 => mult_28_C96_n510, A2 => 
                           mult_28_C96_n645, Z => mult_28_C96_n1086);
   mult_28_C96_U1184 : NOR2D1 port map( A1 => mult_28_C96_n506, A2 => 
                           mult_28_C96_n509, Z => mult_28_C96_n257);
   mult_28_C96_U1183 : AND2D1 port map( A1 => mult_28_C96_n482, A2 => 
                           mult_28_C96_n489, Z => mult_28_C96_n1072);
   mult_28_C96_U1182 : AOI21DL port map( A1 => mult_28_C96_n106, A2 => 
                           mult_28_C96_n1020, B => mult_28_C96_n107, Z => 
                           mult_28_C96_n105);
   mult_28_C96_U1181 : NAN2DL port map( A1 => mult_28_C96_n101, A2 => 
                           mult_28_C96_n279, Z => mult_28_C96_n97);
   mult_28_C96_U1180 : NOR2D1 port map( A1 => mult_28_C96_n1028, A2 => 
                           mult_28_C96_n167, Z => mult_28_C96_n161);
   mult_28_C96_U1179 : NOR2DL port map( A1 => mult_28_C96_n53, A2 => 
                           mult_28_C96_n108, Z => mult_28_C96_n106);
   mult_28_C96_U1178 : EXNOR2D2 port map( A1 => y_12_port, A2 => 
                           coeff_memory_5_port, Z => mult_28_C96_n737);
   mult_28_C96_U1177 : OAI22D1 port map( A1 => mult_28_C96_n947, A2 => 
                           mult_28_C96_n18, B1 => mult_28_C96_n737, B2 => 
                           mult_28_C96_n16, Z => mult_28_C96_n603);
   mult_28_C96_U1176 : EXNOR2D2 port map( A1 => y_14_port, A2 => 
                           coeff_memory_1_port, Z => mult_28_C96_n769);
   mult_28_C96_U1175 : NOR2D2 port map( A1 => mult_28_C96_n416, A2 => 
                           mult_28_C96_n429, Z => mult_28_C96_n206);
   mult_28_C96_U1174 : EXNOR2D2 port map( A1 => n33, A2 => coeff_memory_9_port,
                           Z => mult_28_C96_n710);
   mult_28_C96_U1173 : EXNOR2D2 port map( A1 => y_6_port, A2 => 
                           coeff_memory_11_port, Z => mult_28_C96_n692);
   mult_28_C96_U1172 : EXNOR2D2 port map( A1 => n33, A2 => coeff_memory_11_port
                           , Z => mult_28_C96_n693);
   mult_28_C96_U1171 : NAN2D1 port map( A1 => mult_28_C96_n402, A2 => 
                           mult_28_C96_n415, Z => mult_28_C96_n201);
   mult_28_C96_U1170 : EXNOR2DL port map( A1 => y_6_port, A2 => 
                           coeff_memory_1_port, Z => mult_28_C96_n777);
   mult_28_C96_U1169 : EXNOR2DL port map( A1 => y_6_port, A2 => 
                           coeff_memory_5_port, Z => mult_28_C96_n743);
   mult_28_C96_U1168 : EXNOR2DL port map( A1 => y_6_port, A2 => 
                           coeff_memory_3_port, Z => mult_28_C96_n760);
   mult_28_C96_U1167 : EXOR3DL port map( A1 => mult_28_C96_n381, A2 => 
                           mult_28_C96_n370, A3 => mult_28_C96_n1058, Z => 
                           mult_28_C96_n1064);
   mult_28_C96_U1166 : NAN3D2 port map( A1 => mult_28_C96_n1062, A2 => 
                           mult_28_C96_n1063, A3 => mult_28_C96_n1061, Z => 
                           mult_28_C96_n421);
   mult_28_C96_U1165 : NAN2D1 port map( A1 => mult_28_C96_n1053, A2 => 
                           mult_28_C96_n426, Z => mult_28_C96_n1063);
   mult_28_C96_U1164 : NAN2D1 port map( A1 => mult_28_C96_n1053, A2 => 
                           mult_28_C96_n901, Z => mult_28_C96_n1062);
   mult_28_C96_U1163 : NAN2D1 port map( A1 => mult_28_C96_n426, A2 => 
                           mult_28_C96_n901, Z => mult_28_C96_n1061);
   mult_28_C96_U1162 : EXNOR2DL port map( A1 => y_9_port, A2 => 
                           coeff_memory_1_port, Z => mult_28_C96_n774);
   mult_28_C96_U1161 : EXNOR2DL port map( A1 => y_9_port, A2 => 
                           coeff_memory_15_port, Z => mult_28_C96_n655);
   mult_28_C96_U1160 : BUFDL port map( A => mult_28_C96_n379, Z => 
                           mult_28_C96_n1058);
   mult_28_C96_U1159 : INVDL port map( A => mult_28_C96_n192, Z => 
                           mult_28_C96_n1057);
   mult_28_C96_U1158 : EXNOR2D2 port map( A1 => mult_28_C96_n127, A2 => 
                           mult_28_C96_n1075, Z => m5_11);
   mult_28_C96_U1157 : EXNOR2D2 port map( A1 => n42, A2 => coeff_memory_7_port,
                           Z => mult_28_C96_n722);
   mult_28_C96_U1156 : INVDL port map( A => mult_28_C96_n910, Z => 
                           mult_28_C96_n285);
   mult_28_C96_U1155 : EXNOR2D2 port map( A1 => mult_28_C96_n1082, A2 => 
                           mult_28_C96_n378, Z => mult_28_C96_n376);
   mult_28_C96_U1154 : OR2D2 port map( A1 => mult_28_C96_n529, A2 => 
                           mult_28_C96_n427, Z => mult_28_C96_n413);
   mult_28_C96_U1153 : EXNOR2D2 port map( A1 => n43, A2 => coeff_memory_15_port
                           , Z => mult_28_C96_n662);
   mult_28_C96_U1152 : EXNOR2D2 port map( A1 => n33, A2 => coeff_memory_13_port
                           , Z => mult_28_C96_n676);
   mult_28_C96_U1151 : EXNOR2DL port map( A1 => mult_28_C96_n1020, A2 => 
                           mult_28_C96_n63, Z => m5_6);
   mult_28_C96_U1150 : AOI21DL port map( A1 => mult_28_C96_n1019, A2 => 
                           mult_28_C96_n86, B => mult_28_C96_n87, Z => 
                           mult_28_C96_n85);
   mult_28_C96_U1149 : AO21D1 port map( A1 => mult_28_C96_n12, A2 => 
                           mult_28_C96_n9, B => mult_28_C96_n751, Z => 
                           mult_28_C96_n616);
   mult_28_C96_U1148 : NAN3D2 port map( A1 => mult_28_C96_n1054, A2 => 
                           mult_28_C96_n1055, A3 => mult_28_C96_n1056, Z => 
                           mult_28_C96_n379);
   mult_28_C96_U1147 : NAN2D1 port map( A1 => mult_28_C96_n395, A2 => 
                           mult_28_C96_n616, Z => mult_28_C96_n1056);
   mult_28_C96_U1146 : NAN2D1 port map( A1 => mult_28_C96_n393, A2 => 
                           mult_28_C96_n395, Z => mult_28_C96_n1054);
   mult_28_C96_U1145 : EXNOR2D2 port map( A1 => y_7_port, A2 => 
                           coeff_memory_7_port, Z => mult_28_C96_n725);
   mult_28_C96_U1144 : EXNOR2DL port map( A1 => y_7_port, A2 => 
                           coeff_memory_13_port, Z => mult_28_C96_n674);
   mult_28_C96_U1143 : EXNOR2DL port map( A1 => y_7_port, A2 => 
                           coeff_memory_15_port, Z => mult_28_C96_n657);
   mult_28_C96_U1142 : EXNOR2DL port map( A1 => mult_28_C96_n1042, A2 => 
                           coeff_memory_1_port, Z => mult_28_C96_n776);
   mult_28_C96_U1141 : NOR2D2 port map( A1 => mult_28_C96_n179, A2 => 
                           mult_28_C96_n184, Z => mult_28_C96_n177);
   mult_28_C96_U1140 : ADFULD1 port map( A => mult_28_C96_n544, B => 
                           mult_28_C96_n428, CI => mult_28_C96_n559, CO => 
                           mult_28_C96_n425, S => mult_28_C96_n426);
   mult_28_C96_U1139 : EXNOR2D2 port map( A1 => y_15_port, A2 => 
                           coeff_memory_1_port, Z => mult_28_C96_n768);
   mult_28_C96_U1138 : OAI22D1 port map( A1 => mult_28_C96_n769, A2 => 
                           mult_28_C96_n6, B1 => mult_28_C96_n768, B2 => 
                           mult_28_C96_n824, Z => mult_28_C96_n1053);
   mult_28_C96_U1137 : EXOR3DL port map( A1 => mult_28_C96_n417, A2 => 
                           mult_28_C96_n966, A3 => mult_28_C96_n404, Z => 
                           mult_28_C96_n1052);
   mult_28_C96_U1136 : EXNOR2DL port map( A1 => y_8_port, A2 => 
                           coeff_memory_3_port, Z => mult_28_C96_n758);
   mult_28_C96_U1135 : EXNOR2DL port map( A1 => coeff_memory_1_port, A2 => 
                           y_8_port, Z => mult_28_C96_n775);
   mult_28_C96_U1134 : EXNOR2DL port map( A1 => y_8_port, A2 => 
                           coeff_memory_13_port, Z => mult_28_C96_n673);
   mult_28_C96_U1133 : AND2DL port map( A1 => mult_28_C96_n283, A2 => 
                           mult_28_C96_n168, Z => mult_28_C96_n1049);
   mult_28_C96_U1132 : EXNOR2D2 port map( A1 => mult_28_C96_n169, A2 => 
                           mult_28_C96_n1049, Z => m5_7);
   mult_28_C96_U1131 : AOI21D1 port map( A1 => mult_28_C96_n115, A2 => 
                           mult_28_C96_n1020, B => mult_28_C96_n116, Z => 
                           mult_28_C96_n114);
   mult_28_C96_U1130 : EXOR2D4 port map( A1 => mult_28_C96_n211, A2 => 
                           mult_28_C96_n69, Z => m5_0);
   mult_28_C96_U1129 : OAI22D2 port map( A1 => mult_28_C96_n752, A2 => 
                           mult_28_C96_n12, B1 => mult_28_C96_n751, B2 => 
                           mult_28_C96_n9, Z => mult_28_C96_n617);
   mult_28_C96_U1128 : NAN2D1 port map( A1 => mult_28_C96_n573, A2 => 
                           mult_28_C96_n425, Z => mult_28_C96_n1048);
   mult_28_C96_U1127 : NAN3D2 port map( A1 => mult_28_C96_n1043, A2 => 
                           mult_28_C96_n1045, A3 => mult_28_C96_n1044, Z => 
                           mult_28_C96_n391);
   mult_28_C96_U1126 : NAN2D1 port map( A1 => mult_28_C96_n396, A2 => 
                           mult_28_C96_n617, Z => mult_28_C96_n1045);
   mult_28_C96_U1125 : NAN2D1 port map( A1 => mult_28_C96_n409, A2 => 
                           mult_28_C96_n617, Z => mult_28_C96_n1044);
   mult_28_C96_U1124 : NAN2D1 port map( A1 => mult_28_C96_n396, A2 => 
                           mult_28_C96_n409, Z => mult_28_C96_n1043);
   mult_28_C96_U1123 : EXOR2D4 port map( A1 => mult_28_C96_n188, A2 => 
                           mult_28_C96_n65, Z => m5_4);
   mult_28_C96_U1122 : EXOR2D2 port map( A1 => mult_28_C96_n114, A2 => 
                           mult_28_C96_n57, Z => m5_12);
   mult_28_C96_U1121 : EXNOR2DL port map( A1 => mult_28_C96_n932, A2 => 
                           coeff_memory_15_port, Z => mult_28_C96_n652);
   mult_28_C96_U1120 : EXNOR2DL port map( A1 => mult_28_C96_n932, A2 => 
                           coeff_memory_13_port, Z => mult_28_C96_n669);
   mult_28_C96_U1119 : EXNOR2DL port map( A1 => y_12_port, A2 => 
                           coeff_memory_11_port, Z => mult_28_C96_n686);
   mult_28_C96_U1118 : EXNOR2D2 port map( A1 => y_12_port, A2 => 
                           coeff_memory_7_port, Z => mult_28_C96_n720);
   mult_28_C96_U1117 : EXNOR2D2 port map( A1 => y_3_port, A2 => 
                           coeff_memory_11_port, Z => mult_28_C96_n695);
   mult_28_C96_U1116 : EXNOR2DL port map( A1 => y_7_port, A2 => 
                           coeff_memory_9_port, Z => mult_28_C96_n708);
   mult_28_C96_U1115 : NAN2DL port map( A1 => mult_28_C96_n633, A2 => 
                           mult_28_C96_n423, Z => mult_28_C96_n1039);
   mult_28_C96_U1114 : NAN3D2 port map( A1 => mult_28_C96_n1034, A2 => 
                           mult_28_C96_n1035, A3 => mult_28_C96_n1036, Z => 
                           mult_28_C96_n423);
   mult_28_C96_U1113 : NAN2D1 port map( A1 => mult_28_C96_n439, A2 => 
                           mult_28_C96_n589, Z => mult_28_C96_n1036);
   mult_28_C96_U1112 : NAN2D1 port map( A1 => mult_28_C96_n574, A2 => 
                           mult_28_C96_n589, Z => mult_28_C96_n1035);
   mult_28_C96_U1111 : EXOR3D2 port map( A1 => mult_28_C96_n574, A2 => 
                           mult_28_C96_n439, A3 => mult_28_C96_n589, Z => 
                           mult_28_C96_n424);
   mult_28_C96_U1110 : OAI21D1 port map( A1 => mult_28_C96_n211, A2 => 
                           mult_28_C96_n209, B => mult_28_C96_n210, Z => 
                           mult_28_C96_n208);
   mult_28_C96_U1109 : INVDL port map( A => mult_28_C96_n164, Z => 
                           mult_28_C96_n1033);
   mult_28_C96_U1108 : OAI22DL port map( A1 => mult_28_C96_n674, A2 => 
                           mult_28_C96_n42, B1 => mult_28_C96_n673, B2 => 
                           mult_28_C96_n40, Z => mult_28_C96_n539);
   mult_28_C96_U1107 : NAN3D1 port map( A1 => mult_28_C96_n1030, A2 => 
                           mult_28_C96_n1032, A3 => mult_28_C96_n1031, Z => 
                           mult_28_C96_n359);
   mult_28_C96_U1106 : NAN2DL port map( A1 => mult_28_C96_n569, A2 => 
                           mult_28_C96_n539, Z => mult_28_C96_n1032);
   mult_28_C96_U1105 : NAN2DL port map( A1 => mult_28_C96_n584, A2 => 
                           mult_28_C96_n539, Z => mult_28_C96_n1031);
   mult_28_C96_U1104 : NAN2DL port map( A1 => mult_28_C96_n584, A2 => 
                           mult_28_C96_n569, Z => mult_28_C96_n1030);
   mult_28_C96_U1103 : OAI22D2 port map( A1 => mult_28_C96_n6, A2 => 
                           mult_28_C96_n773, B1 => mult_28_C96_n772, B2 => 
                           mult_28_C96_n824, Z => mult_28_C96_n638);
   mult_28_C96_U1102 : NAN2D1 port map( A1 => mult_28_C96_n189, A2 => 
                           mult_28_C96_n177, Z => mult_28_C96_n175);
   mult_28_C96_U1101 : EXNOR2DL port map( A1 => y_9_port, A2 => 
                           coeff_memory_7_port, Z => mult_28_C96_n723);
   mult_28_C96_U1100 : BUFD1 port map( A => y_14_port, Z => mult_28_C96_n1059);
   mult_28_C96_U1099 : EXNOR2D2 port map( A1 => mult_28_C96_n1059, A2 => 
                           coeff_memory_9_port, Z => mult_28_C96_n701);
   mult_28_C96_U1098 : OAI22D1 port map( A1 => mult_28_C96_n769, A2 => 
                           mult_28_C96_n6, B1 => mult_28_C96_n768, B2 => 
                           mult_28_C96_n824, Z => mult_28_C96_n634);
   mult_28_C96_U1097 : INVD1 port map( A => mult_28_C96_n1041, Z => 
                           mult_28_C96_n1042);
   mult_28_C96_U1096 : EXNOR2D2 port map( A1 => mult_28_C96_n1042, A2 => 
                           coeff_memory_3_port, Z => mult_28_C96_n759);
   mult_28_C96_U1095 : NAN2DL port map( A1 => mult_28_C96_n453, A2 => 
                           mult_28_C96_n442, Z => mult_28_C96_n1027);
   mult_28_C96_U1094 : OAI21D1 port map( A1 => mult_28_C96_n210, A2 => 
                           mult_28_C96_n206, B => mult_28_C96_n207, Z => 
                           mult_28_C96_n205);
   mult_28_C96_U1093 : NAN2D1 port map( A1 => mult_28_C96_n408, A2 => 
                           mult_28_C96_n410, Z => mult_28_C96_n1026);
   mult_28_C96_U1092 : NAN2DL port map( A1 => mult_28_C96_n419, A2 => 
                           mult_28_C96_n410, Z => mult_28_C96_n1025);
   mult_28_C96_U1091 : NAN3D1 port map( A1 => mult_28_C96_n1021, A2 => 
                           mult_28_C96_n1023, A3 => mult_28_C96_n1022, Z => 
                           mult_28_C96_n387);
   mult_28_C96_U1090 : NAN2DL port map( A1 => mult_28_C96_n392, A2 => 
                           mult_28_C96_n390, Z => mult_28_C96_n1023);
   mult_28_C96_U1089 : NAN2DL port map( A1 => mult_28_C96_n403, A2 => 
                           mult_28_C96_n392, Z => mult_28_C96_n1022);
   mult_28_C96_U1088 : NAN2DL port map( A1 => mult_28_C96_n403, A2 => 
                           mult_28_C96_n390, Z => mult_28_C96_n1021);
   mult_28_C96_U1087 : OR2D2 port map( A1 => mult_28_C96_n322, A2 => 
                           mult_28_C96_n327, Z => mult_28_C96_n1078);
   mult_28_C96_U1086 : OAI21D1 port map( A1 => mult_28_C96_n175, A2 => 
                           mult_28_C96_n203, B => mult_28_C96_n176, Z => 
                           mult_28_C96_n51);
   mult_28_C96_U1085 : EXNOR2D2 port map( A1 => mult_28_C96_n1059, A2 => 
                           coeff_memory_7_port, Z => mult_28_C96_n718);
   mult_28_C96_U1084 : BUFD4 port map( A => mult_28_C96_n51, Z => 
                           mult_28_C96_n1020);
   mult_28_C96_U1083 : EXNOR2D2 port map( A1 => y_12_port, A2 => 
                           coeff_memory_9_port, Z => mult_28_C96_n703);
   mult_28_C96_U1082 : INVDL port map( A => mult_28_C96_n1018, Z => 
                           mult_28_C96_n1019);
   mult_28_C96_U1081 : INVDL port map( A => mult_28_C96_n1020, Z => 
                           mult_28_C96_n1018);
   mult_28_C96_U1080 : EXOR2D4 port map( A1 => mult_28_C96_n197, A2 => 
                           mult_28_C96_n66, Z => m5_3);
   mult_28_C96_U1079 : NOR2D2 port map( A1 => mult_28_C96_n344, A2 => 
                           mult_28_C96_n353, Z => mult_28_C96_n167);
   mult_28_C96_U1078 : EXNOR2D2 port map( A1 => n42, A2 => coeff_memory_5_port,
                           Z => mult_28_C96_n1060);
   mult_28_C96_U1077 : NAN2DL port map( A1 => mult_28_C96_n286, A2 => 
                           mult_28_C96_n187, Z => mult_28_C96_n65);
   mult_28_C96_U1076 : ADHALFD2 port map( A => mult_28_C96_n546, B => 
                           mult_28_C96_n514, CO => mult_28_C96_n451, S => 
                           mult_28_C96_n452);
   mult_28_C96_U1075 : EXNOR2D2 port map( A1 => mult_28_C96_n105, A2 => 
                           mult_28_C96_n1017, Z => m5_13);
   mult_28_C96_U1074 : OAI22D1 port map( A1 => mult_28_C96_n742, A2 => 
                           mult_28_C96_n18, B1 => mult_28_C96_n741, B2 => 
                           mult_28_C96_n16, Z => mult_28_C96_n607);
   mult_28_C96_U1073 : NAN2DL port map( A1 => mult_28_C96_n607, A2 => 
                           mult_28_C96_n469, Z => mult_28_C96_n1016);
   mult_28_C96_U1072 : NAN2DL port map( A1 => mult_28_C96_n622, A2 => 
                           mult_28_C96_n469, Z => mult_28_C96_n1015);
   mult_28_C96_U1071 : NAN2DL port map( A1 => mult_28_C96_n622, A2 => 
                           mult_28_C96_n607, Z => mult_28_C96_n1014);
   mult_28_C96_U1070 : NOR2D1 port map( A1 => mult_28_C96_n1051, A2 => 
                           mult_28_C96_n415, Z => mult_28_C96_n200);
   mult_28_C96_U1069 : NAN2D1 port map( A1 => mult_28_C96_n1052, A2 => 
                           mult_28_C96_n415, Z => mult_28_C96_n1066);
   mult_28_C96_U1068 : NAN3D1 port map( A1 => mult_28_C96_n1010, A2 => 
                           mult_28_C96_n1012, A3 => mult_28_C96_n1011, Z => 
                           mult_28_C96_n415);
   mult_28_C96_U1067 : NAN2DL port map( A1 => mult_28_C96_n431, A2 => 
                           mult_28_C96_n420, Z => mult_28_C96_n1012);
   mult_28_C96_U1066 : NAN2D1 port map( A1 => mult_28_C96_n418, A2 => 
                           mult_28_C96_n420, Z => mult_28_C96_n1011);
   mult_28_C96_U1065 : NAN2DL port map( A1 => mult_28_C96_n418, A2 => 
                           mult_28_C96_n431, Z => mult_28_C96_n1010);
   mult_28_C96_U1064 : EXOR2D1 port map( A1 => mult_28_C96_n420, A2 => 
                           mult_28_C96_n431, Z => mult_28_C96_n1009);
   mult_28_C96_U1063 : OR2D2 port map( A1 => mult_28_C96_n474, A2 => 
                           mult_28_C96_n481, Z => mult_28_C96_n1077);
   mult_28_C96_U1062 : AOI21D1 port map( A1 => mult_28_C96_n1020, A2 => 
                           mult_28_C96_n952, B => mult_28_C96_n1033, Z => 
                           mult_28_C96_n160);
   mult_28_C96_U1061 : INVDL port map( A => mult_28_C96_n1007, Z => 
                           mult_28_C96_n1008);
   mult_28_C96_U1060 : INVDL port map( A => y_9_port, Z => mult_28_C96_n1007);
   mult_28_C96_U1059 : EXOR3D1 port map( A1 => mult_28_C96_n616, A2 => 
                           mult_28_C96_n393, A3 => mult_28_C96_n395, Z => 
                           mult_28_C96_n380);
   mult_28_C96_U1058 : EXOR3DL port map( A1 => mult_28_C96_n417, A2 => 
                           mult_28_C96_n406, A3 => mult_28_C96_n404, Z => 
                           mult_28_C96_n1051);
   mult_28_C96_U1057 : NAN3D1 port map( A1 => mult_28_C96_n1004, A2 => 
                           mult_28_C96_n1006, A3 => mult_28_C96_n1005, Z => 
                           mult_28_C96_n429);
   mult_28_C96_U1056 : NAN2DL port map( A1 => mult_28_C96_n432, A2 => 
                           mult_28_C96_n443, Z => mult_28_C96_n1005);
   mult_28_C96_U1055 : NAN2DL port map( A1 => mult_28_C96_n432, A2 => 
                           mult_28_C96_n434, Z => mult_28_C96_n1004);
   mult_28_C96_U1054 : EXOR2D1 port map( A1 => mult_28_C96_n1003, A2 => 
                           mult_28_C96_n432, Z => mult_28_C96_n430);
   mult_28_C96_U1053 : EXOR2D1 port map( A1 => mult_28_C96_n443, A2 => 
                           mult_28_C96_n434, Z => mult_28_C96_n1003);
   mult_28_C96_U1052 : OAI22D1 port map( A1 => mult_28_C96_n758, A2 => 
                           mult_28_C96_n12, B1 => mult_28_C96_n757, B2 => 
                           mult_28_C96_n9, Z => mult_28_C96_n623);
   mult_28_C96_U1051 : EXNOR2DL port map( A1 => n43, A2 => coeff_memory_7_port,
                           Z => mult_28_C96_n730);
   mult_28_C96_U1050 : NAN3D1 port map( A1 => mult_28_C96_n1014, A2 => 
                           mult_28_C96_n1016, A3 => mult_28_C96_n1015, Z => 
                           mult_28_C96_n457);
   mult_28_C96_U1049 : NAN2D1 port map( A1 => mult_28_C96_n288, A2 => 
                           mult_28_C96_n1066, Z => mult_28_C96_n67);
   mult_28_C96_U1048 : EXNOR2DL port map( A1 => n43, A2 => coeff_memory_5_port,
                           Z => mult_28_C96_n747);
   mult_28_C96_U1047 : EXNOR2DL port map( A1 => n43, A2 => coeff_memory_3_port,
                           Z => mult_28_C96_n764);
   mult_28_C96_U1046 : EXNOR2DL port map( A1 => n43, A2 => coeff_memory_1_port,
                           Z => mult_28_C96_n781);
   mult_28_C96_U1045 : EXNOR2DL port map( A1 => y_3_port, A2 => 
                           coeff_memory_13_port, Z => mult_28_C96_n678);
   mult_28_C96_U1044 : EXNOR2D2 port map( A1 => y_3_port, A2 => 
                           coeff_memory_9_port, Z => mult_28_C96_n712);
   mult_28_C96_U1043 : EXNOR2DL port map( A1 => y_3_port, A2 => 
                           coeff_memory_7_port, Z => mult_28_C96_n729);
   mult_28_C96_U1042 : EXNOR2D2 port map( A1 => y_3_port, A2 => 
                           coeff_memory_5_port, Z => mult_28_C96_n746);
   mult_28_C96_U1041 : EXNOR2D2 port map( A1 => y_3_port, A2 => 
                           coeff_memory_1_port, Z => mult_28_C96_n780);
   mult_28_C96_U1040 : EXNOR2D2 port map( A1 => y_3_port, A2 => 
                           coeff_memory_15_port, Z => mult_28_C96_n661);
   mult_28_C96_U1039 : INVDL port map( A => mult_28_C96_n52, Z => 
                           mult_28_C96_n129);
   mult_28_C96_U1038 : OAI21DL port map( A1 => mult_28_C96_n934, A2 => 
                           mult_28_C96_n108, B => mult_28_C96_n109, Z => 
                           mult_28_C96_n107);
   mult_28_C96_U1037 : OA21DL port map( A1 => mult_28_C96_n217, A2 => 
                           mult_28_C96_n223, B => mult_28_C96_n1027, Z => 
                           mult_28_C96_n214);
   mult_28_C96_U1036 : EXNOR2D2 port map( A1 => n33, A2 => coeff_memory_7_port,
                           Z => mult_28_C96_n727);
   mult_28_C96_U1035 : EXNOR2DL port map( A1 => y_11_port, A2 => 
                           coeff_memory_7_port, Z => mult_28_C96_n721);
   mult_28_C96_U1034 : EXNOR2DL port map( A1 => y_7_port, A2 => 
                           coeff_memory_5_port, Z => mult_28_C96_n742);
   mult_28_C96_U1033 : NAN2D1 port map( A1 => mult_28_C96_n437, A2 => 
                           mult_28_C96_n435, Z => mult_28_C96_n1001);
   mult_28_C96_U1032 : NAN2D1 port map( A1 => mult_28_C96_n902, A2 => 
                           mult_28_C96_n435, Z => mult_28_C96_n1000);
   mult_28_C96_U1031 : NAN2D1 port map( A1 => mult_28_C96_n902, A2 => 
                           mult_28_C96_n437, Z => mult_28_C96_n999);
   mult_28_C96_U1030 : EXOR2D1 port map( A1 => mult_28_C96_n619, A2 => 
                           mult_28_C96_n437, Z => mult_28_C96_n998);
   mult_28_C96_U1029 : NAN3D2 port map( A1 => mult_28_C96_n997, A2 => 
                           mult_28_C96_n996, A3 => mult_28_C96_n995, Z => 
                           mult_28_C96_n435);
   mult_28_C96_U1028 : NAN2D1 port map( A1 => mult_28_C96_n605, A2 => 
                           mult_28_C96_n590, Z => mult_28_C96_n997);
   mult_28_C96_U1027 : NAN2D1 port map( A1 => mult_28_C96_n605, A2 => 
                           mult_28_C96_n449, Z => mult_28_C96_n996);
   mult_28_C96_U1026 : EXOR3D1 port map( A1 => mult_28_C96_n449, A2 => 
                           mult_28_C96_n590, A3 => mult_28_C96_n905, Z => 
                           mult_28_C96_n436);
   mult_28_C96_U1025 : EXOR2D1 port map( A1 => mult_28_C96_n539, A2 => 
                           mult_28_C96_n569, Z => mult_28_C96_n1029);
   mult_28_C96_U1024 : EXNOR2D1 port map( A1 => n42, A2 => coeff_memory_1_port,
                           Z => mult_28_C96_n773);
   mult_28_C96_U1023 : EXNOR2DL port map( A1 => n43, A2 => coeff_memory_9_port,
                           Z => mult_28_C96_n713);
   mult_28_C96_U1022 : EXNOR2D2 port map( A1 => n43, A2 => coeff_memory_13_port
                           , Z => mult_28_C96_n679);
   mult_28_C96_U1021 : EXNOR2D2 port map( A1 => n42, A2 => coeff_memory_3_port,
                           Z => mult_28_C96_n756);
   mult_28_C96_U1020 : AOI21DL port map( A1 => mult_28_C96_n202, A2 => 
                           mult_28_C96_n288, B => mult_28_C96_n199, Z => 
                           mult_28_C96_n197);
   mult_28_C96_U1019 : EXNOR2D2 port map( A1 => n43, A2 => coeff_memory_11_port
                           , Z => mult_28_C96_n696);
   mult_28_C96_U1018 : NAN2D1 port map( A1 => mult_28_C96_n354, A2 => 
                           mult_28_C96_n363, Z => mult_28_C96_n173);
   mult_28_C96_U1017 : EXNOR2D1 port map( A1 => n34, A2 => coeff_memory_13_port
                           , Z => mult_28_C96_n680);
   mult_28_C96_U1016 : BUFDL port map( A => mult_28_C96_n680, Z => 
                           mult_28_C96_n994);
   mult_28_C96_U1015 : EXNOR2D2 port map( A1 => y_14_port, A2 => 
                           coeff_memory_5_port, Z => mult_28_C96_n735);
   mult_28_C96_U1014 : EXNOR2D2 port map( A1 => y_13_port, A2 => 
                           coeff_memory_5_port, Z => mult_28_C96_n736);
   mult_28_C96_U1013 : EXOR3D1 port map( A1 => mult_28_C96_n368, A2 => 
                           mult_28_C96_n377, A3 => mult_28_C96_n1064, Z => 
                           mult_28_C96_n1065);
   mult_28_C96_U1012 : NAN3D2 port map( A1 => mult_28_C96_n990, A2 => 
                           mult_28_C96_n991, A3 => mult_28_C96_n992, Z => 
                           mult_28_C96_n377);
   mult_28_C96_U1011 : NAN2DL port map( A1 => mult_28_C96_n391, A2 => 
                           mult_28_C96_n384, Z => mult_28_C96_n992);
   mult_28_C96_U1010 : NAN2DL port map( A1 => mult_28_C96_n382, A2 => 
                           mult_28_C96_n384, Z => mult_28_C96_n991);
   mult_28_C96_U1009 : NAN2DL port map( A1 => mult_28_C96_n391, A2 => 
                           mult_28_C96_n382, Z => mult_28_C96_n990);
   mult_28_C96_U1008 : EXOR3D1 port map( A1 => mult_28_C96_n382, A2 => 
                           mult_28_C96_n384, A3 => mult_28_C96_n979, Z => 
                           mult_28_C96_n378);
   mult_28_C96_U1007 : NOR2D1 port map( A1 => mult_28_C96_n442, A2 => 
                           mult_28_C96_n453, Z => mult_28_C96_n217);
   mult_28_C96_U1006 : EXNOR2DL port map( A1 => y_8_port, A2 => 
                           coeff_memory_11_port, Z => mult_28_C96_n690);
   mult_28_C96_U1005 : NAN3D2 port map( A1 => mult_28_C96_n987, A2 => 
                           mult_28_C96_n989, A3 => mult_28_C96_n988, Z => 
                           mult_28_C96_n385);
   mult_28_C96_U1004 : NAN2D1 port map( A1 => mult_28_C96_n528, A2 => 
                           mult_28_C96_n993, Z => mult_28_C96_n989);
   mult_28_C96_U1003 : NAN2D1 port map( A1 => mult_28_C96_n993, A2 => 
                           mult_28_C96_n541, Z => mult_28_C96_n988);
   mult_28_C96_U1002 : NAN2D1 port map( A1 => mult_28_C96_n541, A2 => 
                           mult_28_C96_n528, Z => mult_28_C96_n987);
   mult_28_C96_U1001 : EXOR2D1 port map( A1 => mult_28_C96_n986, A2 => 
                           mult_28_C96_n541, Z => mult_28_C96_n386);
   mult_28_C96_U1000 : EXOR2D1 port map( A1 => mult_28_C96_n993, A2 => 
                           mult_28_C96_n528, Z => mult_28_C96_n986);
   mult_28_C96_U999 : INVD1 port map( A => mult_28_C96_n150, Z => 
                           mult_28_C96_n148);
   mult_28_C96_U998 : EXOR3D2 port map( A1 => mult_28_C96_n425, A2 => 
                           mult_28_C96_n588, A3 => mult_28_C96_n573, Z => 
                           mult_28_C96_n410);
   mult_28_C96_U997 : NAN2DL port map( A1 => mult_28_C96_n588, A2 => 
                           mult_28_C96_n425, Z => mult_28_C96_n1047);
   mult_28_C96_U996 : NAN2DL port map( A1 => mult_28_C96_n588, A2 => 
                           mult_28_C96_n573, Z => mult_28_C96_n1046);
   mult_28_C96_U995 : EXNOR2DL port map( A1 => y_3_port, A2 => 
                           coeff_memory_3_port, Z => mult_28_C96_n763);
   mult_28_C96_U994 : NAN3D2 port map( A1 => mult_28_C96_n985, A2 => 
                           mult_28_C96_n983, A3 => mult_28_C96_n984, Z => 
                           mult_28_C96_n393);
   mult_28_C96_U993 : NAN2D1 port map( A1 => mult_28_C96_n906, A2 => 
                           mult_28_C96_n587, Z => mult_28_C96_n985);
   mult_28_C96_U992 : NAN2D1 port map( A1 => mult_28_C96_n602, A2 => 
                           mult_28_C96_n953, Z => mult_28_C96_n983);
   mult_28_C96_U991 : EXOR3D2 port map( A1 => mult_28_C96_n398, A2 => 
                           mult_28_C96_n587, A3 => mult_28_C96_n906, Z => 
                           mult_28_C96_n394);
   mult_28_C96_U990 : EXNOR2D2 port map( A1 => y_12_port, A2 => 
                           coeff_memory_3_port, Z => mult_28_C96_n754);
   mult_28_C96_U989 : OAI22D1 port map( A1 => mult_28_C96_n656, A2 => 
                           mult_28_C96_n48, B1 => mult_28_C96_n655, B2 => 
                           mult_28_C96_n46, Z => mult_28_C96_n333);
   mult_28_C96_U988 : OAI22DL port map( A1 => mult_28_C96_n691, A2 => 
                           mult_28_C96_n36, B1 => mult_28_C96_n690, B2 => 
                           mult_28_C96_n34, Z => mult_28_C96_n556);
   mult_28_C96_U987 : EXNOR2D1 port map( A1 => y_11_port, A2 => 
                           coeff_memory_7_port, Z => mult_28_C96_n1002);
   mult_28_C96_U986 : EXNOR2D2 port map( A1 => y_11_port, A2 => 
                           coeff_memory_3_port, Z => mult_28_C96_n755);
   mult_28_C96_U985 : EXOR2D1 port map( A1 => mult_28_C96_n1009, A2 => 
                           mult_28_C96_n418, Z => mult_28_C96_n416);
   mult_28_C96_U984 : ADFULD1 port map( A => mult_28_C96_n561, B => 
                           mult_28_C96_n452, CI => mult_28_C96_n576, CO => 
                           mult_28_C96_n449, S => mult_28_C96_n450);
   mult_28_C96_U983 : NAN2D1 port map( A1 => mult_28_C96_n449, A2 => 
                           mult_28_C96_n590, Z => mult_28_C96_n995);
   mult_28_C96_U982 : NAN3D2 port map( A1 => mult_28_C96_n999, A2 => 
                           mult_28_C96_n1000, A3 => mult_28_C96_n1001, Z => 
                           mult_28_C96_n419);
   mult_28_C96_U981 : OAI22DL port map( A1 => mult_28_C96_n705, A2 => 
                           mult_28_C96_n30, B1 => mult_28_C96_n704, B2 => 
                           mult_28_C96_n28, Z => mult_28_C96_n570);
   mult_28_C96_U980 : NAN3D1 port map( A1 => mult_28_C96_n980, A2 => 
                           mult_28_C96_n982, A3 => mult_28_C96_n981, Z => 
                           mult_28_C96_n369);
   mult_28_C96_U979 : NAN2DL port map( A1 => mult_28_C96_n570, A2 => 
                           mult_28_C96_n600, Z => mult_28_C96_n982);
   mult_28_C96_U978 : NAN2DL port map( A1 => mult_28_C96_n385, A2 => 
                           mult_28_C96_n600, Z => mult_28_C96_n981);
   mult_28_C96_U977 : NAN2DL port map( A1 => mult_28_C96_n385, A2 => 
                           mult_28_C96_n570, Z => mult_28_C96_n980);
   mult_28_C96_U976 : EXOR3D2 port map( A1 => mult_28_C96_n935, A2 => 
                           mult_28_C96_n385, A3 => mult_28_C96_n570, Z => 
                           mult_28_C96_n370);
   mult_28_C96_U975 : OAI21DL port map( A1 => mult_28_C96_n164, A2 => 
                           mult_28_C96_n154, B => mult_28_C96_n155, Z => 
                           mult_28_C96_n153);
   mult_28_C96_U974 : NOR2D1 port map( A1 => mult_28_C96_n163, A2 => 
                           mult_28_C96_n154, Z => mult_28_C96_n152);
   mult_28_C96_U973 : NAN3D1 port map( A1 => mult_28_C96_n1038, A2 => 
                           mult_28_C96_n1039, A3 => mult_28_C96_n1040, Z => 
                           mult_28_C96_n405);
   mult_28_C96_U972 : ADHALFD2 port map( A => mult_28_C96_n513, B => 
                           mult_28_C96_n530, CO => mult_28_C96_n427, S => 
                           mult_28_C96_n428);
   mult_28_C96_U971 : INVD1 port map( A => mult_28_C96_n978, Z => 
                           mult_28_C96_n979);
   mult_28_C96_U970 : INVDL port map( A => mult_28_C96_n391, Z => 
                           mult_28_C96_n978);
   mult_28_C96_U969 : BUFDL port map( A => mult_28_C96_n622, Z => 
                           mult_28_C96_n977);
   mult_28_C96_U968 : EXOR2DL port map( A1 => mult_28_C96_n469, A2 => 
                           mult_28_C96_n607, Z => mult_28_C96_n1013);
   mult_28_C96_U967 : EXOR2D1 port map( A1 => mult_28_C96_n1013, A2 => 
                           mult_28_C96_n977, Z => mult_28_C96_n458);
   mult_28_C96_U966 : ADFULDL port map( A => mult_28_C96_n333, B => 
                           mult_28_C96_n525, CI => mult_28_C96_n550, CO => 
                           mult_28_C96_n325, S => mult_28_C96_n326);
   mult_28_C96_U965 : EXNOR2DL port map( A1 => y_8_port, A2 => 
                           coeff_memory_15_port, Z => mult_28_C96_n656);
   mult_28_C96_U964 : NAN3D1 port map( A1 => mult_28_C96_n974, A2 => 
                           mult_28_C96_n976, A3 => mult_28_C96_n975, Z => 
                           mult_28_C96_n447);
   mult_28_C96_U963 : NAN2DL port map( A1 => mult_28_C96_n591, A2 => 
                           mult_28_C96_n461, Z => mult_28_C96_n975);
   mult_28_C96_U962 : NAN2DL port map( A1 => mult_28_C96_n591, A2 => 
                           mult_28_C96_n606, Z => mult_28_C96_n974);
   mult_28_C96_U961 : OAI21D1 port map( A1 => mult_28_C96_n187, A2 => 
                           mult_28_C96_n179, B => mult_28_C96_n180, Z => 
                           mult_28_C96_n178);
   mult_28_C96_U960 : NAN3D1 port map( A1 => mult_28_C96_n971, A2 => 
                           mult_28_C96_n973, A3 => mult_28_C96_n972, Z => 
                           mult_28_C96_n353);
   mult_28_C96_U959 : NAN2DL port map( A1 => mult_28_C96_n365, A2 => 
                           mult_28_C96_n358, Z => mult_28_C96_n973);
   mult_28_C96_U958 : NAN2DL port map( A1 => mult_28_C96_n356, A2 => 
                           mult_28_C96_n365, Z => mult_28_C96_n971);
   mult_28_C96_U957 : EXOR2D1 port map( A1 => mult_28_C96_n970, A2 => 
                           mult_28_C96_n356, Z => mult_28_C96_n354);
   mult_28_C96_U956 : EXOR2D1 port map( A1 => mult_28_C96_n358, A2 => 
                           mult_28_C96_n365, Z => mult_28_C96_n970);
   mult_28_C96_U955 : EXNOR2DL port map( A1 => y_9_port, A2 => 
                           coeff_memory_11_port, Z => mult_28_C96_n689);
   mult_28_C96_U954 : EXNOR2D2 port map( A1 => n34, A2 => coeff_memory_11_port,
                           Z => mult_28_C96_n697);
   mult_28_C96_U953 : BUFDL port map( A => mult_28_C96_n912, Z => 
                           mult_28_C96_n968);
   mult_28_C96_U952 : EXNOR2D2 port map( A1 => y_12_port, A2 => 
                           coeff_memory_1_port, Z => mult_28_C96_n771);
   mult_28_C96_U951 : INVDL port map( A => mult_28_C96_n396, Z => 
                           mult_28_C96_n967);
   mult_28_C96_U950 : EXOR2D2 port map( A1 => mult_28_C96_n633, A2 => 
                           mult_28_C96_n421, Z => mult_28_C96_n1037);
   mult_28_C96_U949 : NAN3D2 port map( A1 => mult_28_C96_n963, A2 => 
                           mult_28_C96_n965, A3 => mult_28_C96_n964, Z => 
                           mult_28_C96_n357);
   mult_28_C96_U948 : NAN2DL port map( A1 => mult_28_C96_n371, A2 => 
                           mult_28_C96_n599, Z => mult_28_C96_n965);
   mult_28_C96_U947 : NAN2D1 port map( A1 => mult_28_C96_n362, A2 => 
                           mult_28_C96_n599, Z => mult_28_C96_n964);
   mult_28_C96_U946 : NAN2D1 port map( A1 => mult_28_C96_n362, A2 => 
                           mult_28_C96_n371, Z => mult_28_C96_n963);
   mult_28_C96_U945 : EXOR2D1 port map( A1 => mult_28_C96_n599, A2 => 
                           mult_28_C96_n371, Z => mult_28_C96_n962);
   mult_28_C96_U944 : OAI22D1 port map( A1 => mult_28_C96_n708, A2 => 
                           mult_28_C96_n30, B1 => mult_28_C96_n919, B2 => 
                           mult_28_C96_n28, Z => mult_28_C96_n573);
   mult_28_C96_U943 : NAN3D1 port map( A1 => mult_28_C96_n1046, A2 => 
                           mult_28_C96_n1048, A3 => mult_28_C96_n1047, Z => 
                           mult_28_C96_n409);
   mult_28_C96_U942 : NAN2DL port map( A1 => mult_28_C96_n481, A2 => 
                           mult_28_C96_n474, Z => mult_28_C96_n961);
   mult_28_C96_U941 : OA21M20D1 port map( A1 => mult_28_C96_n1077, A2 => 
                           mult_28_C96_n1072, B => mult_28_C96_n961, Z => 
                           mult_28_C96_n232);
   mult_28_C96_U940 : EXNOR2D2 port map( A1 => y_6_port, A2 => 
                           coeff_memory_9_port, Z => mult_28_C96_n709);
   mult_28_C96_U939 : EXNOR2D2 port map( A1 => y_6_port, A2 => 
                           coeff_memory_7_port, Z => mult_28_C96_n726);
   mult_28_C96_U938 : OAI22DL port map( A1 => mult_28_C96_n654, A2 => 
                           mult_28_C96_n46, B1 => mult_28_C96_n655, B2 => 
                           mult_28_C96_n48, Z => mult_28_C96_n525);
   mult_28_C96_U937 : OAI22D1 port map( A1 => mult_28_C96_n775, A2 => 
                           mult_28_C96_n6, B1 => mult_28_C96_n774, B2 => 
                           mult_28_C96_n824, Z => mult_28_C96_n640);
   mult_28_C96_U936 : EXNOR2D2 port map( A1 => y_15_port, A2 => 
                           coeff_memory_5_port, Z => mult_28_C96_n734);
   mult_28_C96_U935 : INVDL port map( A => mult_28_C96_n167, Z => 
                           mult_28_C96_n283);
   mult_28_C96_U934 : OAI22DL port map( A1 => mult_28_C96_n701, A2 => 
                           mult_28_C96_n30, B1 => mult_28_C96_n700, B2 => 
                           mult_28_C96_n28, Z => mult_28_C96_n566);
   mult_28_C96_U933 : NAN3D1 port map( A1 => mult_28_C96_n957, A2 => 
                           mult_28_C96_n959, A3 => mult_28_C96_n958, Z => 
                           mult_28_C96_n329);
   mult_28_C96_U932 : NAN2D1 port map( A1 => mult_28_C96_n341, A2 => 
                           mult_28_C96_n566, Z => mult_28_C96_n959);
   mult_28_C96_U931 : NAN2DL port map( A1 => mult_28_C96_n339, A2 => 
                           mult_28_C96_n566, Z => mult_28_C96_n958);
   mult_28_C96_U930 : NAN2DL port map( A1 => mult_28_C96_n339, A2 => 
                           mult_28_C96_n341, Z => mult_28_C96_n957);
   mult_28_C96_U929 : EXOR2D1 port map( A1 => mult_28_C96_n956, A2 => 
                           mult_28_C96_n339, Z => mult_28_C96_n330);
   mult_28_C96_U928 : EXOR2D1 port map( A1 => mult_28_C96_n566, A2 => 
                           mult_28_C96_n341, Z => mult_28_C96_n956);
   mult_28_C96_U927 : NOR2DL port map( A1 => mult_28_C96_n482, A2 => 
                           mult_28_C96_n489, Z => mult_28_C96_n955);
   mult_28_C96_U926 : NAN2M1D1 port map( A1 => mult_28_C96_n955, A2 => 
                           mult_28_C96_n1077, Z => mult_28_C96_n1068);
   mult_28_C96_U925 : INVD1 port map( A => mult_28_C96_n161, Z => 
                           mult_28_C96_n163);
   mult_28_C96_U924 : EXNOR2D2 port map( A1 => y_9_port, A2 => 
                           coeff_memory_9_port, Z => mult_28_C96_n706);
   mult_28_C96_U923 : EXNOR2D2 port map( A1 => y_9_port, A2 => 
                           coeff_memory_5_port, Z => mult_28_C96_n740);
   mult_28_C96_U922 : OAI21DL port map( A1 => mult_28_C96_n201, A2 => 
                           mult_28_C96_n913, B => mult_28_C96_n196, Z => 
                           mult_28_C96_n954);
   mult_28_C96_U921 : EXOR3D1 port map( A1 => mult_28_C96_n400, A2 => 
                           mult_28_C96_n413, A3 => mult_28_C96_n911, Z => 
                           mult_28_C96_n953);
   mult_28_C96_U920 : EXNOR2D2 port map( A1 => n33, A2 => coeff_memory_5_port, 
                           Z => mult_28_C96_n744);
   mult_28_C96_U919 : BUFDL port map( A => mult_28_C96_n161, Z => 
                           mult_28_C96_n952);
   mult_28_C96_U918 : EXNOR2DL port map( A1 => n42, A2 => coeff_memory_9_port, 
                           Z => mult_28_C96_n705);
   mult_28_C96_U917 : NAN2DL port map( A1 => mult_28_C96_n356, A2 => 
                           mult_28_C96_n358, Z => mult_28_C96_n972);
   mult_28_C96_U916 : EXOR2D4 port map( A1 => mult_28_C96_n962, A2 => 
                           mult_28_C96_n362, Z => mult_28_C96_n358);
   mult_28_C96_U915 : OAI22D1 port map( A1 => mult_28_C96_n717, A2 => 
                           mult_28_C96_n22, B1 => mult_28_C96_n718, B2 => 
                           mult_28_C96_n24, Z => mult_28_C96_n583);
   mult_28_C96_U914 : OAI22D1 port map( A1 => mult_28_C96_n30, A2 => 
                           mult_28_C96_n706, B1 => mult_28_C96_n28, B2 => 
                           mult_28_C96_n705, Z => mult_28_C96_n571);
   mult_28_C96_U913 : NAN3M1D1 port map( A1 => mult_28_C96_n929, A2 => 
                           mult_28_C96_n1094, A3 => mult_28_C96_n1093, Z => 
                           mult_28_C96_n375);
   mult_28_C96_U912 : EXOR3D1 port map( A1 => mult_28_C96_n527, A2 => 
                           mult_28_C96_n373, A3 => mult_28_C96_n554, Z => 
                           mult_28_C96_n362);
   mult_28_C96_U911 : INVDL port map( A => mult_28_C96_n616, Z => 
                           mult_28_C96_n951);
   mult_28_C96_U910 : NAN2M1D1 port map( A1 => mult_28_C96_n951, A2 => 
                           mult_28_C96_n393, Z => mult_28_C96_n1055);
   mult_28_C96_U909 : INVDL port map( A => mult_28_C96_n168, Z => 
                           mult_28_C96_n950);
   mult_28_C96_U908 : INVDL port map( A => mult_28_C96_n173, Z => 
                           mult_28_C96_n949);
   mult_28_C96_U907 : AOI21D1 port map( A1 => mult_28_C96_n283, A2 => 
                           mult_28_C96_n949, B => mult_28_C96_n950, Z => 
                           mult_28_C96_n164);
   mult_28_C96_U906 : INVDL port map( A => mult_28_C96_n454, Z => 
                           mult_28_C96_n948);
   mult_28_C96_U905 : OAI21M10D1 port map( A1 => mult_28_C96_n948, A2 => 
                           mult_28_C96_n463, B => mult_28_C96_n215, Z => 
                           mult_28_C96_n213);
   mult_28_C96_U904 : INVDL port map( A => mult_28_C96_n203, Z => 
                           mult_28_C96_n202);
   mult_28_C96_U903 : BUFD1 port map( A => mult_28_C96_n426, Z => 
                           mult_28_C96_n1050);
   mult_28_C96_U902 : EXNOR2D1 port map( A1 => n34, A2 => coeff_memory_15_port,
                           Z => mult_28_C96_n663);
   mult_28_C96_U901 : EXNOR2D2 port map( A1 => y_13_port, A2 => 
                           coeff_memory_1_port, Z => mult_28_C96_n770);
   mult_28_C96_U900 : EXNOR2D2 port map( A1 => y_13_port, A2 => 
                           coeff_memory_3_port, Z => mult_28_C96_n753);
   mult_28_C96_U899 : NAN2D1 port map( A1 => mult_28_C96_n419, A2 => 
                           mult_28_C96_n408, Z => mult_28_C96_n1024);
   mult_28_C96_U898 : NAN3D2 port map( A1 => mult_28_C96_n1024, A2 => 
                           mult_28_C96_n1026, A3 => mult_28_C96_n1025, Z => 
                           mult_28_C96_n403);
   mult_28_C96_U897 : EXNOR2DL port map( A1 => y_15_port, A2 => 
                           coeff_memory_11_port, Z => mult_28_C96_n683);
   mult_28_C96_U896 : EXNOR2DL port map( A1 => y_15_port, A2 => 
                           coeff_memory_13_port, Z => mult_28_C96_n666);
   mult_28_C96_U895 : EXNOR2D2 port map( A1 => mult_28_C96_n1008, A2 => 
                           coeff_memory_13_port, Z => mult_28_C96_n672);
   mult_28_C96_U894 : NOR2D1 port map( A1 => mult_28_C96_n430, A2 => 
                           mult_28_C96_n441, Z => mult_28_C96_n209);
   mult_28_C96_U893 : EXNOR2DL port map( A1 => y_11_port, A2 => 
                           coeff_memory_5_port, Z => mult_28_C96_n947);
   mult_28_C96_U892 : EXNOR2DL port map( A1 => y_15_port, A2 => 
                           coeff_memory_9_port, Z => mult_28_C96_n700);
   mult_28_C96_U891 : NAN2DL port map( A1 => mult_28_C96_n633, A2 => 
                           mult_28_C96_n421, Z => mult_28_C96_n1038);
   mult_28_C96_U890 : NAN2DL port map( A1 => mult_28_C96_n421, A2 => 
                           mult_28_C96_n423, Z => mult_28_C96_n1040);
   mult_28_C96_U889 : NAN2DL port map( A1 => mult_28_C96_n434, A2 => 
                           mult_28_C96_n443, Z => mult_28_C96_n1006);
   mult_28_C96_U888 : EXOR2D1 port map( A1 => mult_28_C96_n998, A2 => 
                           mult_28_C96_n927, Z => mult_28_C96_n420);
   mult_28_C96_U887 : NAN3D2 port map( A1 => mult_28_C96_n944, A2 => 
                           mult_28_C96_n945, A3 => mult_28_C96_n946, Z => 
                           mult_28_C96_n433);
   mult_28_C96_U886 : NAN2DL port map( A1 => mult_28_C96_n635, A2 => 
                           mult_28_C96_n438, Z => mult_28_C96_n946);
   mult_28_C96_U885 : NAN2DL port map( A1 => mult_28_C96_n620, A2 => 
                           mult_28_C96_n438, Z => mult_28_C96_n945);
   mult_28_C96_U884 : NAN2DL port map( A1 => mult_28_C96_n620, A2 => 
                           mult_28_C96_n635, Z => mult_28_C96_n944);
   mult_28_C96_U883 : NAN3D1 port map( A1 => mult_28_C96_n941, A2 => 
                           mult_28_C96_n942, A3 => mult_28_C96_n943, Z => 
                           mult_28_C96_n437);
   mult_28_C96_U882 : NAN2DL port map( A1 => mult_28_C96_n560, A2 => 
                           mult_28_C96_n440, Z => mult_28_C96_n943);
   mult_28_C96_U881 : NAN2DL port map( A1 => mult_28_C96_n575, A2 => 
                           mult_28_C96_n440, Z => mult_28_C96_n942);
   mult_28_C96_U880 : NAN2DL port map( A1 => mult_28_C96_n575, A2 => 
                           mult_28_C96_n560, Z => mult_28_C96_n941);
   mult_28_C96_U879 : EXOR2D1 port map( A1 => mult_28_C96_n940, A2 => 
                           mult_28_C96_n438, Z => mult_28_C96_n434);
   mult_28_C96_U878 : EXOR2D1 port map( A1 => mult_28_C96_n635, A2 => 
                           mult_28_C96_n620, Z => mult_28_C96_n940);
   mult_28_C96_U877 : INVDL port map( A => mult_28_C96_n217, Z => 
                           mult_28_C96_n215);
   mult_28_C96_U876 : NAN3D1 port map( A1 => mult_28_C96_n937, A2 => 
                           mult_28_C96_n939, A3 => mult_28_C96_n938, Z => 
                           mult_28_C96_n441);
   mult_28_C96_U875 : NAN2DL port map( A1 => mult_28_C96_n455, A2 => 
                           mult_28_C96_n446, Z => mult_28_C96_n939);
   mult_28_C96_U874 : NAN2DL port map( A1 => mult_28_C96_n444, A2 => 
                           mult_28_C96_n446, Z => mult_28_C96_n938);
   mult_28_C96_U873 : NAN2DL port map( A1 => mult_28_C96_n444, A2 => 
                           mult_28_C96_n455, Z => mult_28_C96_n937);
   mult_28_C96_U872 : EXOR2D1 port map( A1 => mult_28_C96_n936, A2 => 
                           mult_28_C96_n444, Z => mult_28_C96_n442);
   mult_28_C96_U871 : EXOR2D1 port map( A1 => mult_28_C96_n446, A2 => 
                           mult_28_C96_n455, Z => mult_28_C96_n936);
   mult_28_C96_U870 : EXNOR2DL port map( A1 => y_9_port, A2 => 
                           coeff_memory_3_port, Z => mult_28_C96_n757);
   mult_28_C96_U869 : EXOR3D2 port map( A1 => mult_28_C96_n410, A2 => 
                           mult_28_C96_n419, A3 => mult_28_C96_n408, Z => 
                           mult_28_C96_n404);
   mult_28_C96_U868 : NAN2D1 port map( A1 => mult_28_C96_n953, A2 => 
                           mult_28_C96_n587, Z => mult_28_C96_n984);
   mult_28_C96_U867 : EXOR3D1 port map( A1 => mult_28_C96_n634, A2 => 
                           mult_28_C96_n604, A3 => mult_28_C96_n1050, Z => 
                           mult_28_C96_n422);
   mult_28_C96_U866 : EXNOR2DL port map( A1 => y_8_port, A2 => 
                           coeff_memory_5_port, Z => mult_28_C96_n741);
   mult_28_C96_U865 : EXNOR2D2 port map( A1 => y_8_port, A2 => 
                           coeff_memory_7_port, Z => mult_28_C96_n724);
   mult_28_C96_U864 : OAI22D1 port map( A1 => mult_28_C96_n735, A2 => 
                           mult_28_C96_n18, B1 => mult_28_C96_n734, B2 => 
                           mult_28_C96_n16, Z => mult_28_C96_n935);
   mult_28_C96_U863 : BUFD2 port map( A => mult_28_C96_n399, Z => 
                           mult_28_C96_n993);
   mult_28_C96_U862 : INVD1 port map( A => mult_28_C96_n399, Z => 
                           mult_28_C96_n400);
   mult_28_C96_U861 : AOI21D1 port map( A1 => mult_28_C96_n162, A2 => 
                           mult_28_C96_n969, B => mult_28_C96_n133, Z => 
                           mult_28_C96_n934);
   mult_28_C96_U860 : EXNOR2D1 port map( A1 => mult_28_C96_n208, A2 => 
                           mult_28_C96_n68, Z => m5_1);
   mult_28_C96_U859 : EXNOR2D2 port map( A1 => y_4_port, A2 => 
                           coeff_memory_15_port, Z => mult_28_C96_n660);
   mult_28_C96_U858 : INVD1 port map( A => mult_28_C96_n931, Z => 
                           mult_28_C96_n932);
   mult_28_C96_U857 : INVDL port map( A => y_12_port, Z => mult_28_C96_n931);
   mult_28_C96_U856 : ADFULD1 port map( A => mult_28_C96_n621, B => 
                           mult_28_C96_n450, CI => mult_28_C96_n636, CO => 
                           mult_28_C96_n445, S => mult_28_C96_n446);
   mult_28_C96_U855 : NOR2DL port map( A1 => mult_28_C96_n464, A2 => 
                           mult_28_C96_n473, Z => mult_28_C96_n930);
   mult_28_C96_U854 : AOI21M10D1 port map( A1 => mult_28_C96_n930, A2 => 
                           mult_28_C96_n230, B => mult_28_C96_n1079, Z => 
                           mult_28_C96_n225);
   mult_28_C96_U853 : NOR2DL port map( A1 => mult_28_C96_n206, A2 => 
                           mult_28_C96_n209, Z => mult_28_C96_n204);
   mult_28_C96_U852 : NAN2M1DL port map( A1 => mult_28_C96_n209, A2 => 
                           mult_28_C96_n210, Z => mult_28_C96_n69);
   mult_28_C96_U851 : NAN2DL port map( A1 => mult_28_C96_n606, A2 => 
                           mult_28_C96_n461, Z => mult_28_C96_n976);
   mult_28_C96_U850 : EXOR3D1 port map( A1 => mult_28_C96_n461, A2 => 
                           mult_28_C96_n591, A3 => mult_28_C96_n606, Z => 
                           mult_28_C96_n448);
   mult_28_C96_U849 : ADHALFD2 port map( A => mult_28_C96_n563, B => 
                           mult_28_C96_n515, CO => mult_28_C96_n471, S => 
                           mult_28_C96_n472);
   mult_28_C96_U848 : AND2DL port map( A1 => mult_28_C96_n389, A2 => 
                           mult_28_C96_n380, Z => mult_28_C96_n929);
   mult_28_C96_U847 : INVDL port map( A => mult_28_C96_n92, Z => 
                           mult_28_C96_n276);
   mult_28_C96_U846 : INVD1 port map( A => mult_28_C96_n56, Z => 
                           mult_28_C96_n1017);
   mult_28_C96_U845 : INVDL port map( A => mult_28_C96_n53, Z => 
                           mult_28_C96_n128);
   mult_28_C96_U844 : NAN2D1 port map( A1 => mult_28_C96_n376, A2 => 
                           mult_28_C96_n387, Z => mult_28_C96_n187);
   mult_28_C96_U843 : OAI22D1 port map( A1 => mult_28_C96_n676, A2 => 
                           mult_28_C96_n42, B1 => mult_28_C96_n675, B2 => 
                           mult_28_C96_n40, Z => mult_28_C96_n541);
   mult_28_C96_U842 : EXOR3D1 port map( A1 => mult_28_C96_n575, A2 => 
                           mult_28_C96_n560, A3 => mult_28_C96_n440, Z => 
                           mult_28_C96_n438);
   mult_28_C96_U841 : INVD1 port map( A => mult_28_C96_n9, Z => 
                           mult_28_C96_n933);
   mult_28_C96_U840 : NOR2D1 port map( A1 => mult_28_C96_n312, A2 => 
                           mult_28_C96_n315, Z => mult_28_C96_n112);
   mult_28_C96_U839 : NAN2D1 port map( A1 => mult_28_C96_n161, A2 => 
                           mult_28_C96_n969, Z => mult_28_C96_n53);
   mult_28_C96_U838 : NOR2D1 port map( A1 => mult_28_C96_n311, A2 => 
                           mult_28_C96_n308, Z => mult_28_C96_n103);
   mult_28_C96_U837 : INVD1 port map( A => mult_28_C96_n118, Z => 
                           mult_28_C96_n960);
   mult_28_C96_U836 : OAI22D1 port map( A1 => mult_28_C96_n686, A2 => 
                           mult_28_C96_n36, B1 => mult_28_C96_n685, B2 => 
                           mult_28_C96_n34, Z => mult_28_C96_n551);
   mult_28_C96_U835 : NOR2D1 port map( A1 => mult_28_C96_n328, A2 => 
                           mult_28_C96_n335, Z => mult_28_C96_n149);
   mult_28_C96_U834 : EXNOR2D2 port map( A1 => mult_28_C96_n529, A2 => 
                           mult_28_C96_n427, Z => mult_28_C96_n414);
   mult_28_C96_U833 : INVBD32 port map( A => mult_28_C96_n933, Z => 
                           mult_28_C96_n928);
   mult_28_C96_U832 : OAI22D1 port map( A1 => mult_28_C96_n928, A2 => 
                           mult_28_C96_n752, B1 => mult_28_C96_n753, B2 => 
                           mult_28_C96_n12, Z => mult_28_C96_n618);
   mult_28_C96_U831 : BUFDL port map( A => mult_28_C96_n435, Z => 
                           mult_28_C96_n927);
   mult_28_C96_U830 : NAN3D1 port map( A1 => mult_28_C96_n924, A2 => 
                           mult_28_C96_n925, A3 => mult_28_C96_n926, Z => 
                           mult_28_C96_n481);
   mult_28_C96_U829 : NAN2DL port map( A1 => mult_28_C96_n486, A2 => 
                           mult_28_C96_n484, Z => mult_28_C96_n926);
   mult_28_C96_U828 : NAN2DL port map( A1 => mult_28_C96_n491, A2 => 
                           mult_28_C96_n484, Z => mult_28_C96_n925);
   mult_28_C96_U827 : NAN2D1 port map( A1 => mult_28_C96_n491, A2 => 
                           mult_28_C96_n486, Z => mult_28_C96_n924);
   mult_28_C96_U826 : NAN3D1 port map( A1 => mult_28_C96_n921, A2 => 
                           mult_28_C96_n922, A3 => mult_28_C96_n923, Z => 
                           mult_28_C96_n483);
   mult_28_C96_U825 : NAN2DL port map( A1 => mult_28_C96_n493, A2 => 
                           mult_28_C96_n640, Z => mult_28_C96_n923);
   mult_28_C96_U824 : NAN2DL port map( A1 => mult_28_C96_n625, A2 => 
                           mult_28_C96_n640, Z => mult_28_C96_n922);
   mult_28_C96_U823 : NAN2DL port map( A1 => mult_28_C96_n625, A2 => 
                           mult_28_C96_n493, Z => mult_28_C96_n921);
   mult_28_C96_U822 : EXOR2D1 port map( A1 => mult_28_C96_n920, A2 => 
                           mult_28_C96_n484, Z => mult_28_C96_n482);
   mult_28_C96_U821 : EXOR2D1 port map( A1 => mult_28_C96_n491, A2 => 
                           mult_28_C96_n486, Z => mult_28_C96_n920);
   mult_28_C96_U820 : EXOR3D2 port map( A1 => mult_28_C96_n625, A2 => 
                           mult_28_C96_n493, A3 => mult_28_C96_n640, Z => 
                           mult_28_C96_n484);
   mult_28_C96_U819 : NAN2D1 port map( A1 => mult_28_C96_n574, A2 => 
                           mult_28_C96_n439, Z => mult_28_C96_n1034);
   mult_28_C96_U818 : EXNOR2DL port map( A1 => y_4_port, A2 => 
                           coeff_memory_7_port, Z => mult_28_C96_n728);
   mult_28_C96_U817 : EXNOR2D2 port map( A1 => y_4_port, A2 => 
                           coeff_memory_11_port, Z => mult_28_C96_n694);
   mult_28_C96_U816 : EXNOR2D2 port map( A1 => y_4_port, A2 => 
                           coeff_memory_13_port, Z => mult_28_C96_n677);
   mult_28_C96_U815 : EXNOR2D2 port map( A1 => y_4_port, A2 => 
                           coeff_memory_9_port, Z => mult_28_C96_n711);
   mult_28_C96_U814 : EXOR2D1 port map( A1 => mult_28_C96_n1029, A2 => 
                           mult_28_C96_n584, Z => mult_28_C96_n360);
   mult_28_C96_U813 : INVD1 port map( A => mult_28_C96_n918, Z => 
                           mult_28_C96_n919);
   mult_28_C96_U812 : INVDL port map( A => mult_28_C96_n908, Z => 
                           mult_28_C96_n918);
   mult_28_C96_U811 : NOR2D1 port map( A1 => mult_28_C96_n354, A2 => 
                           mult_28_C96_n363, Z => mult_28_C96_n1028);
   mult_28_C96_U810 : NOR2D2 port map( A1 => mult_28_C96_n134, A2 => 
                           mult_28_C96_n154, Z => mult_28_C96_n969);
   mult_28_C96_U809 : AND2DL port map( A1 => mult_28_C96_n1078, A2 => 
                           mult_28_C96_n139, Z => mult_28_C96_n917);
   mult_28_C96_U808 : EXNOR2D2 port map( A1 => mult_28_C96_n140, A2 => 
                           mult_28_C96_n917, Z => m5_10);
   mult_28_C96_U807 : INVD1 port map( A => mult_28_C96_n915, Z => 
                           mult_28_C96_n916);
   mult_28_C96_U806 : INVDL port map( A => mult_28_C96_n663, Z => 
                           mult_28_C96_n915);
   mult_28_C96_U805 : INVDL port map( A => mult_28_C96_n286, Z => 
                           mult_28_C96_n914);
   mult_28_C96_U804 : NOR2D1 port map( A1 => mult_28_C96_n909, A2 => 
                           mult_28_C96_n401, Z => mult_28_C96_n195);
   mult_28_C96_U803 : NOR2D2 port map( A1 => mult_28_C96_n388, A2 => 
                           mult_28_C96_n401, Z => mult_28_C96_n913);
   mult_28_C96_U802 : AOI21DL port map( A1 => mult_28_C96_n141, A2 => 
                           mult_28_C96_n1020, B => mult_28_C96_n142, Z => 
                           mult_28_C96_n140);
   mult_28_C96_U801 : INVD1 port map( A => y_7_port, Z => mult_28_C96_n1041);
   mult_28_C96_U800 : EXNOR2D2 port map( A1 => y_7_port, A2 => 
                           coeff_memory_11_port, Z => mult_28_C96_n691);
   mult_28_C96_U799 : EXNOR2D2 port map( A1 => n42, A2 => coeff_memory_11_port,
                           Z => mult_28_C96_n688);
   mult_28_C96_U798 : AO21M20D1 port map( A1 => mult_28_C96_n52, A2 => 
                           mult_28_C96_n117, B => mult_28_C96_n960, Z => 
                           mult_28_C96_n116);
   mult_28_C96_U797 : NOR2DL port map( A1 => mult_28_C96_n913, A2 => 
                           mult_28_C96_n200, Z => mult_28_C96_n912);
   mult_28_C96_U796 : OAI22D1 port map( A1 => mult_28_C96_n677, A2 => 
                           mult_28_C96_n42, B1 => mult_28_C96_n676, B2 => 
                           mult_28_C96_n40, Z => mult_28_C96_n911);
   mult_28_C96_U795 : EXNOR2DL port map( A1 => y_14_port, A2 => 
                           coeff_memory_3_port, Z => mult_28_C96_n752);
   mult_28_C96_U794 : BUFDL port map( A => mult_28_C96_n179, Z => 
                           mult_28_C96_n910);
   mult_28_C96_U793 : EXNOR3D4 port map( A1 => mult_28_C96_n617, A2 => 
                           mult_28_C96_n409, A3 => mult_28_C96_n967, Z => 
                           mult_28_C96_n392);
   mult_28_C96_U792 : EXOR3D1 port map( A1 => mult_28_C96_n392, A2 => 
                           mult_28_C96_n403, A3 => mult_28_C96_n390, Z => 
                           mult_28_C96_n388);
   mult_28_C96_U791 : EXOR3D1 port map( A1 => mult_28_C96_n392, A2 => 
                           mult_28_C96_n403, A3 => mult_28_C96_n390, Z => 
                           mult_28_C96_n909);
   mult_28_C96_U790 : EXNOR2DL port map( A1 => y_6_port, A2 => 
                           coeff_memory_13_port, Z => mult_28_C96_n675);
   mult_28_C96_U789 : EXNOR2D1 port map( A1 => y_11_port, A2 => 
                           coeff_memory_9_port, Z => mult_28_C96_n704);
   mult_28_C96_U788 : EXNOR2D1 port map( A1 => y_8_port, A2 => 
                           coeff_memory_9_port, Z => mult_28_C96_n707);
   mult_28_C96_U787 : INVBD32 port map( A => mult_28_C96_n18, Z => 
                           mult_28_C96_n907);
   mult_28_C96_U786 : OAI22M10D1 port map( A1 => mult_28_C96_n907, A2 => 
                           mult_28_C96_n740, B1 => mult_28_C96_n1060, B2 => 
                           mult_28_C96_n16, Z => mult_28_C96_n605);
   mult_28_C96_U785 : OAI22DL port map( A1 => mult_28_C96_n737, A2 => 
                           mult_28_C96_n18, B1 => mult_28_C96_n736, B2 => 
                           mult_28_C96_n16, Z => mult_28_C96_n602);
   mult_28_C96_U784 : OAI22D1 port map( A1 => mult_28_C96_n737, A2 => 
                           mult_28_C96_n18, B1 => mult_28_C96_n736, B2 => 
                           mult_28_C96_n16, Z => mult_28_C96_n906);
   mult_28_C96_U783 : OAI22DL port map( A1 => mult_28_C96_n781, A2 => 
                           mult_28_C96_n6, B1 => mult_28_C96_n780, B2 => 
                           mult_28_C96_n824, Z => mult_28_C96_n646);
   mult_28_C96_U782 : ADFULD2 port map( A => mult_28_C96_n397, B => 
                           mult_28_C96_n571, CI => mult_28_C96_n556, CO => 
                           mult_28_C96_n383, S => mult_28_C96_n384);
   mult_28_C96_U781 : EXNOR2DL port map( A1 => y_6_port, A2 => 
                           coeff_memory_15_port, Z => mult_28_C96_n658);
   mult_28_C96_U780 : INVD1 port map( A => mult_28_C96_n904, Z => 
                           mult_28_C96_n905);
   mult_28_C96_U779 : INVDL port map( A => mult_28_C96_n605, Z => 
                           mult_28_C96_n904);
   mult_28_C96_U778 : INVBD32 port map( A => mult_28_C96_n24, Z => 
                           mult_28_C96_n903);
   mult_28_C96_U777 : EXOR2D2 port map( A1 => mult_28_C96_n1037, A2 => 
                           mult_28_C96_n423, Z => mult_28_C96_n966);
   mult_28_C96_U776 : EXNOR2DL port map( A1 => y_8_port, A2 => 
                           coeff_memory_9_port, Z => mult_28_C96_n908);
   mult_28_C96_U775 : OAI22D1 port map( A1 => mult_28_C96_n754, A2 => 
                           mult_28_C96_n12, B1 => mult_28_C96_n753, B2 => 
                           mult_28_C96_n9, Z => mult_28_C96_n902);
   mult_28_C96_U774 : EXNOR2D2 port map( A1 => y_11_port, A2 => 
                           coeff_memory_5_port, Z => mult_28_C96_n738);
   mult_28_C96_U773 : OAI22DL port map( A1 => mult_28_C96_n18, A2 => 
                           mult_28_C96_n1060, B1 => mult_28_C96_n738, B2 => 
                           mult_28_C96_n16, Z => mult_28_C96_n604);
   mult_28_C96_U772 : OAI22D1 port map( A1 => mult_28_C96_n18, A2 => 
                           mult_28_C96_n1060, B1 => mult_28_C96_n738, B2 => 
                           mult_28_C96_n16, Z => mult_28_C96_n901);
   mult_28_C96_U771 : EXOR2D1 port map( A1 => mult_28_C96_n1037, A2 => 
                           mult_28_C96_n423, Z => mult_28_C96_n406);
   mult_28_C96_U770 : INVBD32 port map( A => mult_28_C96_n903, Z => 
                           mult_28_C96_n900);
   mult_28_C96_U769 : OAI22D1 port map( A1 => mult_28_C96_n900, A2 => 
                           mult_28_C96_n721, B1 => mult_28_C96_n720, B2 => 
                           mult_28_C96_n22, Z => mult_28_C96_n586);
   mult_28_C96_U768 : NAN2D1 port map( A1 => mult_28_C96_n454, A2 => 
                           mult_28_C96_n463, Z => mult_28_C96_n223);
   mult_28_C96_U767 : OAI22D2 port map( A1 => mult_28_C96_n735, A2 => 
                           mult_28_C96_n18, B1 => mult_28_C96_n734, B2 => 
                           mult_28_C96_n16, Z => mult_28_C96_n600);
   mult_28_C96_U763 : EXOR2D1 port map( A1 => coeff_memory_1_port, A2 => 
                           coeff_memory_0_port, Z => mult_28_C96_n808);
   mult_28_C96_U760 : EXOR2D1 port map( A1 => coeff_memory_3_port, A2 => 
                           coeff_memory_2_port, Z => mult_28_C96_n807);
   mult_28_C96_U757 : EXOR2D1 port map( A1 => coeff_memory_5_port, A2 => 
                           coeff_memory_4_port, Z => mult_28_C96_n806);
   mult_28_C96_U754 : EXOR2D1 port map( A1 => coeff_memory_7_port, A2 => 
                           coeff_memory_6_port, Z => mult_28_C96_n805);
   mult_28_C96_U751 : EXOR2D1 port map( A1 => coeff_memory_9_port, A2 => 
                           coeff_memory_8_port, Z => mult_28_C96_n804);
   mult_28_C96_U748 : EXOR2D1 port map( A1 => coeff_memory_11_port, A2 => 
                           coeff_memory_10_port, Z => mult_28_C96_n803);
   mult_28_C96_U745 : EXOR2D1 port map( A1 => coeff_memory_13_port, A2 => 
                           coeff_memory_12_port, Z => mult_28_C96_n802);
   mult_28_C96_U742 : EXOR2D1 port map( A1 => coeff_memory_15_port, A2 => 
                           coeff_memory_14_port, Z => mult_28_C96_n801);
   mult_28_C96_U717 : NAN2M1D1 port map( A1 => n39, A2 => coeff_memory_1_port, 
                           Z => mult_28_C96_n784);
   mult_28_C96_U716 : EXNOR2D1 port map( A1 => n39, A2 => coeff_memory_1_port, 
                           Z => mult_28_C96_n783);
   mult_28_C96_U712 : EXNOR2D1 port map( A1 => y_4_port, A2 => 
                           coeff_memory_1_port, Z => mult_28_C96_n779);
   mult_28_C96_U699 : OAI22D1 port map( A1 => mult_28_C96_n783, A2 => 
                           mult_28_C96_n6, B1 => mult_28_C96_n782, B2 => 
                           mult_28_C96_n824, Z => mult_28_C96_n648);
   mult_28_C96_U698 : OAI22D1 port map( A1 => mult_28_C96_n782, A2 => 
                           mult_28_C96_n6, B1 => mult_28_C96_n781, B2 => 
                           mult_28_C96_n824, Z => mult_28_C96_n647);
   mult_28_C96_U696 : OAI22D1 port map( A1 => mult_28_C96_n780, A2 => 
                           mult_28_C96_n6, B1 => mult_28_C96_n779, B2 => 
                           mult_28_C96_n824, Z => mult_28_C96_n645);
   mult_28_C96_U695 : OAI22D1 port map( A1 => mult_28_C96_n779, A2 => 
                           mult_28_C96_n6, B1 => mult_28_C96_n778, B2 => 
                           mult_28_C96_n824, Z => mult_28_C96_n644);
   mult_28_C96_U694 : OAI22D1 port map( A1 => mult_28_C96_n778, A2 => 
                           mult_28_C96_n6, B1 => mult_28_C96_n777, B2 => 
                           mult_28_C96_n824, Z => mult_28_C96_n643);
   mult_28_C96_U693 : OAI22D1 port map( A1 => mult_28_C96_n777, A2 => 
                           mult_28_C96_n6, B1 => mult_28_C96_n776, B2 => 
                           mult_28_C96_n824, Z => mult_28_C96_n642);
   mult_28_C96_U692 : OAI22D1 port map( A1 => mult_28_C96_n776, A2 => 
                           mult_28_C96_n6, B1 => mult_28_C96_n775, B2 => 
                           mult_28_C96_n824, Z => mult_28_C96_n641);
   mult_28_C96_U690 : OAI22D1 port map( A1 => mult_28_C96_n773, A2 => 
                           mult_28_C96_n824, B1 => mult_28_C96_n774, B2 => 
                           mult_28_C96_n6, Z => mult_28_C96_n639);
   mult_28_C96_U688 : OAI22D1 port map( A1 => mult_28_C96_n772, A2 => 
                           mult_28_C96_n6, B1 => mult_28_C96_n771, B2 => 
                           mult_28_C96_n824, Z => mult_28_C96_n637);
   mult_28_C96_U683 : OAI22D1 port map( A1 => mult_28_C96_n6, A2 => 
                           mult_28_C96_n832, B1 => mult_28_C96_n784, B2 => 
                           mult_28_C96_n824, Z => mult_28_C96_n520);
   mult_28_C96_U682 : NAN2M1D1 port map( A1 => n39, A2 => coeff_memory_3_port, 
                           Z => mult_28_C96_n767);
   mult_28_C96_U681 : EXNOR2D1 port map( A1 => n39, A2 => coeff_memory_3_port, 
                           Z => mult_28_C96_n766);
   mult_28_C96_U677 : EXNOR2D1 port map( A1 => y_4_port, A2 => 
                           coeff_memory_3_port, Z => mult_28_C96_n762);
   mult_28_C96_U666 : EXNOR2D1 port map( A1 => y_15_port, A2 => 
                           coeff_memory_3_port, Z => mult_28_C96_n751);
   mult_28_C96_U665 : NOR2M1D1 port map( A1 => n39, A2 => mult_28_C96_n9, Z => 
                           mult_28_C96_n632);
   mult_28_C96_U664 : OAI22D1 port map( A1 => mult_28_C96_n766, A2 => 
                           mult_28_C96_n12, B1 => mult_28_C96_n765, B2 => 
                           mult_28_C96_n9, Z => mult_28_C96_n631);
   mult_28_C96_U663 : OAI22D1 port map( A1 => mult_28_C96_n765, A2 => 
                           mult_28_C96_n12, B1 => mult_28_C96_n764, B2 => 
                           mult_28_C96_n9, Z => mult_28_C96_n630);
   mult_28_C96_U662 : OAI22D1 port map( A1 => mult_28_C96_n764, A2 => 
                           mult_28_C96_n12, B1 => mult_28_C96_n763, B2 => 
                           mult_28_C96_n9, Z => mult_28_C96_n629);
   mult_28_C96_U661 : OAI22D1 port map( A1 => mult_28_C96_n763, A2 => 
                           mult_28_C96_n12, B1 => mult_28_C96_n762, B2 => 
                           mult_28_C96_n9, Z => mult_28_C96_n628);
   mult_28_C96_U660 : OAI22D1 port map( A1 => mult_28_C96_n762, A2 => 
                           mult_28_C96_n12, B1 => mult_28_C96_n761, B2 => 
                           mult_28_C96_n9, Z => mult_28_C96_n627);
   mult_28_C96_U659 : OAI22D1 port map( A1 => mult_28_C96_n761, A2 => 
                           mult_28_C96_n12, B1 => mult_28_C96_n760, B2 => 
                           mult_28_C96_n9, Z => mult_28_C96_n626);
   mult_28_C96_U658 : OAI22D1 port map( A1 => mult_28_C96_n760, A2 => 
                           mult_28_C96_n12, B1 => mult_28_C96_n759, B2 => 
                           mult_28_C96_n9, Z => mult_28_C96_n625);
   mult_28_C96_U657 : OAI22D1 port map( A1 => mult_28_C96_n759, A2 => 
                           mult_28_C96_n12, B1 => mult_28_C96_n758, B2 => 
                           mult_28_C96_n9, Z => mult_28_C96_n624);
   mult_28_C96_U655 : OAI22D1 port map( A1 => mult_28_C96_n756, A2 => 
                           mult_28_C96_n9, B1 => mult_28_C96_n757, B2 => 
                           mult_28_C96_n12, Z => mult_28_C96_n622);
   mult_28_C96_U654 : OAI22D1 port map( A1 => mult_28_C96_n756, A2 => 
                           mult_28_C96_n12, B1 => mult_28_C96_n755, B2 => 
                           mult_28_C96_n9, Z => mult_28_C96_n621);
   mult_28_C96_U653 : OAI22D1 port map( A1 => mult_28_C96_n12, A2 => 
                           mult_28_C96_n755, B1 => mult_28_C96_n754, B2 => 
                           mult_28_C96_n9, Z => mult_28_C96_n620);
   mult_28_C96_U652 : OAI22D1 port map( A1 => mult_28_C96_n754, A2 => 
                           mult_28_C96_n12, B1 => mult_28_C96_n753, B2 => 
                           mult_28_C96_n9, Z => mult_28_C96_n619);
   mult_28_C96_U648 : OAI22D1 port map( A1 => mult_28_C96_n12, A2 => 
                           mult_28_C96_n831, B1 => mult_28_C96_n767, B2 => 
                           mult_28_C96_n9, Z => mult_28_C96_n519);
   mult_28_C96_U647 : NAN2M1D1 port map( A1 => n39, A2 => coeff_memory_5_port, 
                           Z => mult_28_C96_n750);
   mult_28_C96_U646 : EXNOR2D1 port map( A1 => n39, A2 => coeff_memory_5_port, 
                           Z => mult_28_C96_n749);
   mult_28_C96_U642 : EXNOR2D1 port map( A1 => y_4_port, A2 => 
                           coeff_memory_5_port, Z => mult_28_C96_n745);
   mult_28_C96_U630 : NOR2M1D1 port map( A1 => n39, A2 => mult_28_C96_n16, Z =>
                           mult_28_C96_n615);
   mult_28_C96_U629 : OAI22D1 port map( A1 => mult_28_C96_n749, A2 => 
                           mult_28_C96_n18, B1 => mult_28_C96_n748, B2 => 
                           mult_28_C96_n16, Z => mult_28_C96_n614);
   mult_28_C96_U628 : OAI22D1 port map( A1 => mult_28_C96_n748, A2 => 
                           mult_28_C96_n18, B1 => mult_28_C96_n747, B2 => 
                           mult_28_C96_n16, Z => mult_28_C96_n613);
   mult_28_C96_U627 : OAI22D1 port map( A1 => mult_28_C96_n747, A2 => 
                           mult_28_C96_n18, B1 => mult_28_C96_n746, B2 => 
                           mult_28_C96_n16, Z => mult_28_C96_n612);
   mult_28_C96_U626 : OAI22D1 port map( A1 => mult_28_C96_n746, A2 => 
                           mult_28_C96_n18, B1 => mult_28_C96_n745, B2 => 
                           mult_28_C96_n16, Z => mult_28_C96_n611);
   mult_28_C96_U625 : OAI22D1 port map( A1 => mult_28_C96_n745, A2 => 
                           mult_28_C96_n18, B1 => mult_28_C96_n744, B2 => 
                           mult_28_C96_n16, Z => mult_28_C96_n610);
   mult_28_C96_U624 : OAI22D1 port map( A1 => mult_28_C96_n744, A2 => 
                           mult_28_C96_n18, B1 => mult_28_C96_n743, B2 => 
                           mult_28_C96_n16, Z => mult_28_C96_n609);
   mult_28_C96_U623 : OAI22D1 port map( A1 => mult_28_C96_n743, A2 => 
                           mult_28_C96_n18, B1 => mult_28_C96_n742, B2 => 
                           mult_28_C96_n16, Z => mult_28_C96_n608);
   mult_28_C96_U621 : OAI22D1 port map( A1 => mult_28_C96_n741, A2 => 
                           mult_28_C96_n18, B1 => mult_28_C96_n740, B2 => 
                           mult_28_C96_n16, Z => mult_28_C96_n606);
   mult_28_C96_U616 : OAI22D1 port map( A1 => mult_28_C96_n736, A2 => 
                           mult_28_C96_n18, B1 => mult_28_C96_n735, B2 => 
                           mult_28_C96_n16, Z => mult_28_C96_n601);
   mult_28_C96_U613 : OAI22D1 port map( A1 => mult_28_C96_n18, A2 => 
                           mult_28_C96_n830, B1 => mult_28_C96_n750, B2 => 
                           mult_28_C96_n16, Z => mult_28_C96_n518);
   mult_28_C96_U612 : NAN2M1D1 port map( A1 => n39, A2 => coeff_memory_7_port, 
                           Z => mult_28_C96_n733);
   mult_28_C96_U611 : EXNOR2D1 port map( A1 => n39, A2 => coeff_memory_7_port, 
                           Z => mult_28_C96_n732);
   mult_28_C96_U596 : EXNOR2D1 port map( A1 => y_15_port, A2 => 
                           coeff_memory_7_port, Z => mult_28_C96_n717);
   mult_28_C96_U595 : NOR2M1D1 port map( A1 => n39, A2 => mult_28_C96_n22, Z =>
                           mult_28_C96_n598);
   mult_28_C96_U594 : OAI22D1 port map( A1 => mult_28_C96_n732, A2 => 
                           mult_28_C96_n24, B1 => mult_28_C96_n731, B2 => 
                           mult_28_C96_n22, Z => mult_28_C96_n597);
   mult_28_C96_U593 : OAI22D1 port map( A1 => mult_28_C96_n731, A2 => 
                           mult_28_C96_n24, B1 => mult_28_C96_n730, B2 => 
                           mult_28_C96_n22, Z => mult_28_C96_n596);
   mult_28_C96_U592 : OAI22D1 port map( A1 => mult_28_C96_n730, A2 => 
                           mult_28_C96_n24, B1 => mult_28_C96_n729, B2 => 
                           mult_28_C96_n22, Z => mult_28_C96_n595);
   mult_28_C96_U591 : OAI22D1 port map( A1 => mult_28_C96_n729, A2 => 
                           mult_28_C96_n24, B1 => mult_28_C96_n728, B2 => 
                           mult_28_C96_n22, Z => mult_28_C96_n594);
   mult_28_C96_U590 : OAI22D1 port map( A1 => mult_28_C96_n728, A2 => 
                           mult_28_C96_n24, B1 => mult_28_C96_n727, B2 => 
                           mult_28_C96_n22, Z => mult_28_C96_n593);
   mult_28_C96_U589 : OAI22D1 port map( A1 => mult_28_C96_n727, A2 => 
                           mult_28_C96_n24, B1 => mult_28_C96_n726, B2 => 
                           mult_28_C96_n22, Z => mult_28_C96_n592);
   mult_28_C96_U588 : OAI22D1 port map( A1 => mult_28_C96_n726, A2 => 
                           mult_28_C96_n24, B1 => mult_28_C96_n725, B2 => 
                           mult_28_C96_n22, Z => mult_28_C96_n591);
   mult_28_C96_U587 : OAI22D1 port map( A1 => mult_28_C96_n24, A2 => 
                           mult_28_C96_n725, B1 => mult_28_C96_n724, B2 => 
                           mult_28_C96_n22, Z => mult_28_C96_n590);
   mult_28_C96_U586 : OAI22D1 port map( A1 => mult_28_C96_n724, A2 => 
                           mult_28_C96_n24, B1 => mult_28_C96_n723, B2 => 
                           mult_28_C96_n22, Z => mult_28_C96_n589);
   mult_28_C96_U585 : OAI22D1 port map( A1 => mult_28_C96_n722, A2 => 
                           mult_28_C96_n22, B1 => mult_28_C96_n723, B2 => 
                           mult_28_C96_n24, Z => mult_28_C96_n588);
   mult_28_C96_U584 : OAI22D1 port map( A1 => mult_28_C96_n722, A2 => 
                           mult_28_C96_n24, B1 => mult_28_C96_n1002, B2 => 
                           mult_28_C96_n22, Z => mult_28_C96_n587);
   mult_28_C96_U582 : OAI22D1 port map( A1 => mult_28_C96_n720, A2 => 
                           mult_28_C96_n24, B1 => mult_28_C96_n719, B2 => 
                           mult_28_C96_n22, Z => mult_28_C96_n585);
   mult_28_C96_U581 : OAI22D1 port map( A1 => mult_28_C96_n719, A2 => 
                           mult_28_C96_n24, B1 => mult_28_C96_n718, B2 => 
                           mult_28_C96_n22, Z => mult_28_C96_n584);
   mult_28_C96_U579 : AO21D2 port map( A1 => mult_28_C96_n24, A2 => 
                           mult_28_C96_n22, B => mult_28_C96_n717, Z => 
                           mult_28_C96_n582);
   mult_28_C96_U578 : OAI22D1 port map( A1 => mult_28_C96_n24, A2 => 
                           mult_28_C96_n829, B1 => mult_28_C96_n733, B2 => 
                           mult_28_C96_n22, Z => mult_28_C96_n517);
   mult_28_C96_U577 : NAN2M1D1 port map( A1 => n39, A2 => coeff_memory_9_port, 
                           Z => mult_28_C96_n716);
   mult_28_C96_U576 : EXNOR2D1 port map( A1 => n39, A2 => coeff_memory_9_port, 
                           Z => mult_28_C96_n715);
   mult_28_C96_U560 : NOR2M1D1 port map( A1 => n39, A2 => mult_28_C96_n28, Z =>
                           mult_28_C96_n581);
   mult_28_C96_U559 : OAI22D1 port map( A1 => mult_28_C96_n715, A2 => 
                           mult_28_C96_n30, B1 => mult_28_C96_n714, B2 => 
                           mult_28_C96_n28, Z => mult_28_C96_n580);
   mult_28_C96_U558 : OAI22D1 port map( A1 => mult_28_C96_n714, A2 => 
                           mult_28_C96_n30, B1 => mult_28_C96_n713, B2 => 
                           mult_28_C96_n28, Z => mult_28_C96_n579);
   mult_28_C96_U557 : OAI22D1 port map( A1 => mult_28_C96_n713, A2 => 
                           mult_28_C96_n30, B1 => mult_28_C96_n712, B2 => 
                           mult_28_C96_n28, Z => mult_28_C96_n578);
   mult_28_C96_U556 : OAI22D1 port map( A1 => mult_28_C96_n712, A2 => 
                           mult_28_C96_n30, B1 => mult_28_C96_n711, B2 => 
                           mult_28_C96_n28, Z => mult_28_C96_n577);
   mult_28_C96_U555 : OAI22D1 port map( A1 => mult_28_C96_n711, A2 => 
                           mult_28_C96_n30, B1 => mult_28_C96_n710, B2 => 
                           mult_28_C96_n28, Z => mult_28_C96_n576);
   mult_28_C96_U554 : OAI22D1 port map( A1 => mult_28_C96_n710, A2 => 
                           mult_28_C96_n30, B1 => mult_28_C96_n709, B2 => 
                           mult_28_C96_n28, Z => mult_28_C96_n575);
   mult_28_C96_U553 : OAI22D1 port map( A1 => mult_28_C96_n709, A2 => 
                           mult_28_C96_n30, B1 => mult_28_C96_n708, B2 => 
                           mult_28_C96_n28, Z => mult_28_C96_n574);
   mult_28_C96_U551 : OAI22D1 port map( A1 => mult_28_C96_n707, A2 => 
                           mult_28_C96_n30, B1 => mult_28_C96_n706, B2 => 
                           mult_28_C96_n28, Z => mult_28_C96_n572);
   mult_28_C96_U548 : OAI22D1 port map( A1 => mult_28_C96_n704, A2 => 
                           mult_28_C96_n30, B1 => mult_28_C96_n703, B2 => 
                           mult_28_C96_n28, Z => mult_28_C96_n569);
   mult_28_C96_U547 : OAI22D1 port map( A1 => mult_28_C96_n703, A2 => 
                           mult_28_C96_n30, B1 => mult_28_C96_n702, B2 => 
                           mult_28_C96_n28, Z => mult_28_C96_n568);
   mult_28_C96_U546 : OAI22D1 port map( A1 => mult_28_C96_n702, A2 => 
                           mult_28_C96_n30, B1 => mult_28_C96_n701, B2 => 
                           mult_28_C96_n28, Z => mult_28_C96_n567);
   mult_28_C96_U544 : AO21D2 port map( A1 => mult_28_C96_n30, A2 => 
                           mult_28_C96_n28, B => mult_28_C96_n700, Z => 
                           mult_28_C96_n565);
   mult_28_C96_U543 : OAI22D1 port map( A1 => mult_28_C96_n30, A2 => 
                           mult_28_C96_n828, B1 => mult_28_C96_n716, B2 => 
                           mult_28_C96_n28, Z => mult_28_C96_n516);
   mult_28_C96_U542 : NAN2M1D1 port map( A1 => n39, A2 => coeff_memory_11_port,
                           Z => mult_28_C96_n699);
   mult_28_C96_U541 : EXNOR2D1 port map( A1 => n39, A2 => coeff_memory_11_port,
                           Z => mult_28_C96_n698);
   mult_28_C96_U525 : NOR2M1D1 port map( A1 => n39, A2 => mult_28_C96_n34, Z =>
                           mult_28_C96_n564);
   mult_28_C96_U524 : OAI22D1 port map( A1 => mult_28_C96_n698, A2 => 
                           mult_28_C96_n36, B1 => mult_28_C96_n697, B2 => 
                           mult_28_C96_n34, Z => mult_28_C96_n563);
   mult_28_C96_U523 : OAI22D1 port map( A1 => mult_28_C96_n697, A2 => 
                           mult_28_C96_n36, B1 => mult_28_C96_n696, B2 => 
                           mult_28_C96_n34, Z => mult_28_C96_n562);
   mult_28_C96_U522 : OAI22D1 port map( A1 => mult_28_C96_n696, A2 => 
                           mult_28_C96_n36, B1 => mult_28_C96_n695, B2 => 
                           mult_28_C96_n34, Z => mult_28_C96_n561);
   mult_28_C96_U521 : OAI22D1 port map( A1 => mult_28_C96_n695, A2 => 
                           mult_28_C96_n36, B1 => mult_28_C96_n694, B2 => 
                           mult_28_C96_n34, Z => mult_28_C96_n560);
   mult_28_C96_U520 : OAI22D1 port map( A1 => mult_28_C96_n694, A2 => 
                           mult_28_C96_n36, B1 => mult_28_C96_n693, B2 => 
                           mult_28_C96_n34, Z => mult_28_C96_n559);
   mult_28_C96_U519 : OAI22D1 port map( A1 => mult_28_C96_n693, A2 => 
                           mult_28_C96_n36, B1 => mult_28_C96_n692, B2 => 
                           mult_28_C96_n34, Z => mult_28_C96_n558);
   mult_28_C96_U518 : OAI22D1 port map( A1 => mult_28_C96_n692, A2 => 
                           mult_28_C96_n36, B1 => mult_28_C96_n691, B2 => 
                           mult_28_C96_n34, Z => mult_28_C96_n557);
   mult_28_C96_U516 : OAI22D1 port map( A1 => mult_28_C96_n690, A2 => 
                           mult_28_C96_n36, B1 => mult_28_C96_n689, B2 => 
                           mult_28_C96_n34, Z => mult_28_C96_n555);
   mult_28_C96_U515 : OAI22D1 port map( A1 => mult_28_C96_n688, A2 => 
                           mult_28_C96_n34, B1 => mult_28_C96_n689, B2 => 
                           mult_28_C96_n36, Z => mult_28_C96_n554);
   mult_28_C96_U513 : OAI22D1 port map( A1 => mult_28_C96_n687, A2 => 
                           mult_28_C96_n36, B1 => mult_28_C96_n686, B2 => 
                           mult_28_C96_n34, Z => mult_28_C96_n552);
   mult_28_C96_U511 : OAI22D1 port map( A1 => mult_28_C96_n685, A2 => 
                           mult_28_C96_n36, B1 => mult_28_C96_n684, B2 => 
                           mult_28_C96_n34, Z => mult_28_C96_n550);
   mult_28_C96_U508 : OAI22D1 port map( A1 => mult_28_C96_n36, A2 => 
                           mult_28_C96_n827, B1 => mult_28_C96_n699, B2 => 
                           mult_28_C96_n34, Z => mult_28_C96_n515);
   mult_28_C96_U507 : NAN2M1D1 port map( A1 => n39, A2 => coeff_memory_13_port,
                           Z => mult_28_C96_n682);
   mult_28_C96_U506 : EXNOR2D1 port map( A1 => n39, A2 => coeff_memory_13_port,
                           Z => mult_28_C96_n681);
   mult_28_C96_U490 : NOR2M1D1 port map( A1 => n39, A2 => mult_28_C96_n40, Z =>
                           mult_28_C96_n547);
   mult_28_C96_U489 : OAI22D1 port map( A1 => mult_28_C96_n681, A2 => 
                           mult_28_C96_n42, B1 => mult_28_C96_n680, B2 => 
                           mult_28_C96_n40, Z => mult_28_C96_n546);
   mult_28_C96_U488 : OAI22D1 port map( A1 => mult_28_C96_n994, A2 => 
                           mult_28_C96_n42, B1 => mult_28_C96_n679, B2 => 
                           mult_28_C96_n40, Z => mult_28_C96_n545);
   mult_28_C96_U487 : OAI22D1 port map( A1 => mult_28_C96_n679, A2 => 
                           mult_28_C96_n42, B1 => mult_28_C96_n678, B2 => 
                           mult_28_C96_n40, Z => mult_28_C96_n544);
   mult_28_C96_U486 : OAI22D1 port map( A1 => mult_28_C96_n678, A2 => 
                           mult_28_C96_n42, B1 => mult_28_C96_n677, B2 => 
                           mult_28_C96_n40, Z => mult_28_C96_n543);
   mult_28_C96_U485 : OAI22D1 port map( A1 => mult_28_C96_n677, A2 => 
                           mult_28_C96_n42, B1 => mult_28_C96_n676, B2 => 
                           mult_28_C96_n40, Z => mult_28_C96_n542);
   mult_28_C96_U483 : OAI22D1 port map( A1 => mult_28_C96_n675, A2 => 
                           mult_28_C96_n42, B1 => mult_28_C96_n674, B2 => 
                           mult_28_C96_n40, Z => mult_28_C96_n540);
   mult_28_C96_U481 : OAI22D1 port map( A1 => mult_28_C96_n673, A2 => 
                           mult_28_C96_n42, B1 => mult_28_C96_n672, B2 => 
                           mult_28_C96_n40, Z => mult_28_C96_n538);
   mult_28_C96_U480 : OAI22D1 port map( A1 => mult_28_C96_n671, A2 => 
                           mult_28_C96_n40, B1 => mult_28_C96_n672, B2 => 
                           mult_28_C96_n42, Z => mult_28_C96_n537);
   mult_28_C96_U479 : OAI22D1 port map( A1 => mult_28_C96_n671, A2 => 
                           mult_28_C96_n42, B1 => mult_28_C96_n670, B2 => 
                           mult_28_C96_n40, Z => mult_28_C96_n536);
   mult_28_C96_U478 : OAI22D1 port map( A1 => mult_28_C96_n670, A2 => 
                           mult_28_C96_n42, B1 => mult_28_C96_n669, B2 => 
                           mult_28_C96_n40, Z => mult_28_C96_n535);
   mult_28_C96_U477 : OAI22D1 port map( A1 => mult_28_C96_n669, A2 => 
                           mult_28_C96_n42, B1 => mult_28_C96_n668, B2 => 
                           mult_28_C96_n40, Z => mult_28_C96_n534);
   mult_28_C96_U476 : OAI22D1 port map( A1 => mult_28_C96_n668, A2 => 
                           mult_28_C96_n42, B1 => mult_28_C96_n667, B2 => 
                           mult_28_C96_n40, Z => mult_28_C96_n533);
   mult_28_C96_U475 : OAI22D1 port map( A1 => mult_28_C96_n667, A2 => 
                           mult_28_C96_n42, B1 => mult_28_C96_n666, B2 => 
                           mult_28_C96_n40, Z => mult_28_C96_n309);
   mult_28_C96_U473 : OAI22D1 port map( A1 => mult_28_C96_n42, A2 => 
                           mult_28_C96_n826, B1 => mult_28_C96_n682, B2 => 
                           mult_28_C96_n40, Z => mult_28_C96_n514);
   mult_28_C96_U472 : NAN2M1D1 port map( A1 => n39, A2 => coeff_memory_15_port,
                           Z => mult_28_C96_n665);
   mult_28_C96_U471 : EXNOR2D1 port map( A1 => n39, A2 => coeff_memory_15_port,
                           Z => mult_28_C96_n664);
   mult_28_C96_U455 : NOR2M1D1 port map( A1 => n39, A2 => mult_28_C96_n46, Z =>
                           mult_28_C96_n531);
   mult_28_C96_U454 : OAI22D1 port map( A1 => mult_28_C96_n664, A2 => 
                           mult_28_C96_n48, B1 => mult_28_C96_n663, B2 => 
                           mult_28_C96_n46, Z => mult_28_C96_n530);
   mult_28_C96_U453 : OAI22D1 port map( A1 => mult_28_C96_n916, A2 => 
                           mult_28_C96_n48, B1 => mult_28_C96_n662, B2 => 
                           mult_28_C96_n46, Z => mult_28_C96_n529);
   mult_28_C96_U452 : OAI22D1 port map( A1 => mult_28_C96_n662, A2 => 
                           mult_28_C96_n48, B1 => mult_28_C96_n661, B2 => 
                           mult_28_C96_n46, Z => mult_28_C96_n399);
   mult_28_C96_U451 : OAI22D1 port map( A1 => mult_28_C96_n661, A2 => 
                           mult_28_C96_n48, B1 => mult_28_C96_n660, B2 => 
                           mult_28_C96_n46, Z => mult_28_C96_n528);
   mult_28_C96_U450 : OAI22D1 port map( A1 => mult_28_C96_n660, A2 => 
                           mult_28_C96_n48, B1 => mult_28_C96_n659, B2 => 
                           mult_28_C96_n46, Z => mult_28_C96_n373);
   mult_28_C96_U449 : OAI22D1 port map( A1 => mult_28_C96_n659, A2 => 
                           mult_28_C96_n48, B1 => mult_28_C96_n658, B2 => 
                           mult_28_C96_n46, Z => mult_28_C96_n527);
   mult_28_C96_U448 : OAI22D1 port map( A1 => mult_28_C96_n658, A2 => 
                           mult_28_C96_n48, B1 => mult_28_C96_n657, B2 => 
                           mult_28_C96_n46, Z => mult_28_C96_n351);
   mult_28_C96_U447 : OAI22D1 port map( A1 => mult_28_C96_n657, A2 => 
                           mult_28_C96_n48, B1 => mult_28_C96_n656, B2 => 
                           mult_28_C96_n46, Z => mult_28_C96_n526);
   mult_28_C96_U444 : OAI22D1 port map( A1 => mult_28_C96_n654, A2 => 
                           mult_28_C96_n48, B1 => mult_28_C96_n653, B2 => 
                           mult_28_C96_n46, Z => mult_28_C96_n319);
   mult_28_C96_U441 : OAI22D1 port map( A1 => mult_28_C96_n651, A2 => 
                           mult_28_C96_n48, B1 => mult_28_C96_n650, B2 => 
                           mult_28_C96_n46, Z => mult_28_C96_n522);
   mult_28_C96_U439 : OAI22D1 port map( A1 => mult_28_C96_n48, A2 => 
                           mult_28_C96_n825, B1 => mult_28_C96_n665, B2 => 
                           mult_28_C96_n46, Z => mult_28_C96_n513);
   mult_28_C96_U437 : ADFULD1 port map( A => mult_28_C96_n511, B => 
                           mult_28_C96_n615, CI => mult_28_C96_n630, CO => 
                           mult_28_C96_n509, S => mult_28_C96_n510);
   mult_28_C96_U436 : ADHALFD1 port map( A => mult_28_C96_n614, B => 
                           mult_28_C96_n518, CO => mult_28_C96_n507, S => 
                           mult_28_C96_n508);
   mult_28_C96_U435 : ADFULD1 port map( A => mult_28_C96_n629, B => 
                           mult_28_C96_n508, CI => mult_28_C96_n644, CO => 
                           mult_28_C96_n505, S => mult_28_C96_n506);
   mult_28_C96_U434 : ADFULD1 port map( A => mult_28_C96_n507, B => 
                           mult_28_C96_n598, CI => mult_28_C96_n613, CO => 
                           mult_28_C96_n503, S => mult_28_C96_n504);
   mult_28_C96_U433 : ADFULD1 port map( A => mult_28_C96_n643, B => 
                           mult_28_C96_n628, CI => mult_28_C96_n504, CO => 
                           mult_28_C96_n501, S => mult_28_C96_n502);
   mult_28_C96_U432 : ADHALFD1 port map( A => mult_28_C96_n597, B => 
                           mult_28_C96_n517, CO => mult_28_C96_n499, S => 
                           mult_28_C96_n500);
   mult_28_C96_U431 : ADFULD1 port map( A => mult_28_C96_n612, B => 
                           mult_28_C96_n500, CI => mult_28_C96_n627, CO => 
                           mult_28_C96_n497, S => mult_28_C96_n498);
   mult_28_C96_U430 : ADFULD1 port map( A => mult_28_C96_n642, B => 
                           mult_28_C96_n503, CI => mult_28_C96_n498, CO => 
                           mult_28_C96_n495, S => mult_28_C96_n496);
   mult_28_C96_U429 : ADFULD1 port map( A => mult_28_C96_n499, B => 
                           mult_28_C96_n581, CI => mult_28_C96_n596, CO => 
                           mult_28_C96_n493, S => mult_28_C96_n494);
   mult_28_C96_U428 : ADFULD1 port map( A => mult_28_C96_n626, B => 
                           mult_28_C96_n611, CI => mult_28_C96_n494, CO => 
                           mult_28_C96_n491, S => mult_28_C96_n492);
   mult_28_C96_U427 : ADFULD1 port map( A => mult_28_C96_n641, B => 
                           mult_28_C96_n497, CI => mult_28_C96_n492, CO => 
                           mult_28_C96_n489, S => mult_28_C96_n490);
   mult_28_C96_U426 : ADHALFD1 port map( A => mult_28_C96_n580, B => 
                           mult_28_C96_n516, CO => mult_28_C96_n487, S => 
                           mult_28_C96_n488);
   mult_28_C96_U425 : ADFULD1 port map( A => mult_28_C96_n595, B => 
                           mult_28_C96_n488, CI => mult_28_C96_n610, CO => 
                           mult_28_C96_n485, S => mult_28_C96_n486);
   mult_28_C96_U422 : ADFULD1 port map( A => mult_28_C96_n487, B => 
                           mult_28_C96_n564, CI => mult_28_C96_n579, CO => 
                           mult_28_C96_n479, S => mult_28_C96_n480);
   mult_28_C96_U421 : ADFULD1 port map( A => mult_28_C96_n609, B => 
                           mult_28_C96_n594, CI => mult_28_C96_n480, CO => 
                           mult_28_C96_n477, S => mult_28_C96_n478);
   mult_28_C96_U420 : ADFULD1 port map( A => mult_28_C96_n639, B => 
                           mult_28_C96_n485, CI => mult_28_C96_n624, CO => 
                           mult_28_C96_n475, S => mult_28_C96_n476);
   mult_28_C96_U419 : ADFULD1 port map( A => mult_28_C96_n483, B => 
                           mult_28_C96_n478, CI => mult_28_C96_n476, CO => 
                           mult_28_C96_n473, S => mult_28_C96_n474);
   mult_28_C96_U417 : ADFULD1 port map( A => mult_28_C96_n578, B => 
                           mult_28_C96_n472, CI => mult_28_C96_n593, CO => 
                           mult_28_C96_n469, S => mult_28_C96_n470);
   mult_28_C96_U416 : ADFULD1 port map( A => mult_28_C96_n608, B => 
                           mult_28_C96_n479, CI => mult_28_C96_n623, CO => 
                           mult_28_C96_n467, S => mult_28_C96_n468);
   mult_28_C96_U415 : ADFULD1 port map( A => mult_28_C96_n470, B => 
                           mult_28_C96_n638, CI => mult_28_C96_n477, CO => 
                           mult_28_C96_n465, S => mult_28_C96_n466);
   mult_28_C96_U414 : ADFULD1 port map( A => mult_28_C96_n468, B => 
                           mult_28_C96_n475, CI => mult_28_C96_n466, CO => 
                           mult_28_C96_n463, S => mult_28_C96_n464);
   mult_28_C96_U413 : ADFULD1 port map( A => mult_28_C96_n471, B => 
                           mult_28_C96_n547, CI => mult_28_C96_n562, CO => 
                           mult_28_C96_n461, S => mult_28_C96_n462);
   mult_28_C96_U412 : ADFULD1 port map( A => mult_28_C96_n592, B => 
                           mult_28_C96_n577, CI => mult_28_C96_n462, CO => 
                           mult_28_C96_n459, S => mult_28_C96_n460);
   mult_28_C96_U410 : ADFULD1 port map( A => mult_28_C96_n460, B => 
                           mult_28_C96_n637, CI => mult_28_C96_n467, CO => 
                           mult_28_C96_n455, S => mult_28_C96_n456);
   mult_28_C96_U409 : ADFULD1 port map( A => mult_28_C96_n458, B => 
                           mult_28_C96_n465, CI => mult_28_C96_n456, CO => 
                           mult_28_C96_n453, S => mult_28_C96_n454);
   mult_28_C96_U404 : ADFULD1 port map( A => mult_28_C96_n457, B => 
                           mult_28_C96_n459, CI => mult_28_C96_n448, CO => 
                           mult_28_C96_n443, S => mult_28_C96_n444);
   mult_28_C96_U402 : ADFULD1 port map( A => mult_28_C96_n451, B => 
                           mult_28_C96_n531, CI => mult_28_C96_n545, CO => 
                           mult_28_C96_n439, S => mult_28_C96_n440);
   mult_28_C96_U398 : ADFULD1 port map( A => mult_28_C96_n445, B => 
                           mult_28_C96_n447, CI => mult_28_C96_n436, CO => 
                           mult_28_C96_n431, S => mult_28_C96_n432);
   mult_28_C96_U391 : ADFULD1 port map( A => mult_28_C96_n433, B => 
                           mult_28_C96_n424, CI => mult_28_C96_n422, CO => 
                           mult_28_C96_n417, S => mult_28_C96_n418);
   mult_28_C96_U387 : ADFULD1 port map( A => mult_28_C96_n414, B => 
                           mult_28_C96_n543, CI => mult_28_C96_n558, CO => 
                           mult_28_C96_n411, S => mult_28_C96_n412);
   mult_28_C96_U385 : ADFULD1 port map( A => mult_28_C96_n618, B => 
                           mult_28_C96_n603, CI => mult_28_C96_n412, CO => 
                           mult_28_C96_n407, S => mult_28_C96_n408);
   mult_28_C96_U382 : ADFULD1 port map( A => mult_28_C96_n417, B => 
                           mult_28_C96_n966, CI => mult_28_C96_n404, CO => 
                           mult_28_C96_n401, S => mult_28_C96_n402);
   mult_28_C96_U380 : ADFULD1 port map( A => mult_28_C96_n413, B => 
                           mult_28_C96_n400, CI => mult_28_C96_n542, CO => 
                           mult_28_C96_n397, S => mult_28_C96_n398);
   mult_28_C96_U379 : ADFULD1 port map( A => mult_28_C96_n572, B => 
                           mult_28_C96_n557, CI => mult_28_C96_n411, CO => 
                           mult_28_C96_n395, S => mult_28_C96_n396);
   mult_28_C96_U376 : ADFULD1 port map( A => mult_28_C96_n394, B => 
                           mult_28_C96_n407, CI => mult_28_C96_n405, CO => 
                           mult_28_C96_n389, S => mult_28_C96_n390);
   mult_28_C96_U372 : ADFULD1 port map( A => mult_28_C96_n601, B => 
                           mult_28_C96_n586, CI => mult_28_C96_n386, CO => 
                           mult_28_C96_n381, S => mult_28_C96_n382);
   mult_28_C96_U367 : ADFULD1 port map( A => mult_28_C96_n540, B => 
                           mult_28_C96_n374, CI => mult_28_C96_n555, CO => 
                           mult_28_C96_n371, S => mult_28_C96_n372);
   mult_28_C96_U365 : ADFULD1 port map( A => mult_28_C96_n383, B => 
                           mult_28_C96_n585, CI => mult_28_C96_n372, CO => 
                           mult_28_C96_n367, S => mult_28_C96_n368);
   mult_28_C96_U364 : ADFULD1 port map( A => mult_28_C96_n381, B => 
                           mult_28_C96_n370, CI => mult_28_C96_n379, CO => 
                           mult_28_C96_n365, S => mult_28_C96_n366);
   mult_28_C96_U363 : ADFULD1 port map( A => mult_28_C96_n377, B => 
                           mult_28_C96_n368, CI => mult_28_C96_n366, CO => 
                           mult_28_C96_n363, S => mult_28_C96_n364);
   mult_28_C96_U362 : ADFULD1 port map( A => mult_28_C96_n527, B => 
                           mult_28_C96_n373, CI => mult_28_C96_n554, CO => 
                           mult_28_C96_n361, S => mult_28_C96_n_1016);
   mult_28_C96_U359 : ADFULD1 port map( A => mult_28_C96_n360, B => 
                           mult_28_C96_n369, CI => mult_28_C96_n367, CO => 
                           mult_28_C96_n355, S => mult_28_C96_n356);
   mult_28_C96_U356 : ADFULD1 port map( A => mult_28_C96_n352, B => 
                           mult_28_C96_n538, CI => mult_28_C96_n553, CO => 
                           mult_28_C96_n349, S => mult_28_C96_n350);
   mult_28_C96_U355 : ADFULD1 port map( A => mult_28_C96_n583, B => 
                           mult_28_C96_n568, CI => mult_28_C96_n361, CO => 
                           mult_28_C96_n347, S => mult_28_C96_n348);
   mult_28_C96_U354 : ADFULD1 port map( A => mult_28_C96_n350, B => 
                           mult_28_C96_n359, CI => mult_28_C96_n357, CO => 
                           mult_28_C96_n345, S => mult_28_C96_n346);
   mult_28_C96_U353 : ADFULD1 port map( A => mult_28_C96_n355, B => 
                           mult_28_C96_n348, CI => mult_28_C96_n346, CO => 
                           mult_28_C96_n343, S => mult_28_C96_n344);
   mult_28_C96_U352 : ADFULD1 port map( A => mult_28_C96_n537, B => 
                           mult_28_C96_n351, CI => mult_28_C96_n526, CO => 
                           mult_28_C96_n341, S => mult_28_C96_n342);
   mult_28_C96_U351 : ADFULD1 port map( A => mult_28_C96_n567, B => 
                           mult_28_C96_n552, CI => mult_28_C96_n582, CO => 
                           mult_28_C96_n339, S => mult_28_C96_n340);
   mult_28_C96_U350 : ADFULD1 port map( A => mult_28_C96_n342, B => 
                           mult_28_C96_n349, CI => mult_28_C96_n347, CO => 
                           mult_28_C96_n337, S => mult_28_C96_n338);
   mult_28_C96_U349 : ADFULD1 port map( A => mult_28_C96_n345, B => 
                           mult_28_C96_n340, CI => mult_28_C96_n338, CO => 
                           mult_28_C96_n335, S => mult_28_C96_n336);
   mult_28_C96_U347 : ADFULD1 port map( A => mult_28_C96_n536, B => 
                           mult_28_C96_n334, CI => mult_28_C96_n551, CO => 
                           mult_28_C96_n331, S => mult_28_C96_n332);
   mult_28_C96_U345 : ADFULD1 port map( A => mult_28_C96_n337, B => 
                           mult_28_C96_n332, CI => mult_28_C96_n330, CO => 
                           mult_28_C96_n327, S => mult_28_C96_n328);
   mult_28_C96_U343 : ADFULD1 port map( A => mult_28_C96_n565, B => 
                           mult_28_C96_n535, CI => mult_28_C96_n331, CO => 
                           mult_28_C96_n323, S => mult_28_C96_n324);
   mult_28_C96_U342 : ADFULD1 port map( A => mult_28_C96_n329, B => 
                           mult_28_C96_n326, CI => mult_28_C96_n324, CO => 
                           mult_28_C96_n321, S => mult_28_C96_n322);
   mult_28_C96_U340 : ADFULD1 port map( A => mult_28_C96_n534, B => 
                           mult_28_C96_n320, CI => mult_28_C96_n549, CO => 
                           mult_28_C96_n317, S => mult_28_C96_n318);
   mult_28_C96_U339 : ADFULD1 port map( A => mult_28_C96_n318, B => 
                           mult_28_C96_n325, CI => mult_28_C96_n323, CO => 
                           mult_28_C96_n315, S => mult_28_C96_n316);
   mult_28_C96_U338 : ADFULD1 port map( A => mult_28_C96_n524, B => 
                           mult_28_C96_n319, CI => mult_28_C96_n548, CO => 
                           mult_28_C96_n313, S => mult_28_C96_n314);
   mult_28_C96_U337 : ADFULD1 port map( A => mult_28_C96_n317, B => 
                           mult_28_C96_n533, CI => mult_28_C96_n314, CO => 
                           mult_28_C96_n311, S => mult_28_C96_n312);
   mult_28_C96_U335 : ADFULD1 port map( A => mult_28_C96_n310, B => 
                           mult_28_C96_n523, CI => mult_28_C96_n313, CO => 
                           mult_28_C96_n307, S => mult_28_C96_n308);
   mult_28_C96_U334 : ADFULD1 port map( A => mult_28_C96_n522, B => 
                           mult_28_C96_n309, CI => mult_28_C96_n532, CO => 
                           mult_28_C96_n305, S => mult_28_C96_n306);
   mult_28_C96_U320 : AOI21D1 port map( A1 => mult_28_C96_n1088, A2 => 
                           mult_28_C96_n1090, B => mult_28_C96_n1089, Z => 
                           mult_28_C96_n267);
   mult_28_C96_U314 : OAI21D1 port map( A1 => mult_28_C96_n267, A2 => 
                           mult_28_C96_n265, B => mult_28_C96_n266, Z => 
                           mult_28_C96_n264);
   mult_28_C96_U306 : AOI21D1 port map( A1 => mult_28_C96_n1086, A2 => 
                           mult_28_C96_n264, B => mult_28_C96_n1087, Z => 
                           mult_28_C96_n259);
   mult_28_C96_U300 : OAI21D1 port map( A1 => mult_28_C96_n257, A2 => 
                           mult_28_C96_n259, B => mult_28_C96_n258, Z => 
                           mult_28_C96_n256);
   mult_28_C96_U292 : AOI21D1 port map( A1 => mult_28_C96_n256, A2 => 
                           mult_28_C96_n1084, B => mult_28_C96_n1085, Z => 
                           mult_28_C96_n251);
   mult_28_C96_U286 : OAI21D1 port map( A1 => mult_28_C96_n249, A2 => 
                           mult_28_C96_n251, B => mult_28_C96_n250, Z => 
                           mult_28_C96_n248);
   mult_28_C96_U278 : AOI21D1 port map( A1 => mult_28_C96_n248, A2 => 
                           mult_28_C96_n1071, B => mult_28_C96_n1083, Z => 
                           mult_28_C96_n243);
   mult_28_C96_U232 : OAI21D1 port map( A1 => mult_28_C96_n225, A2 => 
                           mult_28_C96_n213, B => mult_28_C96_n214, Z => 
                           mult_28_C96_n212);
   mult_28_C96_U217 : AOI21D1 port map( A1 => mult_28_C96_n204, A2 => 
                           mult_28_C96_n212, B => mult_28_C96_n205, Z => 
                           mult_28_C96_n203);
   mult_28_C96_U207 : EXNOR2D1 port map( A1 => mult_28_C96_n202, A2 => 
                           mult_28_C96_n67, Z => m5_2);
   mult_28_C96_U202 : OAI21D1 port map( A1 => mult_28_C96_n201, A2 => 
                           mult_28_C96_n195, B => mult_28_C96_n196, Z => 
                           mult_28_C96_n190);
   mult_28_C96_U193 : NOR2D2 port map( A1 => mult_28_C96_n376, A2 => 
                           mult_28_C96_n387, Z => mult_28_C96_n184);
   mult_28_C96_U183 : NOR2D2 port map( A1 => mult_28_C96_n364, A2 => 
                           mult_28_C96_n375, Z => mult_28_C96_n179);
   mult_28_C96_U178 : AOI21D1 port map( A1 => mult_28_C96_n177, A2 => 
                           mult_28_C96_n190, B => mult_28_C96_n178, Z => 
                           mult_28_C96_n176);
   mult_28_C96_U168 : AOI21D1 port map( A1 => mult_28_C96_n1020, A2 => 
                           mult_28_C96_n284, B => mult_28_C96_n949, Z => 
                           mult_28_C96_n169);
   mult_28_C96_U162 : OAI21D1 port map( A1 => mult_28_C96_n167, A2 => 
                           mult_28_C96_n173, B => mult_28_C96_n168, Z => 
                           mult_28_C96_n162);
   mult_28_C96_U153 : NOR2D2 port map( A1 => mult_28_C96_n336, A2 => 
                           mult_28_C96_n343, Z => mult_28_C96_n154);
   mult_28_C96_U132 : OAI21D1 port map( A1 => mult_28_C96_n164, A2 => 
                           mult_28_C96_n143, B => mult_28_C96_n144, Z => 
                           mult_28_C96_n142);
   mult_28_C96_U120 : OAI21D1 port map( A1 => mult_28_C96_n134, A2 => 
                           mult_28_C96_n155, B => mult_28_C96_n135, Z => 
                           mult_28_C96_n133);
   mult_28_C96_U118 : AOI21D1 port map( A1 => mult_28_C96_n162, A2 => 
                           mult_28_C96_n969, B => mult_28_C96_n133, Z => 
                           mult_28_C96_n52);
   mult_28_C96_U111 : NOR2D2 port map( A1 => mult_28_C96_n316, A2 => 
                           mult_28_C96_n321, Z => mult_28_C96_n117);
   mult_28_C96_U80 : OAI21D1 port map( A1 => mult_28_C96_n113, A2 => 
                           mult_28_C96_n103, B => mult_28_C96_n104, Z => 
                           mult_28_C96_n102);
   mult_28_C96_U78 : AOI21D1 port map( A1 => mult_28_C96_n101, A2 => 
                           mult_28_C96_n960, B => mult_28_C96_n102, Z => 
                           mult_28_C96_n100);
   mult_28_C96_U69 : NOR2D2 port map( A1 => mult_28_C96_n307, A2 => 
                           mult_28_C96_n306, Z => mult_28_C96_n92);
   mult_28_C96_U54 : EXOR2D1 port map( A1 => mult_28_C96_n85, A2 => 
                           mult_28_C96_n54, Z => m5_15);

end flat_sec_par_16_5;
