
library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

package CONV_PACK_siso_gen is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type VHDLOUT_TYPE is array (0 downto 0) of std_logic;

end CONV_PACK_siso_gen;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_siso_gen.all;

architecture hier_sec_par_16_5 of siso_gen_DW_mult_tc_18 is

   component EXNOR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVDL
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22M10D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AO21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA22DL
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22DL
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21M10DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR3DL
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN3D2
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFDL
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component AOI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D4
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22D2
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR3D2
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFD4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFD2
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component EXOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADFULDL
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component NAN2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN3M1D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M10D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFD2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21M10D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INVBD32
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AO21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR3D4
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADFULD2
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component NOR2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AO21D2
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFD1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal n6, n9, n12, n16, n18, n22, n24, n28, n30, n34, n36, n40, n42, n46, 
      n48, n51, n52, n53, n54, n56, n57, n63, n65, n66, n67, n68, n69, n84, n85
      , n86, n87, n92, n93, n95, n96, n97, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n112, n113, n114, n115, n116, n117, n118, n127, 
      n128, n129, n133, n134, n135, n139, n140, n141, n142, n143, n144, n148, 
      n149, n150, n151, n152, n153, n154, n155, n160, n161, n162, n163, n164, 
      n167, n168, n169, n173, n175, n176, n177, n178, n179, n180, n182, n183, 
      n184, n187, n188, n189, n190, n192, n195, n196, n197, n199, n200, n201, 
      n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, 
      n214, n215, n217, n223, n225, n230, n232, n243, n248, n249, n250, n251, 
      n256, n257, n258, n259, n264, n265, n266, n267, n276, n278, n279, n281, 
      n282, n283, n284, n285, n286, n288, n305, n306, n307, n308, n309, n310, 
      n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, 
      n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, 
      n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, 
      n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, 
      n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, 
      n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, 
      n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, 
      n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, 
      n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, 
      n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, 
      n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, 
      n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, 
      n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, 
      n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, 
      n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, 
      n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, 
      n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, 
      n515, n516, n517, n518, n519, n520, n522, n523, n524, n525, n526, n527, 
      n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, 
      n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, 
      n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, 
      n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, 
      n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, 
      n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, 
      n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, 
      n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, 
      n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, 
      n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, 
      n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, 
      n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, 
      n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, 
      n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, 
      n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, 
      n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, 
      n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, 
      n732, n733, n734, n735, n736, n737, n738, n740, n741, n742, n743, n744, 
      n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, 
      n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, 
      n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, 
      n781, n782, n783, n784, n801, n802, n803, n804, n805, n806, n807, n808, 
      n824, n825, n826, n827, n828, n829, n830, n831, n832, n900, n901, n902, 
      n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, 
      n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, 
      n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, 
      n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, 
      n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, 
      n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, 
      n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, 
      n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, 
      n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, 
      n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, 
      n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, 
      n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, 
      n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, 
      n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, 
      n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, 
      n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, 
      n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, 
      n1089, n1090, n1091, n1092, n1093, n1094, n_1016 : std_logic;

begin
   
   U54 : EXOR2D1 port map( A1 => n85, A2 => n54, Z => product(29));
   U69 : NOR2D2 port map( A1 => n307, A2 => n306, Z => n92);
   U78 : AOI21D1 port map( A1 => n101, A2 => n960, B => n102, Z => n100);
   U80 : OAI21D1 port map( A1 => n113, A2 => n103, B => n104, Z => n102);
   U111 : NOR2D2 port map( A1 => n316, A2 => n321, Z => n117);
   U118 : AOI21D1 port map( A1 => n162, A2 => n969, B => n133, Z => n52);
   U120 : OAI21D1 port map( A1 => n134, A2 => n155, B => n135, Z => n133);
   U132 : OAI21D1 port map( A1 => n164, A2 => n143, B => n144, Z => n142);
   U153 : NOR2D2 port map( A1 => n336, A2 => n343, Z => n154);
   U162 : OAI21D1 port map( A1 => n167, A2 => n173, B => n168, Z => n162);
   U168 : AOI21D1 port map( A1 => n1020, A2 => n284, B => n949, Z => n169);
   U178 : AOI21D1 port map( A1 => n177, A2 => n190, B => n178, Z => n176);
   U183 : NOR2D2 port map( A1 => n364, A2 => n375, Z => n179);
   U193 : NOR2D2 port map( A1 => n376, A2 => n387, Z => n184);
   U202 : OAI21D1 port map( A1 => n201, A2 => n195, B => n196, Z => n190);
   U207 : EXNOR2D1 port map( A1 => n202, A2 => n67, Z => product(16));
   U217 : AOI21D1 port map( A1 => n204, A2 => n212, B => n205, Z => n203);
   U232 : OAI21D1 port map( A1 => n225, A2 => n213, B => n214, Z => n212);
   U278 : AOI21D1 port map( A1 => n248, A2 => n1071, B => n1083, Z => n243);
   U286 : OAI21D1 port map( A1 => n249, A2 => n251, B => n250, Z => n248);
   U292 : AOI21D1 port map( A1 => n256, A2 => n1084, B => n1085, Z => n251);
   U300 : OAI21D1 port map( A1 => n257, A2 => n259, B => n258, Z => n256);
   U306 : AOI21D1 port map( A1 => n1086, A2 => n264, B => n1087, Z => n259);
   U314 : OAI21D1 port map( A1 => n267, A2 => n265, B => n266, Z => n264);
   U320 : AOI21D1 port map( A1 => n1088, A2 => n1090, B => n1089, Z => n267);
   U334 : ADFULD1 port map( A => n522, B => n309, CI => n532, CO => n305, S => 
                           n306);
   U335 : ADFULD1 port map( A => n310, B => n523, CI => n313, CO => n307, S => 
                           n308);
   U337 : ADFULD1 port map( A => n317, B => n533, CI => n314, CO => n311, S => 
                           n312);
   U338 : ADFULD1 port map( A => n524, B => n319, CI => n548, CO => n313, S => 
                           n314);
   U339 : ADFULD1 port map( A => n318, B => n325, CI => n323, CO => n315, S => 
                           n316);
   U340 : ADFULD1 port map( A => n534, B => n320, CI => n549, CO => n317, S => 
                           n318);
   U342 : ADFULD1 port map( A => n329, B => n326, CI => n324, CO => n321, S => 
                           n322);
   U343 : ADFULD1 port map( A => n565, B => n535, CI => n331, CO => n323, S => 
                           n324);
   U345 : ADFULD1 port map( A => n337, B => n332, CI => n330, CO => n327, S => 
                           n328);
   U347 : ADFULD1 port map( A => n536, B => n334, CI => n551, CO => n331, S => 
                           n332);
   U349 : ADFULD1 port map( A => n345, B => n340, CI => n338, CO => n335, S => 
                           n336);
   U350 : ADFULD1 port map( A => n342, B => n349, CI => n347, CO => n337, S => 
                           n338);
   U351 : ADFULD1 port map( A => n567, B => n552, CI => n582, CO => n339, S => 
                           n340);
   U352 : ADFULD1 port map( A => n537, B => n351, CI => n526, CO => n341, S => 
                           n342);
   U353 : ADFULD1 port map( A => n355, B => n348, CI => n346, CO => n343, S => 
                           n344);
   U354 : ADFULD1 port map( A => n350, B => n359, CI => n357, CO => n345, S => 
                           n346);
   U355 : ADFULD1 port map( A => n583, B => n568, CI => n361, CO => n347, S => 
                           n348);
   U356 : ADFULD1 port map( A => n352, B => n538, CI => n553, CO => n349, S => 
                           n350);
   U359 : ADFULD1 port map( A => n360, B => n369, CI => n367, CO => n355, S => 
                           n356);
   U362 : ADFULD1 port map( A => n527, B => n373, CI => n554, CO => n361, S => 
                           n_1016);
   U363 : ADFULD1 port map( A => n377, B => n368, CI => n366, CO => n363, S => 
                           n364);
   U364 : ADFULD1 port map( A => n381, B => n370, CI => n379, CO => n365, S => 
                           n366);
   U365 : ADFULD1 port map( A => n383, B => n585, CI => n372, CO => n367, S => 
                           n368);
   U367 : ADFULD1 port map( A => n540, B => n374, CI => n555, CO => n371, S => 
                           n372);
   U372 : ADFULD1 port map( A => n601, B => n586, CI => n386, CO => n381, S => 
                           n382);
   U376 : ADFULD1 port map( A => n394, B => n407, CI => n405, CO => n389, S => 
                           n390);
   U379 : ADFULD1 port map( A => n572, B => n557, CI => n411, CO => n395, S => 
                           n396);
   U380 : ADFULD1 port map( A => n413, B => n400, CI => n542, CO => n397, S => 
                           n398);
   U382 : ADFULD1 port map( A => n417, B => n966, CI => n404, CO => n401, S => 
                           n402);
   U385 : ADFULD1 port map( A => n618, B => n603, CI => n412, CO => n407, S => 
                           n408);
   U387 : ADFULD1 port map( A => n414, B => n543, CI => n558, CO => n411, S => 
                           n412);
   U391 : ADFULD1 port map( A => n433, B => n424, CI => n422, CO => n417, S => 
                           n418);
   U398 : ADFULD1 port map( A => n445, B => n447, CI => n436, CO => n431, S => 
                           n432);
   U402 : ADFULD1 port map( A => n451, B => n531, CI => n545, CO => n439, S => 
                           n440);
   U404 : ADFULD1 port map( A => n457, B => n459, CI => n448, CO => n443, S => 
                           n444);
   U409 : ADFULD1 port map( A => n458, B => n465, CI => n456, CO => n453, S => 
                           n454);
   U410 : ADFULD1 port map( A => n460, B => n637, CI => n467, CO => n455, S => 
                           n456);
   U412 : ADFULD1 port map( A => n592, B => n577, CI => n462, CO => n459, S => 
                           n460);
   U413 : ADFULD1 port map( A => n471, B => n547, CI => n562, CO => n461, S => 
                           n462);
   U414 : ADFULD1 port map( A => n468, B => n475, CI => n466, CO => n463, S => 
                           n464);
   U415 : ADFULD1 port map( A => n470, B => n638, CI => n477, CO => n465, S => 
                           n466);
   U416 : ADFULD1 port map( A => n608, B => n479, CI => n623, CO => n467, S => 
                           n468);
   U417 : ADFULD1 port map( A => n578, B => n472, CI => n593, CO => n469, S => 
                           n470);
   U419 : ADFULD1 port map( A => n483, B => n478, CI => n476, CO => n473, S => 
                           n474);
   U420 : ADFULD1 port map( A => n639, B => n485, CI => n624, CO => n475, S => 
                           n476);
   U421 : ADFULD1 port map( A => n609, B => n594, CI => n480, CO => n477, S => 
                           n478);
   U422 : ADFULD1 port map( A => n487, B => n564, CI => n579, CO => n479, S => 
                           n480);
   U425 : ADFULD1 port map( A => n595, B => n488, CI => n610, CO => n485, S => 
                           n486);
   U426 : ADHALFD1 port map( A => n580, B => n516, CO => n487, S => n488);
   U427 : ADFULD1 port map( A => n641, B => n497, CI => n492, CO => n489, S => 
                           n490);
   U428 : ADFULD1 port map( A => n626, B => n611, CI => n494, CO => n491, S => 
                           n492);
   U429 : ADFULD1 port map( A => n499, B => n581, CI => n596, CO => n493, S => 
                           n494);
   U430 : ADFULD1 port map( A => n642, B => n503, CI => n498, CO => n495, S => 
                           n496);
   U431 : ADFULD1 port map( A => n612, B => n500, CI => n627, CO => n497, S => 
                           n498);
   U432 : ADHALFD1 port map( A => n597, B => n517, CO => n499, S => n500);
   U433 : ADFULD1 port map( A => n643, B => n628, CI => n504, CO => n501, S => 
                           n502);
   U434 : ADFULD1 port map( A => n507, B => n598, CI => n613, CO => n503, S => 
                           n504);
   U435 : ADFULD1 port map( A => n629, B => n508, CI => n644, CO => n505, S => 
                           n506);
   U436 : ADHALFD1 port map( A => n614, B => n518, CO => n507, S => n508);
   U437 : ADFULD1 port map( A => n511, B => n615, CI => n630, CO => n509, S => 
                           n510);
   U439 : OAI22D1 port map( A1 => n48, A2 => n825, B1 => n665, B2 => n46, Z => 
                           n513);
   U441 : OAI22D1 port map( A1 => n651, A2 => n48, B1 => n650, B2 => n46, Z => 
                           n522);
   U444 : OAI22D1 port map( A1 => n654, A2 => n48, B1 => n653, B2 => n46, Z => 
                           n319);
   U447 : OAI22D1 port map( A1 => n657, A2 => n48, B1 => n656, B2 => n46, Z => 
                           n526);
   U448 : OAI22D1 port map( A1 => n658, A2 => n48, B1 => n657, B2 => n46, Z => 
                           n351);
   U449 : OAI22D1 port map( A1 => n659, A2 => n48, B1 => n658, B2 => n46, Z => 
                           n527);
   U450 : OAI22D1 port map( A1 => n660, A2 => n48, B1 => n659, B2 => n46, Z => 
                           n373);
   U451 : OAI22D1 port map( A1 => n661, A2 => n48, B1 => n660, B2 => n46, Z => 
                           n528);
   U452 : OAI22D1 port map( A1 => n662, A2 => n48, B1 => n661, B2 => n46, Z => 
                           n399);
   U453 : OAI22D1 port map( A1 => n916, A2 => n48, B1 => n662, B2 => n46, Z => 
                           n529);
   U454 : OAI22D1 port map( A1 => n664, A2 => n48, B1 => n663, B2 => n46, Z => 
                           n530);
   U455 : NOR2M1D1 port map( A1 => b(0), A2 => n46, Z => n531);
   U471 : EXNOR2D1 port map( A1 => b(0), A2 => a(15), Z => n664);
   U472 : NAN2M1D1 port map( A1 => b(0), A2 => a(15), Z => n665);
   U473 : OAI22D1 port map( A1 => n42, A2 => n826, B1 => n682, B2 => n40, Z => 
                           n514);
   U475 : OAI22D1 port map( A1 => n667, A2 => n42, B1 => n666, B2 => n40, Z => 
                           n309);
   U476 : OAI22D1 port map( A1 => n668, A2 => n42, B1 => n667, B2 => n40, Z => 
                           n533);
   U477 : OAI22D1 port map( A1 => n669, A2 => n42, B1 => n668, B2 => n40, Z => 
                           n534);
   U478 : OAI22D1 port map( A1 => n670, A2 => n42, B1 => n669, B2 => n40, Z => 
                           n535);
   U479 : OAI22D1 port map( A1 => n671, A2 => n42, B1 => n670, B2 => n40, Z => 
                           n536);
   U480 : OAI22D1 port map( A1 => n671, A2 => n40, B1 => n672, B2 => n42, Z => 
                           n537);
   U481 : OAI22D1 port map( A1 => n673, A2 => n42, B1 => n672, B2 => n40, Z => 
                           n538);
   U483 : OAI22D1 port map( A1 => n675, A2 => n42, B1 => n674, B2 => n40, Z => 
                           n540);
   U485 : OAI22D1 port map( A1 => n677, A2 => n42, B1 => n676, B2 => n40, Z => 
                           n542);
   U486 : OAI22D1 port map( A1 => n678, A2 => n42, B1 => n677, B2 => n40, Z => 
                           n543);
   U487 : OAI22D1 port map( A1 => n679, A2 => n42, B1 => n678, B2 => n40, Z => 
                           n544);
   U488 : OAI22D1 port map( A1 => n994, A2 => n42, B1 => n679, B2 => n40, Z => 
                           n545);
   U489 : OAI22D1 port map( A1 => n681, A2 => n42, B1 => n680, B2 => n40, Z => 
                           n546);
   U490 : NOR2M1D1 port map( A1 => b(0), A2 => n40, Z => n547);
   U506 : EXNOR2D1 port map( A1 => b(0), A2 => a(13), Z => n681);
   U507 : NAN2M1D1 port map( A1 => b(0), A2 => a(13), Z => n682);
   U508 : OAI22D1 port map( A1 => n36, A2 => n827, B1 => n699, B2 => n34, Z => 
                           n515);
   U511 : OAI22D1 port map( A1 => n685, A2 => n36, B1 => n684, B2 => n34, Z => 
                           n550);
   U513 : OAI22D1 port map( A1 => n687, A2 => n36, B1 => n686, B2 => n34, Z => 
                           n552);
   U515 : OAI22D1 port map( A1 => n688, A2 => n34, B1 => n689, B2 => n36, Z => 
                           n554);
   U516 : OAI22D1 port map( A1 => n690, A2 => n36, B1 => n689, B2 => n34, Z => 
                           n555);
   U518 : OAI22D1 port map( A1 => n692, A2 => n36, B1 => n691, B2 => n34, Z => 
                           n557);
   U519 : OAI22D1 port map( A1 => n693, A2 => n36, B1 => n692, B2 => n34, Z => 
                           n558);
   U520 : OAI22D1 port map( A1 => n694, A2 => n36, B1 => n693, B2 => n34, Z => 
                           n559);
   U521 : OAI22D1 port map( A1 => n695, A2 => n36, B1 => n694, B2 => n34, Z => 
                           n560);
   U522 : OAI22D1 port map( A1 => n696, A2 => n36, B1 => n695, B2 => n34, Z => 
                           n561);
   U523 : OAI22D1 port map( A1 => n697, A2 => n36, B1 => n696, B2 => n34, Z => 
                           n562);
   U524 : OAI22D1 port map( A1 => n698, A2 => n36, B1 => n697, B2 => n34, Z => 
                           n563);
   U525 : NOR2M1D1 port map( A1 => b(0), A2 => n34, Z => n564);
   U541 : EXNOR2D1 port map( A1 => b(0), A2 => a(11), Z => n698);
   U542 : NAN2M1D1 port map( A1 => b(0), A2 => a(11), Z => n699);
   U543 : OAI22D1 port map( A1 => n30, A2 => n828, B1 => n716, B2 => n28, Z => 
                           n516);
   U544 : AO21D2 port map( A1 => n30, A2 => n28, B => n700, Z => n565);
   U546 : OAI22D1 port map( A1 => n702, A2 => n30, B1 => n701, B2 => n28, Z => 
                           n567);
   U547 : OAI22D1 port map( A1 => n703, A2 => n30, B1 => n702, B2 => n28, Z => 
                           n568);
   U548 : OAI22D1 port map( A1 => n704, A2 => n30, B1 => n703, B2 => n28, Z => 
                           n569);
   U551 : OAI22D1 port map( A1 => n707, A2 => n30, B1 => n706, B2 => n28, Z => 
                           n572);
   U553 : OAI22D1 port map( A1 => n709, A2 => n30, B1 => n708, B2 => n28, Z => 
                           n574);
   U554 : OAI22D1 port map( A1 => n710, A2 => n30, B1 => n709, B2 => n28, Z => 
                           n575);
   U555 : OAI22D1 port map( A1 => n711, A2 => n30, B1 => n710, B2 => n28, Z => 
                           n576);
   U556 : OAI22D1 port map( A1 => n712, A2 => n30, B1 => n711, B2 => n28, Z => 
                           n577);
   U557 : OAI22D1 port map( A1 => n713, A2 => n30, B1 => n712, B2 => n28, Z => 
                           n578);
   U558 : OAI22D1 port map( A1 => n714, A2 => n30, B1 => n713, B2 => n28, Z => 
                           n579);
   U559 : OAI22D1 port map( A1 => n715, A2 => n30, B1 => n714, B2 => n28, Z => 
                           n580);
   U560 : NOR2M1D1 port map( A1 => b(0), A2 => n28, Z => n581);
   U576 : EXNOR2D1 port map( A1 => b(0), A2 => a(9), Z => n715);
   U577 : NAN2M1D1 port map( A1 => b(0), A2 => a(9), Z => n716);
   U578 : OAI22D1 port map( A1 => n24, A2 => n829, B1 => n733, B2 => n22, Z => 
                           n517);
   U579 : AO21D2 port map( A1 => n24, A2 => n22, B => n717, Z => n582);
   U581 : OAI22D1 port map( A1 => n719, A2 => n24, B1 => n718, B2 => n22, Z => 
                           n584);
   U582 : OAI22D1 port map( A1 => n720, A2 => n24, B1 => n719, B2 => n22, Z => 
                           n585);
   U584 : OAI22D1 port map( A1 => n722, A2 => n24, B1 => n1002, B2 => n22, Z =>
                           n587);
   U585 : OAI22D1 port map( A1 => n722, A2 => n22, B1 => n723, B2 => n24, Z => 
                           n588);
   U586 : OAI22D1 port map( A1 => n724, A2 => n24, B1 => n723, B2 => n22, Z => 
                           n589);
   U587 : OAI22D1 port map( A1 => n24, A2 => n725, B1 => n724, B2 => n22, Z => 
                           n590);
   U588 : OAI22D1 port map( A1 => n726, A2 => n24, B1 => n725, B2 => n22, Z => 
                           n591);
   U589 : OAI22D1 port map( A1 => n727, A2 => n24, B1 => n726, B2 => n22, Z => 
                           n592);
   U590 : OAI22D1 port map( A1 => n728, A2 => n24, B1 => n727, B2 => n22, Z => 
                           n593);
   U591 : OAI22D1 port map( A1 => n729, A2 => n24, B1 => n728, B2 => n22, Z => 
                           n594);
   U592 : OAI22D1 port map( A1 => n730, A2 => n24, B1 => n729, B2 => n22, Z => 
                           n595);
   U593 : OAI22D1 port map( A1 => n731, A2 => n24, B1 => n730, B2 => n22, Z => 
                           n596);
   U594 : OAI22D1 port map( A1 => n732, A2 => n24, B1 => n731, B2 => n22, Z => 
                           n597);
   U595 : NOR2M1D1 port map( A1 => b(0), A2 => n22, Z => n598);
   U596 : EXNOR2D1 port map( A1 => b(15), A2 => a(7), Z => n717);
   U611 : EXNOR2D1 port map( A1 => b(0), A2 => a(7), Z => n732);
   U612 : NAN2M1D1 port map( A1 => b(0), A2 => a(7), Z => n733);
   U613 : OAI22D1 port map( A1 => n18, A2 => n830, B1 => n750, B2 => n16, Z => 
                           n518);
   U616 : OAI22D1 port map( A1 => n736, A2 => n18, B1 => n735, B2 => n16, Z => 
                           n601);
   U621 : OAI22D1 port map( A1 => n741, A2 => n18, B1 => n740, B2 => n16, Z => 
                           n606);
   U623 : OAI22D1 port map( A1 => n743, A2 => n18, B1 => n742, B2 => n16, Z => 
                           n608);
   U624 : OAI22D1 port map( A1 => n744, A2 => n18, B1 => n743, B2 => n16, Z => 
                           n609);
   U625 : OAI22D1 port map( A1 => n745, A2 => n18, B1 => n744, B2 => n16, Z => 
                           n610);
   U626 : OAI22D1 port map( A1 => n746, A2 => n18, B1 => n745, B2 => n16, Z => 
                           n611);
   U627 : OAI22D1 port map( A1 => n747, A2 => n18, B1 => n746, B2 => n16, Z => 
                           n612);
   U628 : OAI22D1 port map( A1 => n748, A2 => n18, B1 => n747, B2 => n16, Z => 
                           n613);
   U629 : OAI22D1 port map( A1 => n749, A2 => n18, B1 => n748, B2 => n16, Z => 
                           n614);
   U630 : NOR2M1D1 port map( A1 => b(0), A2 => n16, Z => n615);
   U642 : EXNOR2D1 port map( A1 => b(4), A2 => a(5), Z => n745);
   U646 : EXNOR2D1 port map( A1 => b(0), A2 => a(5), Z => n749);
   U647 : NAN2M1D1 port map( A1 => b(0), A2 => a(5), Z => n750);
   U648 : OAI22D1 port map( A1 => n12, A2 => n831, B1 => n767, B2 => n9, Z => 
                           n519);
   U652 : OAI22D1 port map( A1 => n754, A2 => n12, B1 => n753, B2 => n9, Z => 
                           n619);
   U653 : OAI22D1 port map( A1 => n12, A2 => n755, B1 => n754, B2 => n9, Z => 
                           n620);
   U654 : OAI22D1 port map( A1 => n756, A2 => n12, B1 => n755, B2 => n9, Z => 
                           n621);
   U655 : OAI22D1 port map( A1 => n756, A2 => n9, B1 => n757, B2 => n12, Z => 
                           n622);
   U657 : OAI22D1 port map( A1 => n759, A2 => n12, B1 => n758, B2 => n9, Z => 
                           n624);
   U658 : OAI22D1 port map( A1 => n760, A2 => n12, B1 => n759, B2 => n9, Z => 
                           n625);
   U659 : OAI22D1 port map( A1 => n761, A2 => n12, B1 => n760, B2 => n9, Z => 
                           n626);
   U660 : OAI22D1 port map( A1 => n762, A2 => n12, B1 => n761, B2 => n9, Z => 
                           n627);
   U661 : OAI22D1 port map( A1 => n763, A2 => n12, B1 => n762, B2 => n9, Z => 
                           n628);
   U662 : OAI22D1 port map( A1 => n764, A2 => n12, B1 => n763, B2 => n9, Z => 
                           n629);
   U663 : OAI22D1 port map( A1 => n765, A2 => n12, B1 => n764, B2 => n9, Z => 
                           n630);
   U664 : OAI22D1 port map( A1 => n766, A2 => n12, B1 => n765, B2 => n9, Z => 
                           n631);
   U665 : NOR2M1D1 port map( A1 => b(0), A2 => n9, Z => n632);
   U666 : EXNOR2D1 port map( A1 => b(15), A2 => a(3), Z => n751);
   U677 : EXNOR2D1 port map( A1 => b(4), A2 => a(3), Z => n762);
   U681 : EXNOR2D1 port map( A1 => b(0), A2 => a(3), Z => n766);
   U682 : NAN2M1D1 port map( A1 => b(0), A2 => a(3), Z => n767);
   U683 : OAI22D1 port map( A1 => n6, A2 => n832, B1 => n784, B2 => n824, Z => 
                           n520);
   U688 : OAI22D1 port map( A1 => n772, A2 => n6, B1 => n771, B2 => n824, Z => 
                           n637);
   U690 : OAI22D1 port map( A1 => n773, A2 => n824, B1 => n774, B2 => n6, Z => 
                           n639);
   U692 : OAI22D1 port map( A1 => n776, A2 => n6, B1 => n775, B2 => n824, Z => 
                           n641);
   U693 : OAI22D1 port map( A1 => n777, A2 => n6, B1 => n776, B2 => n824, Z => 
                           n642);
   U694 : OAI22D1 port map( A1 => n778, A2 => n6, B1 => n777, B2 => n824, Z => 
                           n643);
   U695 : OAI22D1 port map( A1 => n779, A2 => n6, B1 => n778, B2 => n824, Z => 
                           n644);
   U696 : OAI22D1 port map( A1 => n780, A2 => n6, B1 => n779, B2 => n824, Z => 
                           n645);
   U698 : OAI22D1 port map( A1 => n782, A2 => n6, B1 => n781, B2 => n824, Z => 
                           n647);
   U699 : OAI22D1 port map( A1 => n783, A2 => n6, B1 => n782, B2 => n824, Z => 
                           n648);
   U712 : EXNOR2D1 port map( A1 => b(4), A2 => a(1), Z => n779);
   U716 : EXNOR2D1 port map( A1 => b(0), A2 => a(1), Z => n783);
   U717 : NAN2M1D1 port map( A1 => b(0), A2 => a(1), Z => n784);
   U742 : EXOR2D1 port map( A1 => a(15), A2 => a(14), Z => n801);
   U745 : EXOR2D1 port map( A1 => a(13), A2 => a(12), Z => n802);
   U748 : EXOR2D1 port map( A1 => a(11), A2 => a(10), Z => n803);
   U751 : EXOR2D1 port map( A1 => a(9), A2 => a(8), Z => n804);
   U754 : EXOR2D1 port map( A1 => a(7), A2 => a(6), Z => n805);
   U757 : EXOR2D1 port map( A1 => a(5), A2 => a(4), Z => n806);
   U760 : EXOR2D1 port map( A1 => a(3), A2 => a(2), Z => n807);
   U763 : EXOR2D1 port map( A1 => a(1), A2 => a(0), Z => n808);
   U767 : OAI22D2 port map( A1 => n735, A2 => n18, B1 => n734, B2 => n16, Z => 
                           n600);
   U768 : NAN2D1 port map( A1 => n454, A2 => n463, Z => n223);
   U769 : OAI22D1 port map( A1 => n900, A2 => n721, B1 => n720, B2 => n22, Z =>
                           n586);
   U770 : INVBD32 port map( A => n903, Z => n900);
   U771 : EXOR2D1 port map( A1 => n1037, A2 => n423, Z => n406);
   U772 : OAI22D1 port map( A1 => n18, A2 => n1060, B1 => n738, B2 => n16, Z =>
                           n901);
   U773 : OAI22DL port map( A1 => n18, A2 => n1060, B1 => n738, B2 => n16, Z =>
                           n604);
   U774 : EXNOR2D2 port map( A1 => b(11), A2 => a(5), Z => n738);
   U775 : OAI22D1 port map( A1 => n754, A2 => n12, B1 => n753, B2 => n9, Z => 
                           n902);
   U776 : EXNOR2DL port map( A1 => b(8), A2 => a(9), Z => n908);
   U777 : EXOR2D2 port map( A1 => n1037, A2 => n423, Z => n966);
   U778 : INVBD32 port map( A => n24, Z => n903);
   U779 : INVDL port map( A => n605, Z => n904);
   U780 : INVD1 port map( A => n904, Z => n905);
   U781 : EXNOR2DL port map( A1 => b(6), A2 => a(15), Z => n658);
   U782 : ADFULD2 port map( A => n397, B => n571, CI => n556, CO => n383, S => 
                           n384);
   U783 : OAI22DL port map( A1 => n781, A2 => n6, B1 => n780, B2 => n824, Z => 
                           n646);
   U784 : OAI22D1 port map( A1 => n737, A2 => n18, B1 => n736, B2 => n16, Z => 
                           n906);
   U785 : OAI22DL port map( A1 => n737, A2 => n18, B1 => n736, B2 => n16, Z => 
                           n602);
   U786 : OAI22M10D1 port map( A1 => n907, A2 => n740, B1 => n1060, B2 => n16, 
                           Z => n605);
   U787 : INVBD32 port map( A => n18, Z => n907);
   U788 : EXNOR2D1 port map( A1 => b(8), A2 => a(9), Z => n707);
   U789 : EXNOR2D1 port map( A1 => b(11), A2 => a(9), Z => n704);
   U790 : EXNOR2DL port map( A1 => b(6), A2 => a(13), Z => n675);
   U791 : EXOR3D1 port map( A1 => n392, A2 => n403, A3 => n390, Z => n909);
   U792 : EXOR3D1 port map( A1 => n392, A2 => n403, A3 => n390, Z => n388);
   U793 : EXNOR3D4 port map( A1 => n617, A2 => n409, A3 => n967, Z => n392);
   U794 : BUFDL port map( A => n179, Z => n910);
   U795 : EXNOR2DL port map( A1 => b(14), A2 => a(3), Z => n752);
   U796 : OAI22D1 port map( A1 => n677, A2 => n42, B1 => n676, B2 => n40, Z => 
                           n911);
   U797 : NOR2DL port map( A1 => n913, A2 => n200, Z => n912);
   U798 : AO21M20D1 port map( A1 => n52, A2 => n117, B => n960, Z => n116);
   U799 : EXNOR2D2 port map( A1 => b(10), A2 => a(11), Z => n688);
   U800 : EXNOR2D2 port map( A1 => b(7), A2 => a(11), Z => n691);
   U801 : INVD1 port map( A => b(7), Z => n1041);
   U802 : AOI21DL port map( A1 => n141, A2 => n1020, B => n142, Z => n140);
   U803 : NOR2D2 port map( A1 => n388, A2 => n401, Z => n913);
   U804 : NOR2D1 port map( A1 => n909, A2 => n401, Z => n195);
   U805 : INVDL port map( A => n286, Z => n914);
   U806 : INVDL port map( A => n663, Z => n915);
   U807 : INVD1 port map( A => n915, Z => n916);
   U808 : EXNOR2D2 port map( A1 => n140, A2 => n917, Z => product(24));
   U809 : AND2DL port map( A1 => n1078, A2 => n139, Z => n917);
   U810 : NOR2D2 port map( A1 => n134, A2 => n154, Z => n969);
   U811 : NOR2D1 port map( A1 => n354, A2 => n363, Z => n1028);
   U812 : INVDL port map( A => n908, Z => n918);
   U813 : INVD1 port map( A => n918, Z => n919);
   U814 : EXOR2D1 port map( A1 => n1029, A2 => n584, Z => n360);
   U815 : EXNOR2D2 port map( A1 => b(4), A2 => a(9), Z => n711);
   U816 : EXNOR2D2 port map( A1 => b(4), A2 => a(13), Z => n677);
   U817 : EXNOR2D2 port map( A1 => b(4), A2 => a(11), Z => n694);
   U818 : EXNOR2DL port map( A1 => b(4), A2 => a(7), Z => n728);
   U819 : NAN2D1 port map( A1 => n574, A2 => n439, Z => n1034);
   U820 : EXOR3D2 port map( A1 => n625, A2 => n493, A3 => n640, Z => n484);
   U821 : EXOR2D1 port map( A1 => n491, A2 => n486, Z => n920);
   U822 : EXOR2D1 port map( A1 => n920, A2 => n484, Z => n482);
   U823 : NAN2DL port map( A1 => n625, A2 => n493, Z => n921);
   U824 : NAN2DL port map( A1 => n625, A2 => n640, Z => n922);
   U825 : NAN2DL port map( A1 => n493, A2 => n640, Z => n923);
   U826 : NAN3D1 port map( A1 => n921, A2 => n922, A3 => n923, Z => n483);
   U827 : NAN2D1 port map( A1 => n491, A2 => n486, Z => n924);
   U828 : NAN2DL port map( A1 => n491, A2 => n484, Z => n925);
   U829 : NAN2DL port map( A1 => n486, A2 => n484, Z => n926);
   U830 : NAN3D1 port map( A1 => n924, A2 => n925, A3 => n926, Z => n481);
   U831 : BUFDL port map( A => n435, Z => n927);
   U832 : OAI22D1 port map( A1 => n928, A2 => n752, B1 => n753, B2 => n12, Z =>
                           n618);
   U833 : INVBD32 port map( A => n933, Z => n928);
   U834 : EXNOR2D2 port map( A1 => n529, A2 => n427, Z => n414);
   U835 : NOR2D1 port map( A1 => n328, A2 => n335, Z => n149);
   U836 : OAI22D1 port map( A1 => n686, A2 => n36, B1 => n685, B2 => n34, Z => 
                           n551);
   U837 : INVD1 port map( A => n118, Z => n960);
   U838 : NOR2D1 port map( A1 => n311, A2 => n308, Z => n103);
   U839 : NAN2D1 port map( A1 => n161, A2 => n969, Z => n53);
   U840 : NOR2D1 port map( A1 => n312, A2 => n315, Z => n112);
   U841 : INVD1 port map( A => n9, Z => n933);
   U842 : EXOR3D1 port map( A1 => n575, A2 => n560, A3 => n440, Z => n438);
   U843 : OAI22D1 port map( A1 => n676, A2 => n42, B1 => n675, B2 => n40, Z => 
                           n541);
   U844 : NAN2D1 port map( A1 => n376, A2 => n387, Z => n187);
   U845 : INVDL port map( A => n53, Z => n128);
   U846 : INVD1 port map( A => n56, Z => n1017);
   U847 : INVDL port map( A => n92, Z => n276);
   U848 : AND2DL port map( A1 => n389, A2 => n380, Z => n929);
   U849 : ADHALFD2 port map( A => n563, B => n515, CO => n471, S => n472);
   U850 : EXOR3D1 port map( A1 => n461, A2 => n591, A3 => n606, Z => n448);
   U851 : NAN2DL port map( A1 => n606, A2 => n461, Z => n976);
   U852 : NAN2M1DL port map( A1 => n209, A2 => n210, Z => n69);
   U853 : NOR2DL port map( A1 => n206, A2 => n209, Z => n204);
   U854 : AOI21M10D1 port map( A1 => n930, A2 => n230, B => n1079, Z => n225);
   U855 : NOR2DL port map( A1 => n464, A2 => n473, Z => n930);
   U856 : ADFULD1 port map( A => n621, B => n450, CI => n636, CO => n445, S => 
                           n446);
   U857 : INVDL port map( A => b(12), Z => n931);
   U858 : INVD1 port map( A => n931, Z => n932);
   U859 : EXNOR2D2 port map( A1 => b(4), A2 => a(15), Z => n660);
   U860 : EXNOR2D1 port map( A1 => n208, A2 => n68, Z => product(15));
   U861 : AOI21D1 port map( A1 => n162, A2 => n969, B => n133, Z => n934);
   U862 : INVD1 port map( A => n399, Z => n400);
   U863 : BUFD2 port map( A => n399, Z => n993);
   U864 : OAI22D1 port map( A1 => n735, A2 => n18, B1 => n734, B2 => n16, Z => 
                           n935);
   U865 : EXNOR2D2 port map( A1 => b(8), A2 => a(7), Z => n724);
   U866 : EXNOR2DL port map( A1 => b(8), A2 => a(5), Z => n741);
   U867 : EXOR3D1 port map( A1 => n634, A2 => n604, A3 => n1050, Z => n422);
   U868 : NAN2D1 port map( A1 => n953, A2 => n587, Z => n984);
   U869 : EXOR3D2 port map( A1 => n410, A2 => n419, A3 => n408, Z => n404);
   U870 : EXNOR2DL port map( A1 => b(9), A2 => a(3), Z => n757);
   U871 : EXOR2D1 port map( A1 => n446, A2 => n455, Z => n936);
   U872 : EXOR2D1 port map( A1 => n936, A2 => n444, Z => n442);
   U873 : NAN2DL port map( A1 => n444, A2 => n455, Z => n937);
   U874 : NAN2DL port map( A1 => n444, A2 => n446, Z => n938);
   U875 : NAN2DL port map( A1 => n455, A2 => n446, Z => n939);
   U876 : NAN3D1 port map( A1 => n937, A2 => n939, A3 => n938, Z => n441);
   U877 : INVDL port map( A => n217, Z => n215);
   U878 : EXOR2D1 port map( A1 => n635, A2 => n620, Z => n940);
   U879 : EXOR2D1 port map( A1 => n940, A2 => n438, Z => n434);
   U880 : NAN2DL port map( A1 => n575, A2 => n560, Z => n941);
   U881 : NAN2DL port map( A1 => n575, A2 => n440, Z => n942);
   U882 : NAN2DL port map( A1 => n560, A2 => n440, Z => n943);
   U883 : NAN3D1 port map( A1 => n941, A2 => n942, A3 => n943, Z => n437);
   U884 : NAN2DL port map( A1 => n620, A2 => n635, Z => n944);
   U885 : NAN2DL port map( A1 => n620, A2 => n438, Z => n945);
   U886 : NAN2DL port map( A1 => n635, A2 => n438, Z => n946);
   U887 : NAN3D2 port map( A1 => n944, A2 => n945, A3 => n946, Z => n433);
   U888 : EXOR2D1 port map( A1 => n998, A2 => n927, Z => n420);
   U889 : NAN2DL port map( A1 => n434, A2 => n443, Z => n1006);
   U890 : NAN2DL port map( A1 => n421, A2 => n423, Z => n1040);
   U891 : NAN2DL port map( A1 => n633, A2 => n421, Z => n1038);
   U892 : EXNOR2DL port map( A1 => b(15), A2 => a(9), Z => n700);
   U893 : EXNOR2DL port map( A1 => b(11), A2 => a(5), Z => n947);
   U894 : NOR2D1 port map( A1 => n430, A2 => n441, Z => n209);
   U895 : EXNOR2D2 port map( A1 => n1008, A2 => a(13), Z => n672);
   U896 : EXNOR2DL port map( A1 => b(15), A2 => a(13), Z => n666);
   U897 : EXNOR2DL port map( A1 => b(15), A2 => a(11), Z => n683);
   U898 : NAN3D2 port map( A1 => n1024, A2 => n1026, A3 => n1025, Z => n403);
   U899 : NAN2D1 port map( A1 => n419, A2 => n408, Z => n1024);
   U900 : EXNOR2D2 port map( A1 => b(13), A2 => a(3), Z => n753);
   U901 : EXNOR2D2 port map( A1 => b(13), A2 => a(1), Z => n770);
   U902 : EXNOR2D1 port map( A1 => b(1), A2 => a(15), Z => n663);
   U903 : BUFD1 port map( A => n426, Z => n1050);
   U904 : INVDL port map( A => n203, Z => n202);
   U905 : OAI21M10D1 port map( A1 => n948, A2 => n463, B => n215, Z => n213);
   U906 : INVDL port map( A => n454, Z => n948);
   U907 : AOI21D1 port map( A1 => n283, A2 => n949, B => n950, Z => n164);
   U908 : INVDL port map( A => n173, Z => n949);
   U909 : INVDL port map( A => n168, Z => n950);
   U910 : NAN2M1D1 port map( A1 => n951, A2 => n393, Z => n1055);
   U911 : INVDL port map( A => n616, Z => n951);
   U912 : EXOR3D1 port map( A1 => n527, A2 => n373, A3 => n554, Z => n362);
   U913 : NAN3M1D1 port map( A1 => n929, A2 => n1094, A3 => n1093, Z => n375);
   U914 : OAI22D1 port map( A1 => n30, A2 => n706, B1 => n28, B2 => n705, Z => 
                           n571);
   U915 : OAI22D1 port map( A1 => n717, A2 => n22, B1 => n718, B2 => n24, Z => 
                           n583);
   U916 : EXOR2D4 port map( A1 => n962, A2 => n362, Z => n358);
   U917 : NAN2DL port map( A1 => n356, A2 => n358, Z => n972);
   U918 : EXNOR2DL port map( A1 => b(10), A2 => a(9), Z => n705);
   U919 : BUFDL port map( A => n161, Z => n952);
   U920 : EXNOR2D2 port map( A1 => b(5), A2 => a(5), Z => n744);
   U921 : EXOR3D1 port map( A1 => n400, A2 => n413, A3 => n911, Z => n953);
   U922 : OAI21DL port map( A1 => n201, A2 => n913, B => n196, Z => n954);
   U923 : EXNOR2D2 port map( A1 => b(9), A2 => a(5), Z => n740);
   U924 : EXNOR2D2 port map( A1 => b(9), A2 => a(9), Z => n706);
   U925 : INVD1 port map( A => n161, Z => n163);
   U926 : NAN2M1D1 port map( A1 => n955, A2 => n1077, Z => n1068);
   U927 : NOR2DL port map( A1 => n482, A2 => n489, Z => n955);
   U928 : EXOR2D1 port map( A1 => n566, A2 => n341, Z => n956);
   U929 : EXOR2D1 port map( A1 => n956, A2 => n339, Z => n330);
   U930 : NAN2DL port map( A1 => n339, A2 => n341, Z => n957);
   U931 : NAN2DL port map( A1 => n339, A2 => n566, Z => n958);
   U932 : NAN2D1 port map( A1 => n341, A2 => n566, Z => n959);
   U933 : NAN3D1 port map( A1 => n957, A2 => n959, A3 => n958, Z => n329);
   U934 : OAI22DL port map( A1 => n701, A2 => n30, B1 => n700, B2 => n28, Z => 
                           n566);
   U935 : INVDL port map( A => n167, Z => n283);
   U936 : EXNOR2D2 port map( A1 => b(15), A2 => a(5), Z => n734);
   U937 : OAI22D1 port map( A1 => n775, A2 => n6, B1 => n774, B2 => n824, Z => 
                           n640);
   U938 : OAI22DL port map( A1 => n654, A2 => n46, B1 => n655, B2 => n48, Z => 
                           n525);
   U939 : EXNOR2D2 port map( A1 => b(6), A2 => a(7), Z => n726);
   U940 : EXNOR2D2 port map( A1 => b(6), A2 => a(9), Z => n709);
   U941 : OA21M20D1 port map( A1 => n1077, A2 => n1072, B => n961, Z => n232);
   U942 : NAN2DL port map( A1 => n481, A2 => n474, Z => n961);
   U943 : NAN3D1 port map( A1 => n1046, A2 => n1048, A3 => n1047, Z => n409);
   U944 : OAI22D1 port map( A1 => n708, A2 => n30, B1 => n919, B2 => n28, Z => 
                           n573);
   U945 : EXOR2D1 port map( A1 => n599, A2 => n371, Z => n962);
   U946 : NAN2D1 port map( A1 => n362, A2 => n371, Z => n963);
   U947 : NAN2D1 port map( A1 => n362, A2 => n599, Z => n964);
   U948 : NAN2DL port map( A1 => n371, A2 => n599, Z => n965);
   U949 : NAN3D2 port map( A1 => n963, A2 => n965, A3 => n964, Z => n357);
   U950 : EXOR2D2 port map( A1 => n633, A2 => n421, Z => n1037);
   U951 : INVDL port map( A => n396, Z => n967);
   U952 : EXNOR2D2 port map( A1 => b(12), A2 => a(1), Z => n771);
   U953 : BUFDL port map( A => n912, Z => n968);
   U954 : EXNOR2D2 port map( A1 => b(1), A2 => a(11), Z => n697);
   U955 : EXNOR2DL port map( A1 => b(9), A2 => a(11), Z => n689);
   U956 : EXOR2D1 port map( A1 => n358, A2 => n365, Z => n970);
   U957 : EXOR2D1 port map( A1 => n970, A2 => n356, Z => n354);
   U958 : NAN2DL port map( A1 => n356, A2 => n365, Z => n971);
   U959 : NAN2DL port map( A1 => n365, A2 => n358, Z => n973);
   U960 : NAN3D1 port map( A1 => n971, A2 => n973, A3 => n972, Z => n353);
   U961 : OAI21D1 port map( A1 => n187, A2 => n179, B => n180, Z => n178);
   U962 : NAN2DL port map( A1 => n591, A2 => n606, Z => n974);
   U963 : NAN2DL port map( A1 => n591, A2 => n461, Z => n975);
   U964 : NAN3D1 port map( A1 => n974, A2 => n976, A3 => n975, Z => n447);
   U965 : EXNOR2DL port map( A1 => b(8), A2 => a(15), Z => n656);
   U966 : ADFULDL port map( A => n333, B => n525, CI => n550, CO => n325, S => 
                           n326);
   U967 : EXOR2D1 port map( A1 => n1013, A2 => n977, Z => n458);
   U968 : EXOR2DL port map( A1 => n469, A2 => n607, Z => n1013);
   U969 : BUFDL port map( A => n622, Z => n977);
   U970 : INVDL port map( A => n391, Z => n978);
   U971 : INVD1 port map( A => n978, Z => n979);
   U972 : ADHALFD2 port map( A => n513, B => n530, CO => n427, S => n428);
   U973 : NAN3D1 port map( A1 => n1038, A2 => n1039, A3 => n1040, Z => n405);
   U974 : NOR2D1 port map( A1 => n163, A2 => n154, Z => n152);
   U975 : OAI21DL port map( A1 => n164, A2 => n154, B => n155, Z => n153);
   U976 : EXOR3D2 port map( A1 => n935, A2 => n385, A3 => n570, Z => n370);
   U977 : NAN2DL port map( A1 => n385, A2 => n570, Z => n980);
   U978 : NAN2DL port map( A1 => n385, A2 => n600, Z => n981);
   U979 : NAN2DL port map( A1 => n570, A2 => n600, Z => n982);
   U980 : NAN3D1 port map( A1 => n980, A2 => n982, A3 => n981, Z => n369);
   U981 : OAI22DL port map( A1 => n705, A2 => n30, B1 => n704, B2 => n28, Z => 
                           n570);
   U982 : NAN3D2 port map( A1 => n999, A2 => n1000, A3 => n1001, Z => n419);
   U983 : NAN2D1 port map( A1 => n449, A2 => n590, Z => n995);
   U984 : ADFULD1 port map( A => n561, B => n452, CI => n576, CO => n449, S => 
                           n450);
   U985 : EXOR2D1 port map( A1 => n1009, A2 => n418, Z => n416);
   U986 : EXNOR2D2 port map( A1 => b(11), A2 => a(3), Z => n755);
   U987 : EXNOR2D1 port map( A1 => b(11), A2 => a(7), Z => n1002);
   U988 : OAI22DL port map( A1 => n691, A2 => n36, B1 => n690, B2 => n34, Z => 
                           n556);
   U989 : OAI22D1 port map( A1 => n656, A2 => n48, B1 => n655, B2 => n46, Z => 
                           n333);
   U990 : EXNOR2D2 port map( A1 => b(12), A2 => a(3), Z => n754);
   U991 : EXOR3D2 port map( A1 => n398, A2 => n587, A3 => n906, Z => n394);
   U992 : NAN2D1 port map( A1 => n602, A2 => n953, Z => n983);
   U993 : NAN2D1 port map( A1 => n906, A2 => n587, Z => n985);
   U994 : NAN3D2 port map( A1 => n985, A2 => n983, A3 => n984, Z => n393);
   U995 : EXNOR2DL port map( A1 => b(3), A2 => a(3), Z => n763);
   U996 : NAN2DL port map( A1 => n588, A2 => n573, Z => n1046);
   U997 : NAN2DL port map( A1 => n588, A2 => n425, Z => n1047);
   U998 : EXOR3D2 port map( A1 => n425, A2 => n588, A3 => n573, Z => n410);
   U999 : INVD1 port map( A => n150, Z => n148);
   U1000 : EXOR2D1 port map( A1 => n993, A2 => n528, Z => n986);
   U1001 : EXOR2D1 port map( A1 => n986, A2 => n541, Z => n386);
   U1002 : NAN2D1 port map( A1 => n541, A2 => n528, Z => n987);
   U1003 : NAN2D1 port map( A1 => n993, A2 => n541, Z => n988);
   U1004 : NAN2D1 port map( A1 => n528, A2 => n993, Z => n989);
   U1005 : NAN3D2 port map( A1 => n987, A2 => n989, A3 => n988, Z => n385);
   U1006 : EXNOR2DL port map( A1 => b(8), A2 => a(11), Z => n690);
   U1007 : NOR2D1 port map( A1 => n442, A2 => n453, Z => n217);
   U1008 : EXOR3D1 port map( A1 => n382, A2 => n384, A3 => n979, Z => n378);
   U1009 : NAN2DL port map( A1 => n391, A2 => n382, Z => n990);
   U1010 : NAN2DL port map( A1 => n382, A2 => n384, Z => n991);
   U1011 : NAN2DL port map( A1 => n391, A2 => n384, Z => n992);
   U1012 : NAN3D2 port map( A1 => n990, A2 => n991, A3 => n992, Z => n377);
   U1013 : EXOR3D1 port map( A1 => n368, A2 => n377, A3 => n1064, Z => n1065);
   U1014 : EXNOR2D2 port map( A1 => b(13), A2 => a(5), Z => n736);
   U1015 : EXNOR2D2 port map( A1 => b(14), A2 => a(5), Z => n735);
   U1016 : BUFDL port map( A => n680, Z => n994);
   U1017 : EXNOR2D1 port map( A1 => b(1), A2 => a(13), Z => n680);
   U1018 : NAN2D1 port map( A1 => n354, A2 => n363, Z => n173);
   U1019 : EXNOR2D2 port map( A1 => b(2), A2 => a(11), Z => n696);
   U1020 : AOI21DL port map( A1 => n202, A2 => n288, B => n199, Z => n197);
   U1021 : EXNOR2D2 port map( A1 => b(10), A2 => a(3), Z => n756);
   U1022 : EXNOR2D2 port map( A1 => b(2), A2 => a(13), Z => n679);
   U1023 : EXNOR2DL port map( A1 => b(2), A2 => a(9), Z => n713);
   U1024 : EXNOR2D1 port map( A1 => b(10), A2 => a(1), Z => n773);
   U1025 : EXOR2D1 port map( A1 => n539, A2 => n569, Z => n1029);
   U1026 : EXOR3D1 port map( A1 => n449, A2 => n590, A3 => n905, Z => n436);
   U1027 : NAN2D1 port map( A1 => n605, A2 => n449, Z => n996);
   U1028 : NAN2D1 port map( A1 => n605, A2 => n590, Z => n997);
   U1029 : NAN3D2 port map( A1 => n997, A2 => n996, A3 => n995, Z => n435);
   U1030 : EXOR2D1 port map( A1 => n619, A2 => n437, Z => n998);
   U1031 : NAN2D1 port map( A1 => n902, A2 => n437, Z => n999);
   U1032 : NAN2D1 port map( A1 => n902, A2 => n435, Z => n1000);
   U1033 : NAN2D1 port map( A1 => n437, A2 => n435, Z => n1001);
   U1034 : EXNOR2DL port map( A1 => b(7), A2 => a(5), Z => n742);
   U1035 : EXNOR2DL port map( A1 => b(11), A2 => a(7), Z => n721);
   U1036 : EXNOR2D2 port map( A1 => b(5), A2 => a(7), Z => n727);
   U1037 : OA21DL port map( A1 => n217, A2 => n223, B => n1027, Z => n214);
   U1038 : OAI21DL port map( A1 => n934, A2 => n108, B => n109, Z => n107);
   U1039 : INVDL port map( A => n52, Z => n129);
   U1040 : EXNOR2D2 port map( A1 => b(3), A2 => a(15), Z => n661);
   U1041 : EXNOR2D2 port map( A1 => b(3), A2 => a(1), Z => n780);
   U1042 : EXNOR2D2 port map( A1 => b(3), A2 => a(5), Z => n746);
   U1043 : EXNOR2DL port map( A1 => b(3), A2 => a(7), Z => n729);
   U1044 : EXNOR2D2 port map( A1 => b(3), A2 => a(9), Z => n712);
   U1045 : EXNOR2DL port map( A1 => b(3), A2 => a(13), Z => n678);
   U1046 : EXNOR2DL port map( A1 => b(2), A2 => a(1), Z => n781);
   U1047 : EXNOR2DL port map( A1 => b(2), A2 => a(3), Z => n764);
   U1048 : EXNOR2DL port map( A1 => b(2), A2 => a(5), Z => n747);
   U1049 : NAN2D1 port map( A1 => n288, A2 => n1066, Z => n67);
   U1050 : NAN3D1 port map( A1 => n1014, A2 => n1016, A3 => n1015, Z => n457);
   U1051 : EXNOR2DL port map( A1 => b(2), A2 => a(7), Z => n730);
   U1052 : OAI22D1 port map( A1 => n758, A2 => n12, B1 => n757, B2 => n9, Z => 
                           n623);
   U1053 : EXOR2D1 port map( A1 => n443, A2 => n434, Z => n1003);
   U1054 : EXOR2D1 port map( A1 => n1003, A2 => n432, Z => n430);
   U1055 : NAN2DL port map( A1 => n432, A2 => n434, Z => n1004);
   U1056 : NAN2DL port map( A1 => n432, A2 => n443, Z => n1005);
   U1057 : NAN3D1 port map( A1 => n1004, A2 => n1006, A3 => n1005, Z => n429);
   U1058 : EXOR3DL port map( A1 => n417, A2 => n406, A3 => n404, Z => n1051);
   U1059 : EXOR3D1 port map( A1 => n616, A2 => n393, A3 => n395, Z => n380);
   U1060 : INVDL port map( A => b(9), Z => n1007);
   U1061 : INVDL port map( A => n1007, Z => n1008);
   U1062 : AOI21D1 port map( A1 => n1020, A2 => n952, B => n1033, Z => n160);
   U1063 : OR2D2 port map( A1 => n474, A2 => n481, Z => n1077);
   U1064 : EXOR2D1 port map( A1 => n420, A2 => n431, Z => n1009);
   U1065 : NAN2DL port map( A1 => n418, A2 => n431, Z => n1010);
   U1066 : NAN2D1 port map( A1 => n418, A2 => n420, Z => n1011);
   U1067 : NAN2DL port map( A1 => n431, A2 => n420, Z => n1012);
   U1068 : NAN3D1 port map( A1 => n1010, A2 => n1012, A3 => n1011, Z => n415);
   U1069 : NAN2D1 port map( A1 => n1052, A2 => n415, Z => n1066);
   U1070 : NOR2D1 port map( A1 => n1051, A2 => n415, Z => n200);
   U1071 : NAN2DL port map( A1 => n622, A2 => n607, Z => n1014);
   U1072 : NAN2DL port map( A1 => n622, A2 => n469, Z => n1015);
   U1073 : NAN2DL port map( A1 => n607, A2 => n469, Z => n1016);
   U1074 : OAI22D1 port map( A1 => n742, A2 => n18, B1 => n741, B2 => n16, Z =>
                           n607);
   U1075 : EXNOR2D2 port map( A1 => n105, A2 => n1017, Z => product(27));
   U1076 : ADHALFD2 port map( A => n546, B => n514, CO => n451, S => n452);
   U1077 : NAN2DL port map( A1 => n286, A2 => n187, Z => n65);
   U1078 : EXNOR2D2 port map( A1 => b(10), A2 => a(5), Z => n1060);
   U1079 : NOR2D2 port map( A1 => n344, A2 => n353, Z => n167);
   U1080 : EXOR2D4 port map( A1 => n197, A2 => n66, Z => product(17));
   U1081 : INVDL port map( A => n1020, Z => n1018);
   U1082 : INVDL port map( A => n1018, Z => n1019);
   U1083 : EXNOR2D2 port map( A1 => b(12), A2 => a(9), Z => n703);
   U1084 : BUFD4 port map( A => n51, Z => n1020);
   U1085 : EXNOR2D2 port map( A1 => n1059, A2 => a(7), Z => n718);
   U1086 : OAI21D1 port map( A1 => n175, A2 => n203, B => n176, Z => n51);
   U1087 : OR2D2 port map( A1 => n322, A2 => n327, Z => n1078);
   U1088 : NAN2DL port map( A1 => n403, A2 => n390, Z => n1021);
   U1089 : NAN2DL port map( A1 => n403, A2 => n392, Z => n1022);
   U1090 : NAN2DL port map( A1 => n392, A2 => n390, Z => n1023);
   U1091 : NAN3D1 port map( A1 => n1021, A2 => n1023, A3 => n1022, Z => n387);
   U1092 : NAN2DL port map( A1 => n419, A2 => n410, Z => n1025);
   U1093 : NAN2D1 port map( A1 => n408, A2 => n410, Z => n1026);
   U1094 : OAI21D1 port map( A1 => n210, A2 => n206, B => n207, Z => n205);
   U1095 : NAN2DL port map( A1 => n453, A2 => n442, Z => n1027);
   U1096 : EXNOR2D2 port map( A1 => n1042, A2 => a(3), Z => n759);
   U1097 : INVD1 port map( A => n1041, Z => n1042);
   U1098 : OAI22D1 port map( A1 => n769, A2 => n6, B1 => n768, B2 => n824, Z =>
                           n634);
   U1099 : EXNOR2D2 port map( A1 => n1059, A2 => a(9), Z => n701);
   U1100 : BUFD1 port map( A => b(14), Z => n1059);
   U1101 : EXNOR2DL port map( A1 => b(9), A2 => a(7), Z => n723);
   U1102 : NAN2D1 port map( A1 => n189, A2 => n177, Z => n175);
   U1103 : OAI22D2 port map( A1 => n6, A2 => n773, B1 => n772, B2 => n824, Z =>
                           n638);
   U1104 : NAN2DL port map( A1 => n584, A2 => n569, Z => n1030);
   U1105 : NAN2DL port map( A1 => n584, A2 => n539, Z => n1031);
   U1106 : NAN2DL port map( A1 => n569, A2 => n539, Z => n1032);
   U1107 : NAN3D1 port map( A1 => n1030, A2 => n1032, A3 => n1031, Z => n359);
   U1108 : OAI22DL port map( A1 => n674, A2 => n42, B1 => n673, B2 => n40, Z =>
                           n539);
   U1109 : INVDL port map( A => n164, Z => n1033);
   U1110 : OAI21D1 port map( A1 => n211, A2 => n209, B => n210, Z => n208);
   U1111 : EXOR3D2 port map( A1 => n574, A2 => n439, A3 => n589, Z => n424);
   U1112 : NAN2D1 port map( A1 => n574, A2 => n589, Z => n1035);
   U1113 : NAN2D1 port map( A1 => n439, A2 => n589, Z => n1036);
   U1114 : NAN3D2 port map( A1 => n1034, A2 => n1035, A3 => n1036, Z => n423);
   U1115 : NAN2DL port map( A1 => n633, A2 => n423, Z => n1039);
   U1116 : EXNOR2DL port map( A1 => b(7), A2 => a(9), Z => n708);
   U1117 : EXNOR2D2 port map( A1 => b(3), A2 => a(11), Z => n695);
   U1118 : EXNOR2D2 port map( A1 => b(12), A2 => a(7), Z => n720);
   U1119 : EXNOR2DL port map( A1 => b(12), A2 => a(11), Z => n686);
   U1120 : EXNOR2DL port map( A1 => n932, A2 => a(13), Z => n669);
   U1121 : EXNOR2DL port map( A1 => n932, A2 => a(15), Z => n652);
   U1122 : EXOR2D2 port map( A1 => n114, A2 => n57, Z => product(26));
   U1123 : EXOR2D4 port map( A1 => n188, A2 => n65, Z => product(18));
   U1124 : NAN2D1 port map( A1 => n396, A2 => n409, Z => n1043);
   U1125 : NAN2D1 port map( A1 => n409, A2 => n617, Z => n1044);
   U1126 : NAN2D1 port map( A1 => n396, A2 => n617, Z => n1045);
   U1127 : NAN3D2 port map( A1 => n1043, A2 => n1045, A3 => n1044, Z => n391);
   U1128 : NAN2D1 port map( A1 => n573, A2 => n425, Z => n1048);
   U1129 : OAI22D2 port map( A1 => n752, A2 => n12, B1 => n751, B2 => n9, Z => 
                           n617);
   U1130 : EXOR2D4 port map( A1 => n211, A2 => n69, Z => product(14));
   U1131 : AOI21D1 port map( A1 => n115, A2 => n1020, B => n116, Z => n114);
   U1132 : EXNOR2D2 port map( A1 => n169, A2 => n1049, Z => product(21));
   U1133 : AND2DL port map( A1 => n283, A2 => n168, Z => n1049);
   U1134 : EXNOR2DL port map( A1 => b(8), A2 => a(13), Z => n673);
   U1135 : EXNOR2DL port map( A1 => a(1), A2 => b(8), Z => n775);
   U1136 : EXNOR2DL port map( A1 => b(8), A2 => a(3), Z => n758);
   U1137 : EXOR3DL port map( A1 => n417, A2 => n966, A3 => n404, Z => n1052);
   U1138 : OAI22D1 port map( A1 => n769, A2 => n6, B1 => n768, B2 => n824, Z =>
                           n1053);
   U1139 : EXNOR2D2 port map( A1 => b(15), A2 => a(1), Z => n768);
   U1140 : ADFULD1 port map( A => n544, B => n428, CI => n559, CO => n425, S =>
                           n426);
   U1141 : NOR2D2 port map( A1 => n179, A2 => n184, Z => n177);
   U1142 : EXNOR2DL port map( A1 => n1042, A2 => a(1), Z => n776);
   U1143 : EXNOR2DL port map( A1 => b(7), A2 => a(15), Z => n657);
   U1144 : EXNOR2DL port map( A1 => b(7), A2 => a(13), Z => n674);
   U1145 : EXNOR2D2 port map( A1 => b(7), A2 => a(7), Z => n725);
   U1146 : NAN2D1 port map( A1 => n393, A2 => n395, Z => n1054);
   U1147 : NAN2D1 port map( A1 => n395, A2 => n616, Z => n1056);
   U1148 : NAN3D2 port map( A1 => n1054, A2 => n1055, A3 => n1056, Z => n379);
   U1149 : AO21D1 port map( A1 => n12, A2 => n9, B => n751, Z => n616);
   U1150 : AOI21DL port map( A1 => n1019, A2 => n86, B => n87, Z => n85);
   U1151 : EXNOR2DL port map( A1 => n1020, A2 => n63, Z => product(20));
   U1152 : EXNOR2D2 port map( A1 => b(5), A2 => a(13), Z => n676);
   U1153 : EXNOR2D2 port map( A1 => b(2), A2 => a(15), Z => n662);
   U1154 : OR2D2 port map( A1 => n529, A2 => n427, Z => n413);
   U1155 : EXNOR2D2 port map( A1 => n1082, A2 => n378, Z => n376);
   U1156 : INVDL port map( A => n910, Z => n285);
   U1157 : EXNOR2D2 port map( A1 => b(10), A2 => a(7), Z => n722);
   U1158 : EXNOR2D2 port map( A1 => n127, A2 => n1075, Z => product(25));
   U1159 : INVDL port map( A => n192, Z => n1057);
   U1160 : BUFDL port map( A => n379, Z => n1058);
   U1161 : EXNOR2DL port map( A1 => b(9), A2 => a(15), Z => n655);
   U1162 : EXNOR2DL port map( A1 => b(9), A2 => a(1), Z => n774);
   U1163 : NAN2D1 port map( A1 => n426, A2 => n901, Z => n1061);
   U1164 : NAN2D1 port map( A1 => n1053, A2 => n901, Z => n1062);
   U1165 : NAN2D1 port map( A1 => n1053, A2 => n426, Z => n1063);
   U1166 : NAN3D2 port map( A1 => n1062, A2 => n1063, A3 => n1061, Z => n421);
   U1167 : EXOR3DL port map( A1 => n381, A2 => n370, A3 => n1058, Z => n1064);
   U1168 : EXNOR2DL port map( A1 => b(6), A2 => a(3), Z => n760);
   U1169 : EXNOR2DL port map( A1 => b(6), A2 => a(5), Z => n743);
   U1170 : EXNOR2DL port map( A1 => b(6), A2 => a(1), Z => n777);
   U1171 : NAN2D1 port map( A1 => n402, A2 => n415, Z => n201);
   U1172 : EXNOR2D2 port map( A1 => b(5), A2 => a(11), Z => n693);
   U1173 : EXNOR2D2 port map( A1 => b(6), A2 => a(11), Z => n692);
   U1174 : EXNOR2D2 port map( A1 => b(5), A2 => a(9), Z => n710);
   U1175 : NOR2D2 port map( A1 => n416, A2 => n429, Z => n206);
   U1176 : EXNOR2D2 port map( A1 => b(14), A2 => a(1), Z => n769);
   U1177 : OAI22D1 port map( A1 => n947, A2 => n18, B1 => n737, B2 => n16, Z =>
                           n603);
   U1178 : EXNOR2D2 port map( A1 => b(12), A2 => a(5), Z => n737);
   U1179 : NOR2DL port map( A1 => n53, A2 => n108, Z => n106);
   U1180 : NOR2D1 port map( A1 => n1028, A2 => n167, Z => n161);
   U1181 : NAN2DL port map( A1 => n101, A2 => n279, Z => n97);
   U1182 : AOI21DL port map( A1 => n106, A2 => n1020, B => n107, Z => n105);
   U1183 : AND2D1 port map( A1 => n482, A2 => n489, Z => n1072);
   U1184 : NOR2D1 port map( A1 => n506, A2 => n509, Z => n257);
   U1185 : OR2D1 port map( A1 => n510, A2 => n645, Z => n1086);
   U1186 : INVDL port map( A => n319, Z => n320);
   U1187 : AND2DL port map( A1 => n281, A2 => n150, Z => n1073);
   U1188 : EXNOR2D2 port map( A1 => n151, A2 => n1073, Z => product(23));
   U1189 : AND2DL port map( A1 => n282, A2 => n155, Z => n1074);
   U1190 : EXNOR2D2 port map( A1 => n160, A2 => n1074, Z => product(22));
   U1191 : EXNOR2D1 port map( A1 => n1067, A2 => n1076, Z => product(19));
   U1192 : AOI21DL port map( A1 => n182, A2 => n202, B => n183, Z => n1067);
   U1193 : NAN2M1DL port map( A1 => n913, A2 => n196, Z => n66);
   U1194 : AOI21M10DL port map( A1 => n155, A2 => n281, B => n148, Z => n144);
   U1195 : INVDL port map( A => n1028, Z => n284);
   U1196 : NAN2D2 port map( A1 => n281, A2 => n1078, Z => n134);
   U1197 : INVD2 port map( A => n117, Z => n279);
   U1198 : NAN2DL port map( A1 => n278, A2 => n113, Z => n57);
   U1199 : NAN2M1DL port map( A1 => n103, A2 => n104, Z => n56);
   U1200 : NAN2M1DL port map( A1 => n206, A2 => n207, Z => n68);
   U1201 : OAI21D1 port map( A1 => n1068, A2 => n243, B => n232, Z => n230);
   U1202 : EXOR2D1 port map( A1 => n1069, A2 => n1070, Z => product(28));
   U1203 : AOI21DL port map( A1 => n1019, A2 => n95, B => n96, Z => n1069);
   U1204 : NAN2DL port map( A1 => n276, A2 => n93, Z => n1070);
   U1205 : NAN2DL port map( A1 => n322, A2 => n327, Z => n139);
   U1206 : INVD1 port map( A => n112, Z => n278);
   U1207 : NAN2DL port map( A1 => n416, A2 => n429, Z => n207);
   U1208 : OR2D1 port map( A1 => n490, A2 => n495, Z => n1071);
   U1209 : AND2DL port map( A1 => n502, A2 => n505, Z => n1085);
   U1210 : OAI22DL port map( A1 => n688, A2 => n36, B1 => n687, B2 => n34, Z =>
                           n553);
   U1211 : OAI22DL port map( A1 => n684, A2 => n36, B1 => n683, B2 => n34, Z =>
                           n549);
   U1212 : OAI22DL port map( A1 => n653, A2 => n48, B1 => n652, B2 => n46, Z =>
                           n524);
   U1213 : OAI22DL port map( A1 => n652, A2 => n48, B1 => n651, B2 => n46, Z =>
                           n523);
   U1214 : OA22DL port map( A1 => n650, A2 => n48, B1 => n649, B2 => n46, Z => 
                           n1092);
   U1215 : NOR2DL port map( A1 => n53, A2 => n97, Z => n95);
   U1216 : INVDL port map( A => n184, Z => n286);
   U1217 : NOR2D1 port map( A1 => n200, A2 => n913, Z => n189);
   U1218 : OA21M20D1 port map( A1 => n148, A2 => n1078, B => n139, Z => n135);
   U1219 : AND2D1 port map( A1 => n279, A2 => n118, Z => n1075);
   U1220 : AND2DL port map( A1 => n285, A2 => n180, Z => n1076);
   U1221 : NOR2D1 port map( A1 => n163, A2 => n143, Z => n141);
   U1222 : NAN2DL port map( A1 => n284, A2 => n173, Z => n63);
   U1223 : INVDL port map( A => n200, Z => n288);
   U1224 : NOR2M1DL port map( A1 => n912, A2 => n914, Z => n182);
   U1225 : NAN2D1 port map( A1 => n282, A2 => n281, Z => n143);
   U1226 : INVDL port map( A => n154, Z => n282);
   U1227 : NOR2DL port map( A1 => n53, A2 => n1081, Z => n86);
   U1228 : NAN2D1 port map( A1 => n279, A2 => n278, Z => n108);
   U1229 : NOR2D1 port map( A1 => n53, A2 => n117, Z => n115);
   U1230 : OA21M20D1 port map( A1 => n960, A2 => n278, B => n113, Z => n109);
   U1231 : INVD2 port map( A => n149, Z => n281);
   U1232 : NAN2D1 port map( A1 => n328, A2 => n335, Z => n150);
   U1233 : NAN2D1 port map( A1 => n344, A2 => n353, Z => n168);
   U1234 : NAN2D1 port map( A1 => n336, A2 => n343, Z => n155);
   U1235 : AND2D1 port map( A1 => n464, A2 => n473, Z => n1079);
   U1236 : OA21DL port map( A1 => n100, A2 => n92, B => n93, Z => n1080);
   U1237 : NAN2D1 port map( A1 => n316, A2 => n321, Z => n118);
   U1238 : OR2D1 port map( A1 => n97, A2 => n92, Z => n1081);
   U1239 : NOR2D1 port map( A1 => n112, A2 => n103, Z => n101);
   U1240 : EXNOR2D1 port map( A1 => n380, A2 => n389, Z => n1082);
   U1241 : NAN2D1 port map( A1 => n430, A2 => n441, Z => n210);
   U1242 : AND2D1 port map( A1 => n490, A2 => n495, Z => n1083);
   U1243 : NAN2DL port map( A1 => n496, A2 => n501, Z => n250);
   U1244 : NOR2DL port map( A1 => n496, A2 => n501, Z => n249);
   U1245 : OR2D1 port map( A1 => n502, A2 => n505, Z => n1084);
   U1246 : NAN2DL port map( A1 => n506, A2 => n509, Z => n258);
   U1247 : AND2D1 port map( A1 => n510, A2 => n645, Z => n1087);
   U1248 : OR2D1 port map( A1 => n647, A2 => n632, Z => n1088);
   U1249 : AND2D1 port map( A1 => n647, A2 => n632, Z => n1089);
   U1250 : NAN2D1 port map( A1 => n312, A2 => n315, Z => n113);
   U1251 : NAN2DL port map( A1 => n311, A2 => n308, Z => n104);
   U1252 : NAN2DL port map( A1 => n307, A2 => n306, Z => n93);
   U1253 : AO21D1 port map( A1 => n6, A2 => n824, B => n768, Z => n633);
   U1254 : AO21D1 port map( A1 => n18, A2 => n16, B => n734, Z => n599);
   U1255 : INVD2 port map( A => n373, Z => n374);
   U1256 : INVD2 port map( A => n351, Z => n352);
   U1257 : INVD2 port map( A => n333, Z => n334);
   U1258 : NAN2D1 port map( A1 => n1091, A2 => n84, Z => n54);
   U1259 : NAN2DL port map( A1 => n305, A2 => n1092, Z => n84);
   U1260 : AO21D1 port map( A1 => n36, A2 => n34, B => n683, Z => n548);
   U1261 : NAN2DL port map( A1 => n646, A2 => n512, Z => n266);
   U1262 : NOR2DL port map( A1 => n646, A2 => n512, Z => n265);
   U1263 : AND2D1 port map( A1 => n648, A2 => n520, Z => n1090);
   U1264 : INVD2 port map( A => n309, Z => n310);
   U1265 : AO21D1 port map( A1 => n42, A2 => n40, B => n666, Z => n532);
   U1266 : OR2D1 port map( A1 => n305, A2 => n1092, Z => n1091);
   U1267 : INVD1 port map( A => a(13), Z => n826);
   U1268 : INVD1 port map( A => a(15), Z => n825);
   U1269 : INVD1 port map( A => a(11), Z => n827);
   U1270 : INVD1 port map( A => a(9), Z => n828);
   U1271 : INVD1 port map( A => a(7), Z => n829);
   U1272 : INVD1 port map( A => a(5), Z => n830);
   U1273 : ADHALFDL port map( A => n631, B => n519, CO => n511, S => n512);
   U1274 : INVD1 port map( A => a(3), Z => n831);
   U1275 : EXNOR2D1 port map( A1 => a(13), A2 => a(14), Z => n46);
   U1276 : NAN2D1 port map( A1 => n801, A2 => n46, Z => n48);
   U1277 : EXNOR2D1 port map( A1 => a(11), A2 => a(12), Z => n40);
   U1278 : NAN2D1 port map( A1 => n802, A2 => n40, Z => n42);
   U1279 : EXNOR2D1 port map( A1 => a(9), A2 => a(10), Z => n34);
   U1280 : NAN2D1 port map( A1 => n803, A2 => n34, Z => n36);
   U1281 : EXNOR2D1 port map( A1 => a(7), A2 => a(8), Z => n28);
   U1282 : NAN2D1 port map( A1 => n804, A2 => n28, Z => n30);
   U1283 : EXNOR2D1 port map( A1 => a(5), A2 => a(6), Z => n22);
   U1284 : NAN2D1 port map( A1 => n805, A2 => n22, Z => n24);
   U1285 : EXNOR2D1 port map( A1 => a(1), A2 => a(2), Z => n9);
   U1286 : NAN2D1 port map( A1 => n807, A2 => n9, Z => n12);
   U1287 : EXNOR2D1 port map( A1 => a(3), A2 => a(4), Z => n16);
   U1288 : NAN2D1 port map( A1 => n806, A2 => n16, Z => n18);
   U1289 : NAN2D1 port map( A1 => n808, A2 => n824, Z => n6);
   U1290 : INVD1 port map( A => a(0), Z => n824);
   U1291 : INVD1 port map( A => a(1), Z => n832);
   U1292 : EXNOR2DL port map( A1 => b(1), A2 => a(1), Z => n782);
   U1293 : EXNOR2DL port map( A1 => b(1), A2 => a(3), Z => n765);
   U1294 : EXNOR2DL port map( A1 => b(1), A2 => a(5), Z => n748);
   U1295 : EXNOR2DL port map( A1 => b(1), A2 => a(7), Z => n731);
   U1296 : EXNOR2DL port map( A1 => b(1), A2 => a(9), Z => n714);
   U1297 : OAI21DL port map( A1 => n192, A2 => n914, B => n187, Z => n183);
   U1298 : INVD1 port map( A => n212, Z => n211);
   U1299 : INVDL port map( A => n954, Z => n192);
   U1300 : OAI22D1 port map( A1 => n771, A2 => n6, B1 => n770, B2 => n824, Z =>
                           n636);
   U1301 : EXNOR2DL port map( A1 => b(5), A2 => a(1), Z => n778);
   U1302 : EXNOR2DL port map( A1 => b(5), A2 => a(3), Z => n761);
   U1303 : EXNOR2DL port map( A1 => b(5), A2 => a(15), Z => n659);
   U1304 : OAI21DL port map( A1 => n52, A2 => n1081, B => n1080, Z => n87);
   U1305 : OAI21DL port map( A1 => n934, A2 => n97, B => n100, Z => n96);
   U1306 : EXNOR2DL port map( A1 => b(15), A2 => a(15), Z => n649);
   U1307 : OAI22M10D1 port map( A1 => a(0), A2 => n769, B1 => n770, B2 => n6, Z
                           => n635);
   U1308 : EXNOR2DL port map( A1 => b(10), A2 => a(15), Z => n654);
   U1309 : EXNOR2DL port map( A1 => b(10), A2 => a(13), Z => n671);
   U1310 : EXNOR2DL port map( A1 => n1059, A2 => a(15), Z => n650);
   U1311 : EXNOR2DL port map( A1 => a(13), A2 => n1059, Z => n667);
   U1312 : EXNOR2DL port map( A1 => n1059, A2 => a(11), Z => n684);
   U1313 : INVDL port map( A => n1066, Z => n199);
   U1314 : NAN2DL port map( A1 => n389, A2 => n378, Z => n1093);
   U1315 : NAN2DL port map( A1 => n378, A2 => n380, Z => n1094);
   U1316 : NAN2D1 port map( A1 => n1065, A2 => n375, Z => n180);
   U1317 : AOI21DL port map( A1 => n128, A2 => n1020, B => n129, Z => n127);
   U1318 : AOI21DL port map( A1 => n1020, A2 => n152, B => n153, Z => n151);
   U1319 : NAN2D1 port map( A1 => n909, A2 => n401, Z => n196);
   U1320 : EXNOR2DL port map( A1 => b(13), A2 => a(15), Z => n651);
   U1321 : EXNOR2DL port map( A1 => b(13), A2 => a(13), Z => n668);
   U1322 : EXNOR2DL port map( A1 => b(13), A2 => a(11), Z => n685);
   U1323 : EXNOR2DL port map( A1 => b(13), A2 => a(9), Z => n702);
   U1324 : EXNOR2DL port map( A1 => b(13), A2 => a(7), Z => n719);
   U1325 : AOI21DL port map( A1 => n202, A2 => n968, B => n1057, Z => n188);
   U1326 : EXNOR2DL port map( A1 => b(11), A2 => a(15), Z => n653);
   U1327 : EXNOR2DL port map( A1 => b(11), A2 => a(13), Z => n670);
   U1328 : EXNOR2DL port map( A1 => b(11), A2 => a(11), Z => n687);
   U1329 : EXNOR2DL port map( A1 => b(11), A2 => a(1), Z => n772);

end hier_sec_par_16_5;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_siso_gen.all;

architecture hier_sec_par_16_5 of siso_gen_DW_mult_tc_17 is

   component EXNOR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INVDL
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AO21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OA22DL
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22DL
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component NAN3D2
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22D2
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFD2
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component EXOR2D4
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR3D2
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR3DL
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFDL
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21M10DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AO21D2
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADFULD2
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component INVBD2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21M20DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFD1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component AOI22M10D1
      port( B1, B2, A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22D4
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21M20DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21M10D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component ADFULDL
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component NOR2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   signal n6, n9, n12, n16, n18, n22, n24, n28, n30, n34, n36, n40, n42, n46, 
      n48, n52, n53, n54, n55, n56, n63, n65, n67, n68, n69, n84, n85, n86, n87
      , n92, n93, n94, n95, n96, n97, n100, n101, n102, n103, n104, n105, n106,
      n107, n108, n109, n112, n113, n114, n115, n116, n117, n118, n124, n127, 
      n128, n129, n135, n139, n140, n141, n142, n148, n160, n167, n168, n169, 
      n171, n172, n173, n182, n183, n188, n192, n195, n196, n197, n199, n200, 
      n201, n202, n206, n207, n208, n209, n210, n211, n212, n213, n214, n225, 
      n230, n231, n232, n243, n248, n249, n250, n251, n256, n257, n258, n259, 
      n264, n265, n266, n267, n278, n279, n283, n284, n285, n287, n288, n305, 
      n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, 
      n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, 
      n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, 
      n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, 
      n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, 
      n366, n367, n368, n369, n370, n371, n372, n373, n374, n379, n381, n382, 
      n383, n385, n386, n388, n393, n394, n397, n398, n399, n400, n401, n402, 
      n403, n404, n407, n408, n410, n413, n415, n416, n417, n418, n419, n420, 
      n422, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, 
      n436, n437, n438, n441, n442, n443, n444, n445, n446, n447, n448, n449, 
      n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, 
      n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, 
      n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, 
      n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, 
      n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, 
      n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n522, 
      n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n544, n546, n547, n548, 
      n549, n550, n551, n552, n553, n554, n555, n556, n559, n560, n561, n562, 
      n563, n564, n565, n566, n567, n568, n569, n570, n571, n573, n574, n575, 
      n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, 
      n588, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, 
      n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, 
      n613, n614, n615, n616, n618, n619, n620, n621, n622, n623, n624, n625, 
      n626, n627, n628, n629, n630, n631, n632, n635, n636, n637, n638, n639, 
      n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, 
      n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, 
      n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, 
      n676, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, 
      n690, n691, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, 
      n704, n705, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, 
      n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, 
      n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, 
      n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, 
      n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, 
      n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, 
      n778, n779, n780, n781, n782, n783, n784, n801, n805, n806, n807, n808, 
      n824, n826, n827, n828, n829, n830, n831, n832, net11025, net11083, 
      net11172, net11509, net11507, net11503, net11662, net11667, net11666, 
      net11693, net11746, net11745, net11829, net12033, net12055, net12054, 
      net12079, net12078, net12095, net12127, net12126, net12125, net12153, 
      net12152, net12151, net12183, net12250, net12249, net12257, net12285, 
      n804, net12065, n205, n204, n203, n187, n180, n384, n380, n378, n377, n51
      , n161, n132, net11587, net11586, net11585, n387, n802, n678, n677, n803,
      n707, n693, n692, n617, n572, n558, n557, n543, n414, n412, n411, n409, 
      n396, n395, n392, n391, n634, n633, n589, n545, n440, n439, n424, n423, 
      n421, n406, n405, n390, n389, net12019, n376, n375, n184, n179, net11675,
      net11621, net11096, net10037, n282, n164, n163, n162, n155, n154, n153, 
      n152, n151, n150, n144, n143, n134, n189, n178, n177, n176, n175, n706, 
      n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, 
      n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, 
      n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, 
      n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, 
      n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, 
      n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, 
      n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, 
      n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, 
      n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, 
      n1007, n1008, n1009, n1010, n1011, n1012, n1013, n_1033 : std_logic;

begin
   
   U54 : EXOR2D1 port map( A1 => n85, A2 => n54, Z => product(29));
   U59 : EXOR2D1 port map( A1 => n94, A2 => n55, Z => product(28));
   U78 : AOI21D1 port map( A1 => n101, A2 => n124, B => n102, Z => n100);
   U80 : OAI21D1 port map( A1 => n113, A2 => n103, B => n104, Z => n102);
   U114 : AOI21D1 port map( A1 => net12285, A2 => n128, B => n129, Z => n127);
   U165 : NOR2D2 port map( A1 => n344, A2 => n353, Z => n167);
   U205 : NOR2D2 port map( A1 => n388, A2 => n401, Z => n195);
   U207 : EXNOR2D1 port map( A1 => n202, A2 => n67, Z => product(16));
   U222 : NOR2D2 port map( A1 => n416, A2 => n429, Z => n206);
   U224 : EXOR2D1 port map( A1 => n211, A2 => n69, Z => product(14));
   U228 : NOR2D2 port map( A1 => n430, A2 => n441, Z => n209);
   U232 : OAI21D1 port map( A1 => n225, A2 => n213, B => n214, Z => n212);
   U234 : AOI21D1 port map( A1 => n990, A2 => n992, B => n994, Z => n214);
   U259 : OAI21D1 port map( A1 => n231, A2 => n243, B => n232, Z => n230);
   U278 : AOI21D1 port map( A1 => n248, A2 => n1000, B => n1001, Z => n243);
   U286 : OAI21D1 port map( A1 => n249, A2 => n251, B => n250, Z => n248);
   U292 : AOI21D1 port map( A1 => n256, A2 => n1002, B => n1003, Z => n251);
   U300 : OAI21D1 port map( A1 => n257, A2 => n259, B => n258, Z => n256);
   U306 : AOI21D1 port map( A1 => n1004, A2 => n264, B => n1005, Z => n259);
   U314 : OAI21D1 port map( A1 => n267, A2 => n265, B => n266, Z => n264);
   U320 : AOI21D1 port map( A1 => n1006, A2 => n1008, B => n1007, Z => n267);
   U334 : ADFULD1 port map( A => n522, B => n309, CI => n532, CO => n305, S => 
                           n306);
   U335 : ADFULD1 port map( A => n310, B => n523, CI => n313, CO => n307, S => 
                           n308);
   U337 : ADFULD1 port map( A => n317, B => n533, CI => n314, CO => n311, S => 
                           n312);
   U338 : ADFULD1 port map( A => n524, B => n319, CI => n548, CO => n313, S => 
                           n314);
   U339 : ADFULD1 port map( A => n318, B => n325, CI => n323, CO => n315, S => 
                           n316);
   U340 : ADFULD1 port map( A => n534, B => n549, CI => n320, CO => n317, S => 
                           n318);
   U342 : ADFULD1 port map( A => n329, B => n326, CI => n324, CO => n321, S => 
                           n322);
   U343 : ADFULD1 port map( A => n565, B => n535, CI => n331, CO => n323, S => 
                           n324);
   U344 : ADFULD1 port map( A => n333, B => n525, CI => n550, CO => n325, S => 
                           n326);
   U345 : ADFULD1 port map( A => n337, B => n332, CI => n330, CO => n327, S => 
                           n328);
   U346 : ADFULD1 port map( A => n341, B => n566, CI => n339, CO => n329, S => 
                           n330);
   U347 : ADFULD1 port map( A => n536, B => n334, CI => n551, CO => n331, S => 
                           n332);
   U349 : ADFULD1 port map( A => n345, B => n340, CI => n338, CO => n335, S => 
                           n336);
   U350 : ADFULD1 port map( A => n342, B => n349, CI => n347, CO => n337, S => 
                           n338);
   U351 : ADFULD1 port map( A => n567, B => n552, CI => n582, CO => n339, S => 
                           n340);
   U352 : ADFULD1 port map( A => n537, B => n351, CI => n526, CO => n341, S => 
                           n342);
   U353 : ADFULD1 port map( A => n355, B => n348, CI => n346, CO => n343, S => 
                           n344);
   U354 : ADFULD1 port map( A => n350, B => n359, CI => n357, CO => n345, S => 
                           n346);
   U355 : ADFULD1 port map( A => n568, B => n583, CI => n361, CO => n347, S => 
                           n348);
   U356 : ADFULD1 port map( A => n352, B => n538, CI => n553, CO => n349, S => 
                           n350);
   U358 : ADFULD1 port map( A => n365, B => n358, CI => n356, CO => n353, S => 
                           n354);
   U359 : ADFULD1 port map( A => n360, B => n369, CI => n367, CO => n355, S => 
                           n356);
   U360 : ADFULD1 port map( A => n371, B => n599, CI => n362, CO => n357, S => 
                           n358);
   U361 : ADFULD1 port map( A => n569, B => n539, CI => n584, CO => n359, S => 
                           n360);
   U362 : ADFULD1 port map( A => n527, B => n373, CI => n554, CO => n361, S => 
                           n362);
   U365 : ADFULD1 port map( A => n383, B => n585, CI => n372, CO => n367, S => 
                           n368);
   U366 : ADFULD1 port map( A => n570, B => n385, CI => n600, CO => n369, S => 
                           n370);
   U367 : ADFULD1 port map( A => n540, B => n374, CI => n555, CO => n371, S => 
                           n372);
   U372 : ADFULD1 port map( A => n386, B => n586, CI => n601, CO => n381, S => 
                           n382);
   U374 : ADFULD1 port map( A => n528, B => n399, CI => n541, CO => n385, S => 
                           n386);
   U378 : ADFULD1 port map( A => n398, B => n587, CI => n602, CO => n393, S => 
                           n394);
   U380 : ADFULD1 port map( A => n400, B => n413, CI => n542, CO => n397, S => 
                           n398);
   U390 : ADFULD1 port map( A => n431, B => n420, CI => n418, CO => n415, S => 
                           n416);
   U397 : ADFULD1 port map( A => n443, B => n434, CI => n432, CO => n429, S => 
                           n430);
   U398 : ADFULD1 port map( A => n447, B => n445, CI => n436, CO => n431, S => 
                           n432);
   U405 : ADFULD1 port map( A => n450, B => n621, CI => n636, CO => n445, S => 
                           n446);
   U407 : ADFULD1 port map( A => n561, B => n452, CI => n576, CO => n449, S => 
                           n450);
   U409 : ADFULD1 port map( A => n458, B => n465, CI => n456, CO => n453, S => 
                           n454);
   U410 : ADFULD1 port map( A => n460, B => n637, CI => n467, CO => n455, S => 
                           n456);
   U412 : ADFULD1 port map( A => n592, B => n577, CI => n462, CO => n459, S => 
                           n460);
   U413 : ADFULD1 port map( A => n471, B => n547, CI => n562, CO => n461, S => 
                           n462);
   U414 : ADFULD1 port map( A => n468, B => n475, CI => n466, CO => n463, S => 
                           n464);
   U415 : ADFULD1 port map( A => n470, B => n638, CI => n477, CO => n465, S => 
                           n466);
   U416 : ADFULD1 port map( A => n608, B => n479, CI => n623, CO => n467, S => 
                           n468);
   U421 : ADFULD1 port map( A => n609, B => n594, CI => n480, CO => n477, S => 
                           n478);
   U422 : ADFULD1 port map( A => n487, B => n564, CI => n579, CO => n479, S => 
                           n480);
   U423 : ADFULD1 port map( A => n491, B => n486, CI => n484, CO => n481, S => 
                           n482);
   U424 : ADFULD1 port map( A => n625, B => n493, CI => n640, CO => n483, S => 
                           n484);
   U425 : ADFULD1 port map( A => n595, B => n488, CI => n610, CO => n485, S => 
                           n486);
   U427 : ADFULD1 port map( A => n641, B => n497, CI => n492, CO => n489, S => 
                           n490);
   U428 : ADFULD1 port map( A => n626, B => n611, CI => n494, CO => n491, S => 
                           n492);
   U429 : ADFULD1 port map( A => n499, B => n581, CI => n596, CO => n493, S => 
                           n494);
   U430 : ADFULD1 port map( A => n642, B => n503, CI => n498, CO => n495, S => 
                           n496);
   U431 : ADFULD1 port map( A => n612, B => n500, CI => n627, CO => n497, S => 
                           n498);
   U433 : ADFULD1 port map( A => n643, B => n628, CI => n504, CO => n501, S => 
                           n502);
   U434 : ADFULD1 port map( A => n507, B => n598, CI => n613, CO => n503, S => 
                           n504);
   U435 : ADFULD1 port map( A => n629, B => n508, CI => n644, CO => n505, S => 
                           n506);
   U439 : OAI22D1 port map( A1 => n48, A2 => n920, B1 => n665, B2 => n46, Z => 
                           n513);
   U441 : OAI22D1 port map( A1 => n651, A2 => n48, B1 => n650, B2 => n46, Z => 
                           n522);
   U444 : OAI22D1 port map( A1 => n654, A2 => n48, B1 => n653, B2 => n46, Z => 
                           n319);
   U445 : OAI22D1 port map( A1 => n654, A2 => n46, B1 => n655, B2 => n48, Z => 
                           n525);
   U448 : OAI22D1 port map( A1 => n658, A2 => n48, B1 => n657, B2 => n46, Z => 
                           n351);
   U449 : OAI22D1 port map( A1 => n659, A2 => n48, B1 => n658, B2 => n46, Z => 
                           n527);
   U450 : OAI22D1 port map( A1 => n660, A2 => n48, B1 => n659, B2 => n46, Z => 
                           n373);
   U451 : OAI22D1 port map( A1 => n661, A2 => n48, B1 => n660, B2 => n46, Z => 
                           n528);
   U454 : OAI22D1 port map( A1 => n664, A2 => n48, B1 => n663, B2 => n46, Z => 
                           n530);
   U455 : NOR2M1D1 port map( A1 => b(0), A2 => n46, Z => n531);
   U471 : EXNOR2D1 port map( A1 => b(0), A2 => a(15), Z => n664);
   U472 : NAN2M1D1 port map( A1 => b(0), A2 => a(15), Z => n665);
   U473 : OAI22D1 port map( A1 => n42, A2 => n826, B1 => n682, B2 => n40, Z => 
                           n514);
   U475 : OAI22D1 port map( A1 => n667, A2 => n42, B1 => n666, B2 => n40, Z => 
                           n309);
   U477 : OAI22D1 port map( A1 => n669, A2 => n42, B1 => n668, B2 => n40, Z => 
                           n534);
   U479 : OAI22D1 port map( A1 => n42, A2 => n671, B1 => n670, B2 => n40, Z => 
                           n536);
   U480 : OAI22D1 port map( A1 => n671, A2 => n40, B1 => n672, B2 => n42, Z => 
                           n537);
   U481 : OAI22D1 port map( A1 => n673, A2 => n42, B1 => n672, B2 => n40, Z => 
                           n538);
   U482 : OAI22D1 port map( A1 => n674, A2 => n42, B1 => n673, B2 => n40, Z => 
                           n539);
   U483 : OAI22D1 port map( A1 => n675, A2 => n42, B1 => n674, B2 => n40, Z => 
                           n540);
   U484 : OAI22D1 port map( A1 => n676, A2 => n42, B1 => n675, B2 => n40, Z => 
                           n541);
   U489 : OAI22D1 port map( A1 => n681, A2 => n42, B1 => n680, B2 => n40, Z => 
                           n546);
   U490 : NOR2M1D1 port map( A1 => b(0), A2 => n40, Z => n547);
   U506 : EXNOR2D1 port map( A1 => b(0), A2 => a(13), Z => n681);
   U507 : NAN2M1D1 port map( A1 => b(0), A2 => a(13), Z => n682);
   U508 : OAI22D1 port map( A1 => n36, A2 => n827, B1 => n699, B2 => n34, Z => 
                           n515);
   U511 : OAI22D1 port map( A1 => n685, A2 => n36, B1 => n684, B2 => n34, Z => 
                           n550);
   U512 : OAI22D1 port map( A1 => n686, A2 => n36, B1 => n685, B2 => n34, Z => 
                           n551);
   U513 : OAI22D1 port map( A1 => n687, A2 => n36, B1 => n686, B2 => n34, Z => 
                           n552);
   U515 : OAI22D1 port map( A1 => n688, A2 => n34, B1 => n689, B2 => n36, Z => 
                           n554);
   U516 : OAI22D1 port map( A1 => n690, A2 => n36, B1 => n689, B2 => n34, Z => 
                           n555);
   U517 : OAI22D1 port map( A1 => n691, A2 => n36, B1 => n690, B2 => n34, Z => 
                           n556);
   U521 : OAI22D1 port map( A1 => n695, A2 => n36, B1 => n694, B2 => n34, Z => 
                           n560);
   U522 : OAI22D1 port map( A1 => n696, A2 => n36, B1 => n695, B2 => n34, Z => 
                           n561);
   U524 : OAI22D1 port map( A1 => n698, A2 => n36, B1 => n697, B2 => n34, Z => 
                           n563);
   U525 : NOR2M1D1 port map( A1 => b(0), A2 => n34, Z => n564);
   U537 : EXNOR2D1 port map( A1 => b(4), A2 => a(11), Z => n694);
   U541 : EXNOR2D1 port map( A1 => b(0), A2 => a(11), Z => n698);
   U542 : NAN2M1D1 port map( A1 => b(0), A2 => a(11), Z => n699);
   U543 : OAI22D1 port map( A1 => n30, A2 => n828, B1 => n716, B2 => n28, Z => 
                           n516);
   U546 : OAI22D1 port map( A1 => n702, A2 => n30, B1 => n701, B2 => n28, Z => 
                           n567);
   U547 : OAI22D1 port map( A1 => n703, A2 => n30, B1 => n702, B2 => n28, Z => 
                           n568);
   U548 : OAI22D1 port map( A1 => n704, A2 => n30, B1 => n703, B2 => n28, Z => 
                           n569);
   U549 : OAI22D1 port map( A1 => n30, A2 => n705, B1 => n704, B2 => n28, Z => 
                           n570);
   U550 : OAI22D1 port map( A1 => n705, A2 => n28, B1 => n706, B2 => n30, Z => 
                           n571);
   U553 : OAI22D1 port map( A1 => n709, A2 => n30, B1 => n708, B2 => n28, Z => 
                           n574);
   U554 : OAI22D1 port map( A1 => n710, A2 => n30, B1 => n709, B2 => n28, Z => 
                           n575);
   U555 : OAI22D1 port map( A1 => n711, A2 => n30, B1 => n710, B2 => n28, Z => 
                           n576);
   U556 : OAI22D1 port map( A1 => n712, A2 => n30, B1 => n711, B2 => n28, Z => 
                           n577);
   U559 : OAI22D1 port map( A1 => n715, A2 => n30, B1 => n714, B2 => n28, Z => 
                           n580);
   U560 : NOR2M1D1 port map( A1 => b(0), A2 => n28, Z => n581);
   U572 : EXNOR2D1 port map( A1 => b(4), A2 => a(9), Z => n711);
   U576 : EXNOR2D1 port map( A1 => b(0), A2 => a(9), Z => n715);
   U577 : NAN2M1D1 port map( A1 => b(0), A2 => a(9), Z => n716);
   U578 : OAI22D1 port map( A1 => n24, A2 => n829, B1 => n733, B2 => n22, Z => 
                           n517);
   U581 : OAI22D1 port map( A1 => n719, A2 => n24, B1 => n718, B2 => n22, Z => 
                           n584);
   U582 : OAI22D1 port map( A1 => n720, A2 => n24, B1 => n719, B2 => n22, Z => 
                           n585);
   U583 : OAI22D1 port map( A1 => n721, A2 => n24, B1 => n720, B2 => n22, Z => 
                           n586);
   U584 : OAI22D1 port map( A1 => n722, A2 => n24, B1 => n721, B2 => n22, Z => 
                           n587);
   U585 : OAI22D1 port map( A1 => n722, A2 => n22, B1 => n723, B2 => n24, Z => 
                           n588);
   U587 : OAI22D1 port map( A1 => n725, A2 => n24, B1 => n724, B2 => n22, Z => 
                           n590);
   U589 : OAI22D1 port map( A1 => n727, A2 => n24, B1 => n726, B2 => n22, Z => 
                           n592);
   U591 : OAI22D1 port map( A1 => n729, A2 => n24, B1 => n728, B2 => n22, Z => 
                           n594);
   U594 : OAI22D1 port map( A1 => n732, A2 => n24, B1 => n731, B2 => n22, Z => 
                           n597);
   U595 : NOR2M1D1 port map( A1 => b(0), A2 => n22, Z => n598);
   U607 : EXNOR2D1 port map( A1 => b(4), A2 => a(7), Z => n728);
   U611 : EXNOR2D1 port map( A1 => b(0), A2 => a(7), Z => n732);
   U612 : NAN2M1D1 port map( A1 => b(0), A2 => a(7), Z => n733);
   U613 : OAI22D1 port map( A1 => n18, A2 => n830, B1 => n750, B2 => n16, Z => 
                           n518);
   U616 : OAI22D1 port map( A1 => n736, A2 => n18, B1 => n735, B2 => n16, Z => 
                           n601);
   U617 : OAI22D1 port map( A1 => n737, A2 => n18, B1 => n736, B2 => n16, Z => 
                           n602);
   U620 : OAI22D1 port map( A1 => n739, A2 => n16, B1 => n740, B2 => n18, Z => 
                           n605);
   U623 : OAI22D1 port map( A1 => n743, A2 => n18, B1 => n742, B2 => n16, Z => 
                           n608);
   U624 : OAI22D1 port map( A1 => n744, A2 => n18, B1 => n743, B2 => n16, Z => 
                           n609);
   U625 : OAI22D1 port map( A1 => n745, A2 => n18, B1 => n744, B2 => n16, Z => 
                           n610);
   U626 : OAI22D1 port map( A1 => n746, A2 => n18, B1 => n745, B2 => n16, Z => 
                           n611);
   U629 : OAI22D1 port map( A1 => n749, A2 => n18, B1 => n748, B2 => n16, Z => 
                           n614);
   U630 : NOR2M1D1 port map( A1 => b(0), A2 => n16, Z => n615);
   U642 : EXNOR2D1 port map( A1 => b(4), A2 => a(5), Z => n745);
   U646 : EXNOR2D1 port map( A1 => b(0), A2 => a(5), Z => n749);
   U647 : NAN2M1D1 port map( A1 => b(0), A2 => a(5), Z => n750);
   U648 : OAI22D1 port map( A1 => n12, A2 => n831, B1 => n767, B2 => n9, Z => 
                           n519);
   U649 : AO21D2 port map( A1 => n12, A2 => n9, B => n751, Z => n616);
   U651 : OAI22D1 port map( A1 => n753, A2 => n12, B1 => n752, B2 => n9, Z => 
                           n618);
   U653 : OAI22D1 port map( A1 => n755, A2 => n12, B1 => n754, B2 => n9, Z => 
                           n620);
   U654 : OAI22D1 port map( A1 => n756, A2 => n12, B1 => n755, B2 => n9, Z => 
                           n621);
   U655 : OAI22D1 port map( A1 => n756, A2 => n9, B1 => n757, B2 => n12, Z => 
                           n622);
   U656 : OAI22D1 port map( A1 => n758, A2 => n12, B1 => n757, B2 => n9, Z => 
                           n623);
   U657 : OAI22D1 port map( A1 => n759, A2 => n12, B1 => n758, B2 => n9, Z => 
                           n624);
   U658 : OAI22D1 port map( A1 => n760, A2 => n12, B1 => n759, B2 => n9, Z => 
                           n625);
   U659 : OAI22D1 port map( A1 => n761, A2 => n12, B1 => n760, B2 => n9, Z => 
                           n626);
   U660 : OAI22D1 port map( A1 => n762, A2 => n12, B1 => n761, B2 => n9, Z => 
                           n627);
   U661 : OAI22D1 port map( A1 => n763, A2 => n12, B1 => n762, B2 => n9, Z => 
                           n628);
   U664 : OAI22D1 port map( A1 => n766, A2 => n12, B1 => n765, B2 => n9, Z => 
                           n631);
   U665 : NOR2M1D1 port map( A1 => b(0), A2 => n9, Z => n632);
   U681 : EXNOR2D1 port map( A1 => b(0), A2 => a(3), Z => n766);
   U682 : NAN2M1D1 port map( A1 => b(0), A2 => a(3), Z => n767);
   U683 : OAI22D1 port map( A1 => n6, A2 => n832, B1 => n784, B2 => n824, Z => 
                           n520);
   U686 : OAI22D1 port map( A1 => n770, A2 => n6, B1 => n769, B2 => n824, Z => 
                           n635);
   U687 : OAI22D1 port map( A1 => n771, A2 => n6, B1 => n770, B2 => n824, Z => 
                           n636);
   U688 : OAI22D1 port map( A1 => n772, A2 => n6, B1 => n771, B2 => n824, Z => 
                           n637);
   U689 : OAI22D1 port map( A1 => n773, A2 => n6, B1 => n772, B2 => n824, Z => 
                           n638);
   U691 : OAI22D1 port map( A1 => n775, A2 => n6, B1 => n774, B2 => n824, Z => 
                           n640);
   U692 : OAI22D1 port map( A1 => n776, A2 => n6, B1 => n775, B2 => n824, Z => 
                           n641);
   U693 : OAI22D1 port map( A1 => n777, A2 => n6, B1 => n776, B2 => n824, Z => 
                           n642);
   U694 : OAI22D1 port map( A1 => n778, A2 => n6, B1 => n777, B2 => n824, Z => 
                           n643);
   U695 : OAI22D1 port map( A1 => n779, A2 => n6, B1 => n778, B2 => n824, Z => 
                           n644);
   U696 : OAI22D1 port map( A1 => n780, A2 => n6, B1 => n779, B2 => n824, Z => 
                           n645);
   U698 : OAI22D1 port map( A1 => n782, A2 => n6, B1 => n781, B2 => n824, Z => 
                           n647);
   U699 : OAI22D1 port map( A1 => n783, A2 => n6, B1 => n782, B2 => n824, Z => 
                           n648);
   U716 : EXNOR2D1 port map( A1 => b(0), A2 => a(1), Z => n783);
   U717 : NAN2M1D1 port map( A1 => b(0), A2 => a(1), Z => n784);
   U742 : EXOR2D1 port map( A1 => a(15), A2 => a(14), Z => n801);
   U754 : EXOR2D1 port map( A1 => a(7), A2 => a(6), Z => n805);
   U757 : EXOR2D1 port map( A1 => a(5), A2 => a(4), Z => n806);
   U760 : EXOR2D1 port map( A1 => a(3), A2 => a(2), Z => n807);
   U763 : EXOR2D1 port map( A1 => a(1), A2 => a(0), Z => n808);
   U751 : EXOR2D1 port map( A1 => a(9), A2 => a(8), Z => n804);
   U217 : AOI21D1 port map( A1 => n204, A2 => n212, B => n205, Z => n203);
   U485 : OAI22D1 port map( A1 => n677, A2 => n42, B1 => n676, B2 => n40, Z => 
                           n542);
   U502 : EXNOR2D1 port map( A1 => b(4), A2 => a(13), Z => n677);
   U745 : EXOR2D1 port map( A1 => a(13), A2 => a(12), Z => n802);
   U487 : OAI22D1 port map( A1 => n679, A2 => n42, B1 => n678, B2 => n40, Z => 
                           n544);
   U748 : EXOR2D1 port map( A1 => a(11), A2 => a(10), Z => n803);
   U520 : OAI22D1 port map( A1 => n694, A2 => n36, B1 => n693, B2 => n34, Z => 
                           n559);
   U518 : OAI22D1 port map( A1 => n692, A2 => n36, B1 => n691, B2 => n34, Z => 
                           n557);
   U486 : OAI22D1 port map( A1 => n678, A2 => n42, B1 => n677, B2 => n40, Z => 
                           n543);
   U519 : OAI22D1 port map( A1 => n693, A2 => n36, B1 => n692, B2 => n34, Z => 
                           n558);
   U387 : ADFULD1 port map( A => n414, B => n543, CI => n558, CO => n411, S => 
                           n412);
   U379 : ADFULD1 port map( A => n572, B => n557, CI => n411, CO => n395, S => 
                           n396);
   U370 : ADFULD1 port map( A => n382, B => n384, CI => n391, CO => n377, S => 
                           n378);
   U402 : ADFULD1 port map( A => n451, B => n531, CI => n545, CO => n439, S => 
                           n440);
   U586 : OAI22D1 port map( A1 => n24, A2 => n724, B1 => n723, B2 => n22, Z => 
                           n589);
   U391 : ADFULD1 port map( A => n433, B => n424, CI => n422, CO => n417, S => 
                           n418);
   U384 : ADFULD1 port map( A => n423, B => n633, CI => n421, CO => n405, S => 
                           n406);
   U183 : NOR2D2 port map( A1 => n364, A2 => n375, Z => n179);
   U193 : NOR2D2 port map( A1 => n376, A2 => n387, Z => n184);
   U162 : OAI21D1 port map( A1 => n167, A2 => n173, B => n168, Z => n162);
   U132 : OAI21D1 port map( A1 => n164, A2 => n143, B => n144, Z => n142);
   U144 : AOI21D1 port map( A1 => net11621, A2 => n152, B => n153, Z => n151);
   U178 : AOI21D1 port map( A1 => n177, A2 => net12065, B => n178, Z => n176);
   U551 : OAI22D1 port map( A1 => n707, A2 => n30, B1 => n706, B2 => n28, Z => 
                           n572);
   U767 : EXOR2D1 port map( A1 => net11503, A2 => n404, Z => n402);
   U768 : OAI22D1 port map( A1 => n680, A2 => n42, B1 => n679, B2 => n40, Z => 
                           n545);
   U769 : EXNOR2D2 port map( A1 => b(1), A2 => a(13), Z => n680);
   U770 : OAI22DL port map( A1 => n714, A2 => n30, B1 => n713, B2 => n28, Z => 
                           n579);
   U771 : OAI22DL port map( A1 => n713, A2 => n30, B1 => n712, B2 => n28, Z => 
                           n578);
   U772 : OAI22DL port map( A1 => n663, A2 => n48, B1 => n662, B2 => n46, Z => 
                           n529);
   U773 : OAI22DL port map( A1 => n765, A2 => n12, B1 => n764, B2 => n9, Z => 
                           n630);
   U774 : OAI22DL port map( A1 => n764, A2 => n12, B1 => n763, B2 => n9, Z => 
                           n629);
   U775 : OAI22DL port map( A1 => n731, A2 => n24, B1 => n730, B2 => n22, Z => 
                           n596);
   U776 : OAI22DL port map( A1 => n730, A2 => n24, B1 => n729, B2 => n22, Z => 
                           n595);
   U777 : OAI22DL port map( A1 => n748, A2 => n18, B1 => n747, B2 => n16, Z => 
                           n613);
   U778 : OAI22DL port map( A1 => n747, A2 => n18, B1 => n746, B2 => n16, Z => 
                           n612);
   U779 : OAI22DL port map( A1 => n781, A2 => n6, B1 => n780, B2 => n824, Z => 
                           n646);
   U780 : EXNOR2D1 port map( A1 => n529, A2 => n427, Z => n414);
   U781 : OR2D1 port map( A1 => n529, A2 => n427, Z => n413);
   U782 : ADFULDL port map( A => n511, B => n615, CI => n630, CO => n509, S => 
                           n510);
   U783 : OR2DL port map( A1 => n647, A2 => n632, Z => n1006);
   U784 : EXNOR2D1 port map( A1 => b(10), A2 => a(13), Z => n671);
   U785 : AOI21M10D1 port map( A1 => n163, A2 => net11621, B => n904, Z => n160
                           );
   U786 : EXOR2D2 port map( A1 => n973, A2 => n379, Z => n366);
   U787 : INVDL port map( A => n284, Z => n900);
   U788 : OAI21DL port map( A1 => n195, A2 => n201, B => n196, Z => n901);
   U789 : EXOR3D1 port map( A1 => n382, A2 => n384, A3 => n391, Z => n902);
   U790 : EXNOR2D2 port map( A1 => b(6), A2 => a(7), Z => n726);
   U791 : EXNOR2D2 port map( A1 => b(9), A2 => a(9), Z => n706);
   U792 : OAI21DL port map( A1 => n134, A2 => n155, B => n135, Z => n903);
   U793 : OA21M20DL port map( A1 => net11083, A2 => n148, B => n139, Z => n135)
                           ;
   U794 : BUFDL port map( A => n162, Z => n904);
   U795 : OAI21DL port map( A1 => n164, A2 => n154, B => n155, Z => n153);
   U796 : EXNOR2D2 port map( A1 => b(9), A2 => a(15), Z => n655);
   U797 : INVDL port map( A => n203, Z => n202);
   U798 : EXNOR2D2 port map( A1 => b(7), A2 => a(13), Z => n674);
   U799 : NAN3D2 port map( A1 => n907, A2 => n909, A3 => n908, Z => n391);
   U800 : EXNOR2D2 port map( A1 => b(1), A2 => a(11), Z => n697);
   U801 : EXNOR2D2 port map( A1 => b(8), A2 => a(7), Z => n724);
   U802 : OAI22D1 port map( A1 => n16, A2 => n734, B1 => n18, B2 => n735, Z => 
                           n600);
   U803 : OAI22D1 port map( A1 => n726, A2 => n24, B1 => n725, B2 => n22, Z => 
                           n591);
   U804 : EXNOR2D1 port map( A1 => b(15), A2 => a(5), Z => n734);
   U805 : EXNOR2D2 port map( A1 => b(7), A2 => a(9), Z => n708);
   U806 : EXNOR2DL port map( A1 => b(4), A2 => a(15), Z => n660);
   U807 : EXNOR2DL port map( A1 => b(4), A2 => a(1), Z => n779);
   U808 : EXNOR2DL port map( A1 => b(4), A2 => a(3), Z => n762);
   U809 : OAI22D1 port map( A1 => n739, A2 => n18, B1 => n738, B2 => n16, Z => 
                           n905);
   U810 : OAI22DL port map( A1 => n739, A2 => n18, B1 => n738, B2 => n16, Z => 
                           n604);
   U811 : EXNOR2D2 port map( A1 => b(11), A2 => a(5), Z => n738);
   U812 : NAN2D2 port map( A1 => n354, A2 => n363, Z => n173);
   U813 : EXNOR2D1 port map( A1 => b(12), A2 => a(5), Z => n737);
   U814 : INVD4 port map( A => n399, Z => n400);
   U815 : OAI22D4 port map( A1 => n662, A2 => n48, B1 => n661, B2 => n46, Z => 
                           n399);
   U816 : EXOR2D1 port map( A1 => n617, A2 => n409, Z => n906);
   U817 : EXOR2D1 port map( A1 => n906, A2 => n396, Z => n392);
   U818 : NAN2D1 port map( A1 => n396, A2 => n409, Z => n907);
   U819 : NAN2D1 port map( A1 => n396, A2 => n617, Z => n908);
   U820 : NAN2DL port map( A1 => n409, A2 => n617, Z => n909);
   U821 : OAI22D2 port map( A1 => n752, A2 => n12, B1 => n751, B2 => n9, Z => 
                           n617);
   U822 : OAI22DL port map( A1 => n688, A2 => n36, B1 => n687, B2 => n34, Z => 
                           n553);
   U823 : OAI22DL port map( A1 => n741, A2 => n18, B1 => n740, B2 => n16, Z => 
                           n606);
   U824 : EXOR2D1 port map( A1 => n934, A2 => n559, Z => n426);
   U825 : INVD1 port map( A => n56, Z => n947);
   U826 : INVD1 port map( A => n377, Z => n915);
   U827 : INVD1 port map( A => a(15), Z => n920);
   U828 : EXNOR2D2 port map( A1 => n197, A2 => n910, Z => product(17));
   U829 : AND2DL port map( A1 => n287, A2 => n196, Z => n910);
   U830 : EXNOR2D1 port map( A1 => b(11), A2 => a(7), Z => n721);
   U831 : OR2DL port map( A1 => n482, A2 => n489, Z => n998);
   U832 : AOI21D1 port map( A1 => n991, A2 => n999, B => n911, Z => n232);
   U833 : AND2DL port map( A1 => n474, A2 => n481, Z => n911);
   U834 : EXOR2D2 port map( A1 => n455, A2 => n446, Z => n958);
   U835 : EXOR3DL port map( A1 => n424, A2 => n433, A3 => n422, Z => n912);
   U836 : NAN2M1D1 port map( A1 => n206, A2 => n207, Z => n68);
   U837 : OR2D2 port map( A1 => n474, A2 => n481, Z => n991);
   U838 : EXNOR2D2 port map( A1 => b(10), A2 => a(3), Z => n756);
   U839 : EXNOR2DL port map( A1 => b(3), A2 => a(1), Z => n780);
   U840 : AOI22M10D1 port map( B1 => n995, B2 => n230, A1 => n923, A2 => n464, 
                           Z => n225);
   U841 : NOR2DL port map( A1 => n364, A2 => n375, Z => n913);
   U842 : NAN3D1 port map( A1 => net11666, A2 => net11667, A3 => n972, Z => 
                           n379);
   U843 : NAN2D1 port map( A1 => n605, A2 => n449, Z => n984);
   U844 : EXOR3D2 port map( A1 => n979, A2 => n905, A3 => n426, Z => n422);
   U845 : EXNOR2DL port map( A1 => b(2), A2 => a(1), Z => n781);
   U846 : OAI22D1 port map( A1 => n769, A2 => n6, B1 => n768, B2 => n824, Z => 
                           n634);
   U847 : BUFDL port map( A => b(11), Z => n914);
   U848 : EXNOR2DL port map( A1 => b(6), A2 => a(3), Z => n760);
   U849 : EXNOR2D2 port map( A1 => n208, A2 => n68, Z => product(15));
   U850 : EXNOR2D2 port map( A1 => n169, A2 => n989, Z => product(21));
   U851 : EXNOR2DL port map( A1 => b(2), A2 => a(5), Z => n747);
   U852 : ADFULD2 port map( A => n380, B => n389, CI => n378, CO => n375, S => 
                           n_1033);
   U853 : ADFULD2 port map( A => n574, B => n439, CI => n589, CO => n423, S => 
                           n424);
   U854 : NAN2DL port map( A1 => n377, A2 => n368, Z => n917);
   U855 : NAN2D1 port map( A1 => n915, A2 => n916, Z => n918);
   U856 : NAN2D1 port map( A1 => n917, A2 => n918, Z => net11025);
   U857 : INVDL port map( A => n368, Z => n916);
   U858 : NAN2D1 port map( A1 => b(1), A2 => a(15), Z => n921);
   U859 : NAN2D2 port map( A1 => n919, A2 => n920, Z => n922);
   U860 : NAN2D2 port map( A1 => n921, A2 => n922, Z => n663);
   U861 : INVD2 port map( A => b(1), Z => n919);
   U862 : INVBD2 port map( A => net10037, Z => net11621);
   U863 : AOI21DL port map( A1 => n288, A2 => n202, B => n199, Z => n197);
   U864 : NAN2D1 port map( A1 => n990, A2 => n993, Z => n213);
   U865 : ADHALFD1 port map( A => n580, B => n516, CO => n487, S => n488);
   U866 : EXNOR2D2 port map( A1 => b(1), A2 => a(9), Z => n714);
   U867 : NAN2M1D1 port map( A1 => n209, A2 => n931, Z => n69);
   U868 : NAN2D1 port map( A1 => n605, A2 => n590, Z => n985);
   U869 : AOI21M20DL port map( A1 => n336, A2 => n343, B => n163, Z => n152);
   U870 : INVDL port map( A => n473, Z => n923);
   U871 : OA21M20D1 port map( A1 => n283, A2 => n924, B => n168, Z => n164);
   U872 : INVDL port map( A => n173, Z => n924);
   U873 : EXOR3D1 port map( A1 => n389, A2 => n380, A3 => n902, Z => n376);
   U874 : EXNOR2D2 port map( A1 => b(5), A2 => a(11), Z => n693);
   U875 : NAN2D1 port map( A1 => n177, A2 => n189, Z => n175);
   U876 : OAI21D1 port map( A1 => n175, A2 => n203, B => n176, Z => n51);
   U877 : NOR2D2 port map( A1 => n184, A2 => n179, Z => n177);
   U878 : NOR2D1 port map( A1 => n195, A2 => n200, Z => n189);
   U879 : BUFDL port map( A => n189, Z => net12127);
   U880 : NOR2M1DL port map( A1 => n189, A2 => net12055, Z => n182);
   U881 : INVDL port map( A => n184, Z => net12054);
   U882 : OAI21D1 port map( A1 => n187, A2 => n179, B => n180, Z => n178);
   U883 : INVDL port map( A => n195, Z => n287);
   U884 : OAI21D1 port map( A1 => n195, A2 => n201, B => n196, Z => net12065);
   U885 : INVDL port map( A => n200, Z => n288);
   U886 : EXNOR2D2 port map( A1 => n151, A2 => net11675, Z => product(23));
   U887 : AND2DL port map( A1 => net11096, A2 => n150, Z => net11675);
   U888 : INVDL port map( A => n161, Z => n163);
   U889 : NOR2DL port map( A1 => n163, A2 => n143, Z => n141);
   U890 : EXNOR2DL port map( A1 => net11621, A2 => n63, Z => product(20));
   U891 : INVD2 port map( A => n51, Z => net10037);
   U892 : INVBD2 port map( A => net10037, Z => net12285);
   U893 : OR2D1 port map( A1 => n328, A2 => n335, Z => net11096);
   U894 : NAN2DL port map( A1 => n282, A2 => net11096, Z => n143);
   U895 : NAN2D1 port map( A1 => net11096, A2 => net11083, Z => n134);
   U896 : AOI21M10DL port map( A1 => n155, A2 => net11096, B => n148, Z => n144
                           );
   U897 : NAN2DL port map( A1 => n328, A2 => n335, Z => n150);
   U898 : INVD1 port map( A => n150, Z => n148);
   U899 : NOR2D1 port map( A1 => n336, A2 => n343, Z => n154);
   U900 : INVD1 port map( A => n154, Z => n282);
   U901 : NOR2D1 port map( A1 => n134, A2 => n154, Z => n132);
   U902 : NAN2D1 port map( A1 => n336, A2 => n343, Z => n155);
   U903 : AND2DL port map( A1 => n282, A2 => n155, Z => net11662);
   U904 : AOI21DL port map( A1 => n132, A2 => n162, B => n903, Z => net12183);
   U905 : AOI21DL port map( A1 => n132, A2 => n162, B => n903, Z => n52);
   U906 : NOR2D1 port map( A1 => n172, A2 => n167, Z => n161);
   U907 : NAN2D1 port map( A1 => n375, A2 => n364, Z => n180);
   U908 : NAN2D1 port map( A1 => net12019, A2 => n387, Z => n187);
   U909 : EXOR3DL port map( A1 => n389, A2 => n380, A3 => n902, Z => net12019);
   U910 : ADFULD2 port map( A => n394, B => n407, CI => n405, CO => n389, S => 
                           n390);
   U911 : INVDL port map( A => n390, Z => net12152);
   U912 : NAN2D1 port map( A1 => net11693, A2 => n390, Z => net12153);
   U913 : NAN2DL port map( A1 => n390, A2 => n403, Z => net11585);
   U914 : NAN2D1 port map( A1 => n390, A2 => n392, Z => net11586);
   U915 : NAN2DL port map( A1 => n406, A2 => n404, Z => net11509);
   U916 : NAN2DL port map( A1 => n417, A2 => n406, Z => net11507);
   U917 : EXOR2D2 port map( A1 => n417, A2 => n406, Z => net11503);
   U918 : NAN3D2 port map( A1 => n925, A2 => n927, A3 => n926, Z => n421);
   U919 : NAN2D1 port map( A1 => n634, A2 => n905, Z => n926);
   U920 : INVD1 port map( A => a(0), Z => n824);
   U921 : NAN2D1 port map( A1 => n634, A2 => n426, Z => n927);
   U922 : NAN2DL port map( A1 => n604, A2 => n426, Z => n925);
   U923 : AO21D2 port map( A1 => n6, A2 => n824, B => n768, Z => n633);
   U924 : NAN2DL port map( A1 => n560, A2 => n440, Z => net12079);
   U925 : NAN2DL port map( A1 => n575, A2 => n440, Z => net12078);
   U926 : EXOR3D2 port map( A1 => n575, A2 => n560, A3 => n440, Z => n438);
   U927 : EXNOR2D1 port map( A1 => n392, A2 => n403, Z => net11693);
   U928 : NAN2DL port map( A1 => n403, A2 => n392, Z => net11587);
   U929 : EXOR3D1 port map( A1 => n395, A2 => n616, A3 => n393, Z => n380);
   U930 : NAN2DL port map( A1 => n395, A2 => n393, Z => net11667);
   U931 : NAN2D1 port map( A1 => n395, A2 => n616, Z => net11666);
   U932 : NAN2DL port map( A1 => n603, A2 => n412, Z => net12126);
   U933 : NAN2DL port map( A1 => n618, A2 => n412, Z => net12125);
   U934 : EXOR3D2 port map( A1 => n412, A2 => n618, A3 => n603, Z => n408);
   U935 : EXNOR2D1 port map( A1 => b(8), A2 => a(9), Z => n707);
   U936 : NAN3D1 port map( A1 => n928, A2 => n930, A3 => n929, Z => n409);
   U937 : NAN2DL port map( A1 => n588, A2 => n573, Z => n929);
   U938 : NAN2DL port map( A1 => n425, A2 => n573, Z => n930);
   U939 : NAN2DL port map( A1 => n588, A2 => n425, Z => n928);
   U940 : NAN2D1 port map( A1 => n803, A2 => n34, Z => n36);
   U941 : EXNOR2D2 port map( A1 => b(6), A2 => a(11), Z => n692);
   U942 : EXNOR2D1 port map( A1 => a(9), A2 => a(10), Z => n34);
   U943 : EXNOR2D2 port map( A1 => b(3), A2 => a(13), Z => n678);
   U944 : NAN2D1 port map( A1 => n802, A2 => n40, Z => n42);
   U945 : EXNOR2D1 port map( A1 => a(11), A2 => a(12), Z => n40);
   U946 : NAN3D1 port map( A1 => net11585, A2 => net11587, A3 => net11586, Z =>
                           n387);
   U947 : NAN2D1 port map( A1 => n161, A2 => n132, Z => n53);
   U948 : AOI21M10DL port map( A1 => n900, A2 => n51, B => n171, Z => n169);
   U949 : EXOR2D1 port map( A1 => net11829, A2 => n571, Z => n384);
   U950 : OAI21D1 port map( A1 => n206, A2 => n210, B => n207, Z => n205);
   U951 : NOR2D1 port map( A1 => n206, A2 => n209, Z => n204);
   U952 : INVDL port map( A => n901, Z => n192);
   U953 : INVDL port map( A => n187, Z => net11745);
   U954 : AND2D1 port map( A1 => n285, A2 => n180, Z => net11172);
   U955 : INVD1 port map( A => n212, Z => n211);
   U956 : BUFDL port map( A => n210, Z => n931);
   U957 : OAI21D1 port map( A1 => n211, A2 => n209, B => n931, Z => n208);
   U958 : NAN2D1 port map( A1 => n804, A2 => n28, Z => n30);
   U959 : EXNOR2D1 port map( A1 => a(7), A2 => a(8), Z => n28);
   U960 : EXNOR2D2 port map( A1 => b(11), A2 => a(9), Z => n704);
   U961 : EXNOR2D2 port map( A1 => net12250, A2 => a(13), Z => n672);
   U962 : EXNOR2DL port map( A1 => b(6), A2 => a(1), Z => n777);
   U963 : INVDL port map( A => n915, Z => net12257);
   U964 : OAI22D1 port map( A1 => n656, A2 => n48, B1 => n655, B2 => n46, Z => 
                           n333);
   U965 : EXOR3D1 port map( A1 => n590, A2 => n449, A3 => n605, Z => n436);
   U966 : NAN2DL port map( A1 => n606, A2 => n461, Z => n967);
   U967 : INVDL port map( A => b(9), Z => net12249);
   U968 : INVDL port map( A => net12249, Z => net12250);
   U969 : EXNOR2DL port map( A1 => b(6), A2 => a(15), Z => n658);
   U970 : EXNOR2D2 port map( A1 => b(10), A2 => a(7), Z => n722);
   U971 : OAI22DL port map( A1 => n728, A2 => n24, B1 => n727, B2 => n22, Z => 
                           n593);
   U972 : EXNOR2DL port map( A1 => b(2), A2 => a(7), Z => n730);
   U973 : NAN2D1 port map( A1 => net12151, A2 => net12152, Z => n932);
   U974 : NAN2D2 port map( A1 => net12153, A2 => n932, Z => n388);
   U975 : INVD1 port map( A => net11693, Z => net12151);
   U976 : NAN2DL port map( A1 => n618, A2 => n603, Z => n933);
   U977 : NAN3D1 port map( A1 => n933, A2 => net12126, A3 => net12125, Z => 
                           n407);
   U978 : OAI22DL port map( A1 => n738, A2 => n18, B1 => n737, B2 => n16, Z => 
                           n603);
   U979 : EXOR2D1 port map( A1 => n544, A2 => n428, Z => n934);
   U980 : NAN2DL port map( A1 => n559, A2 => n544, Z => n935);
   U981 : NAN2DL port map( A1 => n559, A2 => n428, Z => n936);
   U982 : NAN2DL port map( A1 => n544, A2 => n428, Z => n937);
   U983 : NAN3D1 port map( A1 => n935, A2 => n937, A3 => n936, Z => n425);
   U984 : ADHALFD2 port map( A => n513, B => n530, CO => n427, S => n428);
   U985 : OAI22D1 port map( A1 => n742, A2 => n18, B1 => n741, B2 => n16, Z => 
                           n607);
   U986 : EXNOR2D1 port map( A1 => a(3), A2 => b(9), Z => n757);
   U987 : EXNOR2D2 port map( A1 => b(7), A2 => a(11), Z => n691);
   U988 : EXNOR2D2 port map( A1 => b(7), A2 => a(7), Z => n725);
   U989 : INVDL port map( A => n171, Z => net12095);
   U990 : EXOR2D1 port map( A1 => n620, A2 => n635, Z => n938);
   U991 : EXOR2D1 port map( A1 => n938, A2 => n438, Z => n434);
   U992 : NAN2DL port map( A1 => n575, A2 => n560, Z => n939);
   U993 : NAN3D1 port map( A1 => n939, A2 => net12078, A3 => net12079, Z => 
                           n437);
   U994 : NAN2D1 port map( A1 => n620, A2 => n635, Z => n940);
   U995 : NAN2D1 port map( A1 => n620, A2 => n438, Z => n941);
   U996 : NAN2D1 port map( A1 => n635, A2 => n438, Z => n942);
   U997 : NAN3D2 port map( A1 => n940, A2 => n941, A3 => n942, Z => n433);
   U998 : EXOR3DL port map( A1 => n431, A2 => n420, A3 => n912, Z => n943);
   U999 : EXNOR2D2 port map( A1 => b(13), A2 => a(3), Z => n753);
   U1000 : INVDL port map( A => n373, Z => n374);
   U1001 : INVD1 port map( A => net12054, Z => net12055);
   U1002 : EXNOR2DL port map( A1 => b(8), A2 => a(11), Z => n690);
   U1003 : INVD2 port map( A => n351, Z => n352);
   U1004 : OAI22D2 port map( A1 => n657, A2 => n48, B1 => n656, B2 => n46, Z =>
                           n526);
   U1005 : INVDL port map( A => n192, Z => net12033);
   U1006 : AOI21DL port map( A1 => net12285, A2 => n106, B => n107, Z => n105);
   U1007 : EXNOR2DL port map( A1 => b(8), A2 => a(15), Z => n656);
   U1008 : EXNOR2DL port map( A1 => b(8), A2 => a(5), Z => n741);
   U1009 : EXNOR2D2 port map( A1 => b(11), A2 => a(3), Z => n755);
   U1010 : OAI22DL port map( A1 => n697, A2 => n36, B1 => n696, B2 => n34, Z =>
                           n562);
   U1011 : ADHALFD2 port map( A => n563, B => n515, CO => n471, S => n472);
   U1012 : EXNOR2DL port map( A1 => b(2), A2 => a(3), Z => n764);
   U1013 : EXNOR2D2 port map( A1 => b(13), A2 => a(1), Z => n770);
   U1014 : OAI21DL port map( A1 => n192, A2 => net12055, B => net11746, Z => 
                           n183);
   U1015 : EXNOR2D2 port map( A1 => b(3), A2 => a(15), Z => n661);
   U1016 : EXNOR2DL port map( A1 => b(3), A2 => a(3), Z => n763);
   U1017 : EXNOR2D2 port map( A1 => b(3), A2 => a(5), Z => n746);
   U1018 : EXNOR2D2 port map( A1 => b(3), A2 => a(7), Z => n729);
   U1019 : EXNOR2D2 port map( A1 => b(3), A2 => a(9), Z => n712);
   U1020 : EXNOR2D2 port map( A1 => b(3), A2 => a(11), Z => n695);
   U1021 : EXOR2D1 port map( A1 => n556, A2 => n397, Z => net11829);
   U1022 : NAN2D1 port map( A1 => n571, A2 => n397, Z => n944);
   U1023 : NAN2DL port map( A1 => n571, A2 => n556, Z => n945);
   U1024 : NAN2DL port map( A1 => n397, A2 => n556, Z => n946);
   U1025 : NAN3D1 port map( A1 => n944, A2 => n946, A3 => n945, Z => n383);
   U1026 : EXNOR2D2 port map( A1 => n105, A2 => n947, Z => product(27));
   U1027 : EXNOR2D2 port map( A1 => b(12), A2 => a(1), Z => n771);
   U1028 : INVD1 port map( A => net11745, Z => net11746);
   U1029 : EXNOR2D2 port map( A1 => n140, A2 => n948, Z => product(24));
   U1030 : AND2DL port map( A1 => net11083, A2 => n139, Z => n948);
   U1031 : NAN2D1 port map( A1 => n943, A2 => n429, Z => n207);
   U1032 : EXNOR2D2 port map( A1 => b(6), A2 => a(9), Z => n709);
   U1033 : EXNOR2D2 port map( A1 => n127, A2 => n949, Z => product(25));
   U1034 : AND2DL port map( A1 => n279, A2 => n118, Z => n949);
   U1035 : EXOR2D1 port map( A1 => n483, A2 => n478, Z => n950);
   U1036 : EXOR2D1 port map( A1 => n950, A2 => n476, Z => n474);
   U1037 : NAN2DL port map( A1 => n476, A2 => n478, Z => n951);
   U1038 : NAN2DL port map( A1 => n476, A2 => n483, Z => n952);
   U1039 : NAN2DL port map( A1 => n478, A2 => n483, Z => n953);
   U1040 : NAN3D1 port map( A1 => n951, A2 => n953, A3 => n952, Z => n473);
   U1041 : EXOR2D1 port map( A1 => n624, A2 => n485, Z => n954);
   U1042 : EXOR2D1 port map( A1 => n954, A2 => n639, Z => n476);
   U1043 : NAN2DL port map( A1 => n639, A2 => n485, Z => n955);
   U1044 : NAN2DL port map( A1 => n639, A2 => n624, Z => n956);
   U1045 : NAN2DL port map( A1 => n485, A2 => n624, Z => n957);
   U1046 : NAN3D1 port map( A1 => n955, A2 => n957, A3 => n956, Z => n475);
   U1047 : OAI22DL port map( A1 => n773, A2 => n824, B1 => n774, B2 => n6, Z =>
                           n639);
   U1048 : EXOR3D1 port map( A1 => n457, A2 => n459, A3 => n448, Z => n444);
   U1049 : EXOR2D1 port map( A1 => n958, A2 => n444, Z => n442);
   U1050 : NAN2DL port map( A1 => n457, A2 => n459, Z => n959);
   U1051 : NAN2DL port map( A1 => n457, A2 => n448, Z => n960);
   U1052 : NAN2D1 port map( A1 => n459, A2 => n448, Z => n961);
   U1053 : NAN3D2 port map( A1 => n959, A2 => n960, A3 => n961, Z => n443);
   U1054 : NAN2DL port map( A1 => n446, A2 => n455, Z => n962);
   U1055 : NAN2DL port map( A1 => n444, A2 => n455, Z => n963);
   U1056 : NAN2DL port map( A1 => n446, A2 => n444, Z => n964);
   U1057 : NAN3D1 port map( A1 => n962, A2 => n963, A3 => n964, Z => n441);
   U1058 : EXOR2D1 port map( A1 => n461, A2 => n591, Z => n965);
   U1059 : EXOR2D1 port map( A1 => n965, A2 => n606, Z => n448);
   U1060 : NAN2DL port map( A1 => n606, A2 => n591, Z => n966);
   U1061 : NAN2DL port map( A1 => n591, A2 => n461, Z => n968);
   U1062 : NAN3D1 port map( A1 => n966, A2 => n968, A3 => n967, Z => n447);
   U1063 : EXOR3D2 port map( A1 => n622, A2 => n469, A3 => n607, Z => n458);
   U1064 : NAN2D1 port map( A1 => n469, A2 => n607, Z => n969);
   U1065 : NAN2D1 port map( A1 => n469, A2 => n622, Z => n970);
   U1066 : NAN2D1 port map( A1 => n607, A2 => n622, Z => n971);
   U1067 : NAN3D2 port map( A1 => n969, A2 => n971, A3 => n970, Z => n457);
   U1068 : ADFULD1 port map( A => n578, B => n472, CI => n593, CO => n469, S =>
                           n470);
   U1069 : NAN2D1 port map( A1 => n430, A2 => n441, Z => n210);
   U1070 : INVD1 port map( A => n167, Z => n283);
   U1071 : OAI22D1 port map( A1 => n769, A2 => n6, B1 => n768, B2 => n824, Z =>
                           n979);
   U1072 : NAN2DL port map( A1 => n616, A2 => n393, Z => n972);
   U1073 : EXOR2D1 port map( A1 => n370, A2 => n381, Z => n973);
   U1074 : NAN2DL port map( A1 => n370, A2 => n381, Z => n974);
   U1075 : NAN2DL port map( A1 => n370, A2 => n379, Z => n975);
   U1076 : NAN2DL port map( A1 => n381, A2 => n379, Z => n976);
   U1077 : NAN3D2 port map( A1 => n974, A2 => n975, A3 => n976, Z => n365);
   U1078 : EXNOR2D2 port map( A1 => b(10), A2 => a(11), Z => n688);
   U1079 : EXNOR2D2 port map( A1 => n160, A2 => net11662, Z => product(22));
   U1080 : EXNOR2DL port map( A1 => b(9), A2 => a(5), Z => n740);
   U1081 : EXNOR2DL port map( A1 => b(9), A2 => a(7), Z => n723);
   U1082 : EXOR2D1 port map( A1 => n573, A2 => n425, Z => n977);
   U1083 : EXOR2D1 port map( A1 => n977, A2 => n588, Z => n410);
   U1084 : OAI22D1 port map( A1 => n708, A2 => n30, B1 => n978, B2 => n28, Z =>
                           n573);
   U1085 : EXNOR2DL port map( A1 => b(2), A2 => a(15), Z => n662);
   U1086 : EXNOR2DL port map( A1 => b(2), A2 => a(11), Z => n696);
   U1087 : EXNOR2DL port map( A1 => b(12), A2 => a(3), Z => n754);
   U1088 : EXNOR2DL port map( A1 => b(12), A2 => a(9), Z => n703);
   U1089 : EXNOR2DL port map( A1 => b(12), A2 => a(11), Z => n686);
   U1090 : EXNOR2DL port map( A1 => b(12), A2 => a(13), Z => n669);
   U1091 : EXNOR2DL port map( A1 => b(12), A2 => a(15), Z => n652);
   U1092 : EXNOR2D2 port map( A1 => b(5), A2 => a(13), Z => n676);
   U1093 : EXNOR2D2 port map( A1 => b(12), A2 => a(7), Z => n720);
   U1094 : EXOR2D4 port map( A1 => n188, A2 => n65, Z => product(18));
   U1095 : ADHALFD2 port map( A => n546, B => n514, CO => n451, S => n452);
   U1096 : EXNOR2DL port map( A1 => b(8), A2 => a(13), Z => n673);
   U1097 : EXNOR2DL port map( A1 => b(8), A2 => a(1), Z => n775);
   U1098 : EXNOR2DL port map( A1 => b(8), A2 => a(3), Z => n758);
   U1099 : OAI22DL port map( A1 => n668, A2 => n42, B1 => n667, B2 => n40, Z =>
                           n533);
   U1100 : OAI22D2 port map( A1 => n684, A2 => n36, B1 => n683, B2 => n34, Z =>
                           n549);
   U1101 : OAI22DL port map( A1 => n701, A2 => n30, B1 => n700, B2 => n28, Z =>
                           n566);
   U1102 : OAI22D2 port map( A1 => n718, A2 => n24, B1 => n717, B2 => n22, Z =>
                           n583);
   U1103 : EXNOR2DL port map( A1 => b(7), A2 => a(1), Z => n776);
   U1104 : EXNOR2DL port map( A1 => b(7), A2 => a(3), Z => n759);
   U1105 : EXNOR2DL port map( A1 => b(7), A2 => a(15), Z => n657);
   U1106 : EXNOR2DL port map( A1 => a(7), A2 => b(14), Z => n718);
   U1107 : EXNOR2DL port map( A1 => b(7), A2 => a(5), Z => n742);
   U1108 : EXNOR2DL port map( A1 => b(8), A2 => a(9), Z => n978);
   U1109 : EXNOR2D2 port map( A1 => b(15), A2 => a(1), Z => n768);
   U1110 : EXOR3D1 port map( A1 => n419, A2 => n410, A3 => n408, Z => n404);
   U1111 : NAN2D1 port map( A1 => n419, A2 => n410, Z => n980);
   U1112 : NAN2D1 port map( A1 => n419, A2 => n408, Z => n981);
   U1113 : NAN2D1 port map( A1 => n410, A2 => n408, Z => n982);
   U1114 : NAN3D2 port map( A1 => n980, A2 => n981, A3 => n982, Z => n403);
   U1115 : NAN2DL port map( A1 => n417, A2 => n404, Z => n983);
   U1116 : NAN3D1 port map( A1 => net11507, A2 => n983, A3 => net11509, Z => 
                           n401);
   U1117 : NAN2D1 port map( A1 => n449, A2 => n590, Z => n986);
   U1118 : NAN3D2 port map( A1 => n984, A2 => n986, A3 => n985, Z => n435);
   U1119 : ADFULD1 port map( A => n619, B => n437, CI => n435, CO => n419, S =>
                           n420);
   U1120 : EXNOR2D2 port map( A1 => b(5), A2 => a(9), Z => n710);
   U1121 : EXNOR2DL port map( A1 => a(1), A2 => b(9), Z => n774);
   U1122 : EXNOR2DL port map( A1 => b(9), A2 => a(11), Z => n689);
   U1123 : EXNOR2DL port map( A1 => b(6), A2 => a(5), Z => n743);
   U1124 : EXNOR2D2 port map( A1 => b(6), A2 => a(13), Z => n675);
   U1125 : EXNOR2D2 port map( A1 => b(14), A2 => a(1), Z => n769);
   U1126 : EXNOR2DL port map( A1 => b(14), A2 => a(5), Z => n735);
   U1127 : EXNOR2DL port map( A1 => b(14), A2 => a(3), Z => n752);
   U1128 : NAN2D2 port map( A1 => n402, A2 => n415, Z => n201);
   U1129 : EXNOR2D2 port map( A1 => b(10), A2 => a(5), Z => n739);
   U1130 : EXNOR2DL port map( A1 => b(2), A2 => a(9), Z => n713);
   U1131 : EXNOR2DL port map( A1 => b(2), A2 => a(13), Z => n679);
   U1132 : INVDL port map( A => n53, Z => n128);
   U1133 : NOR2DL port map( A1 => n53, A2 => n108, Z => n106);
   U1134 : AND2DL port map( A1 => n283, A2 => n168, Z => n989);
   U1135 : NAN2DL port map( A1 => n284, A2 => net12095, Z => n63);
   U1136 : NAN2M1DL port map( A1 => net12055, A2 => net11746, Z => n65);
   U1137 : EXNOR2D1 port map( A1 => n987, A2 => net11172, Z => product(19));
   U1138 : AOI21DL port map( A1 => n182, A2 => n202, B => n183, Z => n987);
   U1139 : INVDL port map( A => n173, Z => n171);
   U1140 : INVDL port map( A => n117, Z => n279);
   U1141 : INVDL port map( A => n118, Z => n124);
   U1142 : NAN2M1DL port map( A1 => n103, A2 => n104, Z => n56);
   U1143 : EXNOR2D2 port map( A1 => n114, A2 => n988, Z => product(26));
   U1144 : AND2DL port map( A1 => n278, A2 => n113, Z => n988);
   U1145 : NAN2M1DL port map( A1 => n92, A2 => n93, Z => n55);
   U1146 : NAN2DL port map( A1 => n322, A2 => n327, Z => n139);
   U1147 : INVDL port map( A => n112, Z => n278);
   U1148 : NOR2DL port map( A1 => n112, A2 => n103, Z => n101);
   U1149 : EXNOR2D2 port map( A1 => net11025, A2 => n366, Z => n364);
   U1150 : AND2DL port map( A1 => n502, A2 => n505, Z => n1003);
   U1151 : NOR2D1 port map( A1 => n506, A2 => n509, Z => n257);
   U1152 : OR2DL port map( A1 => n510, A2 => n645, Z => n1004);
   U1153 : AND2DL port map( A1 => n647, A2 => n632, Z => n1007);
   U1154 : OAI22D1 port map( A1 => n754, A2 => n12, B1 => n753, B2 => n9, Z => 
                           n619);
   U1155 : OAI22DL port map( A1 => n670, A2 => n42, B1 => n669, B2 => n40, Z =>
                           n535);
   U1156 : OAI22DL port map( A1 => n653, A2 => n48, B1 => n652, B2 => n46, Z =>
                           n524);
   U1157 : OAI22DL port map( A1 => n652, A2 => n48, B1 => n651, B2 => n46, Z =>
                           n523);
   U1158 : OA22DL port map( A1 => n650, A2 => n48, B1 => n649, B2 => n46, Z => 
                           n1010);
   U1159 : NOR2DL port map( A1 => n53, A2 => n97, Z => n95);
   U1160 : INVDL port map( A => n172, Z => n284);
   U1161 : NOR2DL port map( A1 => n53, A2 => n997, Z => n86);
   U1162 : NAN2D1 port map( A1 => n279, A2 => n278, Z => n108);
   U1163 : NAN2DL port map( A1 => n101, A2 => n279, Z => n97);
   U1164 : NOR2DL port map( A1 => n53, A2 => n117, Z => n115);
   U1165 : OR2D1 port map( A1 => n442, A2 => n453, Z => n990);
   U1166 : NOR2D1 port map( A1 => n402, A2 => n415, Z => n200);
   U1167 : OA21M20D1 port map( A1 => n124, A2 => n278, B => n113, Z => n109);
   U1168 : NAN2D1 port map( A1 => n991, A2 => n998, Z => n231);
   U1169 : AND2D1 port map( A1 => n454, A2 => n463, Z => n992);
   U1170 : OR2D1 port map( A1 => n454, A2 => n463, Z => n993);
   U1171 : AND2DL port map( A1 => n442, A2 => n453, Z => n994);
   U1172 : NAN2D1 port map( A1 => n344, A2 => n353, Z => n168);
   U1173 : OR2D1 port map( A1 => n322, A2 => n327, Z => net11083);
   U1174 : OR2D1 port map( A1 => n464, A2 => n473, Z => n995);
   U1175 : OA21DL port map( A1 => n100, A2 => n92, B => n93, Z => n996);
   U1176 : NOR2D1 port map( A1 => n316, A2 => n321, Z => n117);
   U1177 : NAN2D1 port map( A1 => n316, A2 => n321, Z => n118);
   U1178 : OR2D1 port map( A1 => n97, A2 => n92, Z => n997);
   U1179 : AND2D1 port map( A1 => n482, A2 => n489, Z => n999);
   U1180 : OR2D1 port map( A1 => n490, A2 => n495, Z => n1000);
   U1181 : NAN2DL port map( A1 => n496, A2 => n501, Z => n250);
   U1182 : NOR2DL port map( A1 => n496, A2 => n501, Z => n249);
   U1183 : AND2D1 port map( A1 => n490, A2 => n495, Z => n1001);
   U1184 : OR2D1 port map( A1 => n502, A2 => n505, Z => n1002);
   U1185 : NAN2DL port map( A1 => n506, A2 => n509, Z => n258);
   U1186 : AND2D1 port map( A1 => n510, A2 => n645, Z => n1005);
   U1187 : NOR2D1 port map( A1 => n312, A2 => n315, Z => n112);
   U1188 : NAN2D1 port map( A1 => n312, A2 => n315, Z => n113);
   U1189 : NOR2D1 port map( A1 => n311, A2 => n308, Z => n103);
   U1190 : NAN2DL port map( A1 => n311, A2 => n308, Z => n104);
   U1191 : NOR2D1 port map( A1 => n307, A2 => n306, Z => n92);
   U1192 : NAN2DL port map( A1 => n307, A2 => n306, Z => n93);
   U1193 : AO21D1 port map( A1 => n18, A2 => n16, B => n734, Z => n599);
   U1194 : AO21D1 port map( A1 => n30, A2 => n28, B => n700, Z => n565);
   U1195 : INVDL port map( A => n333, Z => n334);
   U1196 : AO21D1 port map( A1 => n24, A2 => n22, B => n717, Z => n582);
   U1197 : NAN2D1 port map( A1 => n1009, A2 => n84, Z => n54);
   U1198 : NAN2DL port map( A1 => n305, A2 => n1010, Z => n84);
   U1199 : INVDL port map( A => n319, Z => n320);
   U1200 : AO21D1 port map( A1 => n36, A2 => n34, B => n683, Z => n548);
   U1201 : NAN2DL port map( A1 => n646, A2 => n512, Z => n266);
   U1202 : NOR2DL port map( A1 => n646, A2 => n512, Z => n265);
   U1203 : AND2D1 port map( A1 => n648, A2 => n520, Z => n1008);
   U1204 : INVDL port map( A => n309, Z => n310);
   U1205 : AO21D1 port map( A1 => n42, A2 => n40, B => n666, Z => n532);
   U1206 : OR2D1 port map( A1 => n305, A2 => n1010, Z => n1009);
   U1207 : INVD1 port map( A => a(13), Z => n826);
   U1208 : EXNOR2DL port map( A1 => b(5), A2 => a(7), Z => n727);
   U1209 : INVD1 port map( A => a(11), Z => n827);
   U1210 : EXNOR2DL port map( A1 => b(10), A2 => a(1), Z => n773);
   U1211 : INVD1 port map( A => a(9), Z => n828);
   U1212 : ADHALFDL port map( A => n597, B => n517, CO => n499, S => n500);
   U1213 : INVD1 port map( A => a(7), Z => n829);
   U1214 : ADHALFDL port map( A => n614, B => n518, CO => n507, S => n508);
   U1215 : INVD1 port map( A => a(5), Z => n830);
   U1216 : ADHALFDL port map( A => n631, B => n519, CO => n511, S => n512);
   U1217 : INVD1 port map( A => a(3), Z => n831);
   U1218 : EXNOR2D1 port map( A1 => a(13), A2 => a(14), Z => n46);
   U1219 : NAN2D1 port map( A1 => n801, A2 => n46, Z => n48);
   U1220 : EXNOR2D1 port map( A1 => a(5), A2 => a(6), Z => n22);
   U1221 : NAN2D1 port map( A1 => n805, A2 => n22, Z => n24);
   U1222 : EXNOR2D1 port map( A1 => a(1), A2 => a(2), Z => n9);
   U1223 : NAN2D1 port map( A1 => n807, A2 => n9, Z => n12);
   U1224 : EXNOR2D1 port map( A1 => a(3), A2 => a(4), Z => n16);
   U1225 : NAN2D1 port map( A1 => n806, A2 => n16, Z => n18);
   U1226 : NAN2D1 port map( A1 => n808, A2 => n824, Z => n6);
   U1227 : INVD1 port map( A => a(1), Z => n832);
   U1228 : INVDL port map( A => n201, Z => n199);
   U1229 : EXNOR2DL port map( A1 => b(1), A2 => a(1), Z => n782);
   U1230 : EXNOR2DL port map( A1 => b(1), A2 => a(3), Z => n765);
   U1231 : EXNOR2DL port map( A1 => b(1), A2 => a(5), Z => n748);
   U1232 : EXNOR2DL port map( A1 => b(1), A2 => a(7), Z => n731);
   U1233 : AOI21DL port map( A1 => n202, A2 => net12127, B => net12033, Z => 
                           n188);
   U1234 : INVDL port map( A => n913, Z => n285);
   U1235 : OAI21DL port map( A1 => n997, A2 => net12183, B => n996, Z => n87);
   U1236 : OAI21DL port map( A1 => net12183, A2 => n97, B => n100, Z => n96);
   U1237 : EXNOR2DL port map( A1 => b(5), A2 => a(1), Z => n778);
   U1238 : EXNOR2DL port map( A1 => b(5), A2 => a(3), Z => n761);
   U1239 : EXNOR2DL port map( A1 => b(5), A2 => a(15), Z => n659);
   U1240 : EXNOR2DL port map( A1 => b(5), A2 => a(5), Z => n744);
   U1241 : EXNOR2DL port map( A1 => b(15), A2 => a(3), Z => n751);
   U1242 : EXNOR2DL port map( A1 => b(15), A2 => a(7), Z => n717);
   U1243 : EXNOR2DL port map( A1 => b(15), A2 => a(9), Z => n700);
   U1244 : EXNOR2DL port map( A1 => b(15), A2 => a(11), Z => n683);
   U1245 : EXNOR2DL port map( A1 => b(15), A2 => a(13), Z => n666);
   U1246 : EXNOR2DL port map( A1 => b(15), A2 => a(15), Z => n649);
   U1247 : EXNOR2DL port map( A1 => b(10), A2 => a(15), Z => n654);
   U1248 : EXNOR2DL port map( A1 => b(10), A2 => a(9), Z => n705);
   U1249 : NAN2DL port map( A1 => n366, A2 => net12257, Z => n1011);
   U1250 : NAN2DL port map( A1 => n366, A2 => n368, Z => n1012);
   U1251 : NAN2DL port map( A1 => n368, A2 => net12257, Z => n1013);
   U1252 : NAN3D1 port map( A1 => n1011, A2 => n1013, A3 => n1012, Z => n363);
   U1253 : NOR2D1 port map( A1 => n354, A2 => n363, Z => n172);
   U1254 : NAN2D1 port map( A1 => n388, A2 => n401, Z => n196);
   U1255 : EXNOR2DL port map( A1 => b(14), A2 => a(15), Z => n650);
   U1256 : EXNOR2DL port map( A1 => b(14), A2 => a(13), Z => n667);
   U1257 : EXNOR2DL port map( A1 => b(14), A2 => a(11), Z => n684);
   U1258 : EXNOR2DL port map( A1 => b(14), A2 => a(9), Z => n701);
   U1259 : OAI21DL port map( A1 => n52, A2 => n117, B => n118, Z => n116);
   U1260 : INVDL port map( A => net12183, Z => n129);
   U1261 : OAI21DL port map( A1 => n52, A2 => n108, B => n109, Z => n107);
   U1262 : AOI21D1 port map( A1 => net12285, A2 => n141, B => n142, Z => n140);
   U1263 : AOI21DL port map( A1 => net12285, A2 => n86, B => n87, Z => n85);
   U1264 : AOI21DL port map( A1 => net12285, A2 => n95, B => n96, Z => n94);
   U1265 : AOI21DL port map( A1 => net12285, A2 => n115, B => n116, Z => n114);
   U1266 : NAN2DL port map( A1 => n288, A2 => n201, Z => n67);
   U1267 : EXNOR2DL port map( A1 => b(13), A2 => a(15), Z => n651);
   U1268 : EXNOR2DL port map( A1 => b(13), A2 => a(13), Z => n668);
   U1269 : EXNOR2DL port map( A1 => b(13), A2 => a(11), Z => n685);
   U1270 : EXNOR2DL port map( A1 => b(13), A2 => a(9), Z => n702);
   U1271 : EXNOR2DL port map( A1 => b(13), A2 => a(7), Z => n719);
   U1272 : EXNOR2D2 port map( A1 => b(13), A2 => a(5), Z => n736);
   U1273 : EXNOR2DL port map( A1 => n914, A2 => a(15), Z => n653);
   U1274 : EXNOR2DL port map( A1 => n914, A2 => a(13), Z => n670);
   U1275 : EXNOR2DL port map( A1 => b(11), A2 => a(11), Z => n687);
   U1276 : EXNOR2DL port map( A1 => b(11), A2 => a(1), Z => n772);

end hier_sec_par_16_5;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_siso_gen.all;

architecture hier_sec_par_16_5 of siso_gen_DW01_add_13 is

   component INVBD2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D4
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21M20DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVDL
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFDL
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21M10D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n9, n10, n12, n13, n14, n15, n16, n17, 
      n19, n20, n21, n22, n23, n26, n27, n28, n30, n31, n32, n33, n34, n35, n36
      , n37, n38, n39, n42, n43, n44, n45, n47, n50, n51, n52, n53, n55, n56, 
      n58, n59, n71, n80, n81, n82, n89, n90, n91, n92, n93, n94, n95, n96, n97
      , n98, n100, n101, n102, n104, n105, n106, n107, n108, n112, n113, n115, 
      n117, n118, n119, n120, n129, net11329, net11441, net11439, net11615, 
      net11859, net12242, net12241, n78, n60, net12276, net11486, net11440, n88
      , n87, n86, n84, n8, n79, n75, n73, n70, n66, n64, n63, n62, n61, n122, 
      n83, n72, n67, n65, n123, n187, n188, n189, n190, n191, n192, n193, n194,
      n195, n196, n197, n198, n199, n200, n201, n202 : std_logic;

begin
   
   U10 : OAI21D1 port map( A1 => n31, A2 => n23, B => n26, Z => n22);
   U15 : NOR2D2 port map( A1 => B(14), A2 => A(14), Z => n23);
   U22 : AOI21D1 port map( A1 => n32, A2 => n45, B => n33, Z => n31);
   U37 : NOR2D2 port map( A1 => B(12), A2 => A(12), Z => n39);
   U46 : OAI21D1 port map( A1 => n50, A2 => n56, B => n51, Z => n45);
   U49 : NOR2D2 port map( A1 => B(11), A2 => A(11), Z => n50);
   U58 : NAN2D2 port map( A1 => B(10), A2 => A(10), Z => n56);
   U106 : NOR2D2 port map( A1 => B(5), A2 => A(5), Z => n89);
   U109 : OAI21D1 port map( A1 => n94, A2 => n92, B => n93, Z => n91);
   U112 : NOR2D2 port map( A1 => B(4), A2 => A(4), Z => n92);
   U113 : NAN2D2 port map( A1 => B(4), A2 => A(4), Z => n93);
   U116 : OAI21D1 port map( A1 => n96, A2 => n108, B => n97, Z => n95);
   U123 : NOR2D2 port map( A1 => B(3), A2 => A(3), Z => n100);
   U131 : NOR2D2 port map( A1 => B(2), A2 => A(2), Z => n105);
   U132 : NAN2D2 port map( A1 => B(2), A2 => A(2), Z => n106);
   U89 : NOR2D2 port map( A1 => B(7), A2 => A(7), Z => n78);
   U103 : OAI21D1 port map( A1 => n89, A2 => n93, B => n90, Z => n88);
   U101 : AOI21D1 port map( A1 => n95, A2 => n87, B => n88, Z => n86);
   U62 : AOI21D1 port map( A1 => n60, A2 => n73, B => n61, Z => n59);
   U67 : NOR2D2 port map( A1 => B(9), A2 => A(9), Z => n62);
   U86 : OAI21D1 port map( A1 => n78, A2 => n84, B => n79, Z => n73);
   U63 : NOR2D2 port map( A1 => n67, A2 => n62, Z => n60);
   U77 : NOR2D2 port map( A1 => B(8), A2 => A(8), Z => n67);
   U151 : NOR2D1 port map( A1 => B(13), A2 => A(13), Z => n34);
   U152 : OAI21D1 port map( A1 => n75, A2 => net12276, B => n70, Z => n66);
   U153 : NAN2M1D1 port map( A1 => B(1), A2 => n194, Z => n187);
   U154 : NAN2M1DL port map( A1 => B(1), A2 => n194, Z => n202);
   U155 : AND2D1 port map( A1 => n72, A2 => n123, Z => n65);
   U156 : INVD1 port map( A => A(7), Z => n192);
   U157 : NAN2DL port map( A1 => n122, A2 => n63, Z => n8);
   U158 : NAN2DL port map( A1 => n120, A2 => n51, Z => n6);
   U159 : NAN2DL port map( A1 => n118, A2 => n35, Z => n4);
   U160 : INVD1 port map( A => A(1), Z => n194);
   U161 : OR2D1 port map( A1 => A(7), A2 => net12242, Z => n188);
   U162 : INVD2 port map( A => n58, Z => net11439);
   U163 : INVD1 port map( A => n115, Z => n113);
   U164 : INVD1 port map( A => n108, Z => n107);
   U165 : INVDL port map( A => n129, Z => n189);
   U166 : INVD1 port map( A => n189, Z => n190);
   U167 : INVBD2 port map( A => n100, Z => n98);
   U168 : NOR2D2 port map( A1 => B(10), A2 => A(10), Z => n55);
   U169 : AOI21M10D1 port map( A1 => n55, A2 => n1, B => n191, Z => n52);
   U170 : INVDL port map( A => n56, Z => n191);
   U171 : EXNOR2D2 port map( A1 => n91, A2 => n12, Z => SUM(5));
   U172 : AOI21DL port map( A1 => n65, A2 => net11440, B => n66, Z => n64);
   U173 : INVDL port map( A => n67, Z => n123);
   U174 : NAN2DL port map( A1 => n123, A2 => n70, Z => n9);
   U175 : NOR2D1 port map( A1 => n78, A2 => n83, Z => n72);
   U176 : NAN2D2 port map( A1 => n72, A2 => n60, Z => n58);
   U177 : AOI21DL port map( A1 => net11440, A2 => n72, B => net11486, Z => n71)
                           ;
   U178 : BUFDL port map( A => n67, Z => net12276);
   U179 : INVDL port map( A => n83, Z => n81);
   U180 : NAN2D1 port map( A1 => A(8), A2 => B(8), Z => n70);
   U181 : NOR2D2 port map( A1 => B(6), A2 => A(6), Z => n83);
   U182 : NAN2DL port map( A1 => A(6), A2 => B(6), Z => net11615);
   U183 : NAN2D1 port map( A1 => B(6), A2 => A(6), Z => n84);
   U184 : EXOR2D4 port map( A1 => n64, A2 => n8, Z => SUM(9));
   U185 : INVDL port map( A => n62, Z => n122);
   U186 : INVDL port map( A => n73, Z => n75);
   U187 : INVDL port map( A => n75, Z => net11486);
   U188 : INVD2 port map( A => n86, Z => net11440);
   U189 : AOI21DL port map( A1 => net11440, A2 => n81, B => n82, Z => n80);
   U190 : NAN2D2 port map( A1 => net11439, A2 => net11440, Z => net11441);
   U191 : NAN2D1 port map( A1 => B(9), A2 => A(9), Z => n63);
   U192 : OAI21DL port map( A1 => n70, A2 => n62, B => n63, Z => n61);
   U193 : NAN2M1DL port map( A1 => n192, A2 => B(7), Z => n79);
   U194 : EXOR2D4 port map( A1 => n86, A2 => net11329, Z => SUM(6));
   U195 : NOR2D1 port map( A1 => n89, A2 => n92, Z => n87);
   U196 : INVDL port map( A => B(7), Z => net12241);
   U197 : NAN2DL port map( A1 => A(7), A2 => net12242, Z => net11859);
   U198 : INVDL port map( A => net12241, Z => net12242);
   U199 : INVDL port map( A => n47, Z => n193);
   U200 : NAN2DL port map( A1 => n119, A2 => n42, Z => n5);
   U201 : OAI21DL port map( A1 => n47, A2 => n39, B => n42, Z => n38);
   U202 : OAI21DL port map( A1 => n34, A2 => n42, B => n35, Z => n33);
   U203 : INVD2 port map( A => n106, Z => n104);
   U204 : INVDL port map( A => net11615, Z => n82);
   U205 : NAN2M1DL port map( A1 => n194, A2 => B(1), Z => n112);
   U206 : NAN2D1 port map( A1 => n117, A2 => n26, Z => n3);
   U207 : AOI21D1 port map( A1 => n107, A2 => n190, B => n104, Z => n102);
   U208 : NAN2D1 port map( A1 => n199, A2 => n15, Z => n197);
   U209 : NAN2D2 port map( A1 => n196, A2 => n195, Z => n198);
   U210 : NAN2D2 port map( A1 => n198, A2 => n197, Z => SUM(2));
   U211 : INVD2 port map( A => n15, Z => n195);
   U212 : INVD1 port map( A => n199, Z => n196);
   U213 : INVDL port map( A => n108, Z => n199);
   U214 : NAN2D1 port map( A1 => n81, A2 => net11615, Z => net11329);
   U215 : NAN2D1 port map( A1 => n129, A2 => n98, Z => n96);
   U216 : INVDL port map( A => n17, Z => SUM(0));
   U217 : NAN2D2 port map( A1 => net11441, A2 => n59, Z => n1);
   U218 : NAN2DL port map( A1 => n200, A2 => n115, Z => n17);
   U219 : OR2DL port map( A1 => B(0), A2 => A(0), Z => n200);
   U220 : INVDL port map( A => n30, Z => n28);
   U221 : NAN2M1DL port map( A1 => n89, A2 => n90, Z => n12);
   U222 : INVDL port map( A => n55, Z => n53);
   U223 : NAN2M1DL port map( A1 => n92, A2 => n93, Z => n13);
   U224 : NOR2DL port map( A1 => n30, A2 => n23, Z => n21);
   U225 : NAN2D1 port map( A1 => B(13), A2 => A(13), Z => n35);
   U226 : NAN2D1 port map( A1 => B(14), A2 => A(14), Z => n26);
   U227 : NAN2D1 port map( A1 => n32, A2 => n44, Z => n30);
   U228 : INVDL port map( A => n50, Z => n120);
   U229 : INVDL port map( A => n23, Z => n117);
   U230 : OA21M20D1 port map( A1 => n187, A2 => n113, B => n112, Z => n108);
   U231 : OA21M20D1 port map( A1 => n98, A2 => n104, B => n101, Z => n97);
   U232 : INVDL port map( A => n39, Z => n119);
   U233 : INVDL port map( A => n34, Z => n118);
   U234 : NOR2M1DL port map( A1 => n44, A2 => n39, Z => n37);
   U235 : INVDL port map( A => n45, Z => n47);
   U236 : NAN2D1 port map( A1 => n201, A2 => n19, Z => n2);
   U237 : NAN2DL port map( A1 => B(15), A2 => A(15), Z => n19);
   U238 : NAN2D1 port map( A1 => B(11), A2 => A(11), Z => n51);
   U239 : NAN2D1 port map( A1 => A(0), A2 => B(0), Z => n115);
   U240 : NAN2D1 port map( A1 => B(12), A2 => A(12), Z => n42);
   U241 : OR2D1 port map( A1 => B(15), A2 => A(15), Z => n201);
   U242 : NAN2D1 port map( A1 => B(5), A2 => A(5), Z => n90);
   U243 : AOI21DL port map( A1 => n1, A2 => n37, B => n38, Z => n36);
   U244 : INVD1 port map( A => n95, Z => n94);
   U245 : EXNOR2D1 port map( A1 => n1, A2 => n7, Z => SUM(10));
   U246 : OA21M20DL port map( A1 => n1, A2 => n28, B => n31, Z => n27);
   U247 : NOR2D1 port map( A1 => n39, A2 => n34, Z => n32);
   U248 : NAN2DL port map( A1 => n53, A2 => n56, Z => n7);
   U249 : NAN2DL port map( A1 => n202, A2 => n112, Z => n16);
   U250 : NAN2D1 port map( A1 => n188, A2 => net11859, Z => n10);
   U251 : EXNOR2D2 port map( A1 => n16, A2 => n113, Z => SUM(1));
   U252 : EXOR2D4 port map( A1 => n94, A2 => n13, Z => SUM(4));
   U253 : NAN2D1 port map( A1 => A(3), A2 => B(3), Z => n101);
   U254 : NAN2DL port map( A1 => n101, A2 => n98, Z => n14);
   U255 : NAN2D1 port map( A1 => n129, A2 => n106, Z => n15);
   U256 : EXOR2D4 port map( A1 => n102, A2 => n14, Z => SUM(3));
   U257 : NOR2D1 port map( A1 => n55, A2 => n50, Z => n44);
   U258 : EXOR2D4 port map( A1 => n80, A2 => n10, Z => SUM(7));
   U259 : EXOR2D4 port map( A1 => n36, A2 => n4, Z => SUM(13));
   U260 : EXOR2D4 port map( A1 => n20, A2 => n2, Z => SUM(15));
   U261 : AOI21DL port map( A1 => n1, A2 => n21, B => n22, Z => n20);
   U262 : EXOR2D4 port map( A1 => n71, A2 => n9, Z => SUM(8));
   U263 : EXOR2D4 port map( A1 => n43, A2 => n5, Z => SUM(12));
   U264 : EXOR2D4 port map( A1 => n27, A2 => n3, Z => SUM(14));
   U265 : EXOR2D4 port map( A1 => n52, A2 => n6, Z => SUM(11));
   U266 : AOI21DL port map( A1 => n1, A2 => n44, B => n193, Z => n43);
   U267 : INVBD2 port map( A => n105, Z => n129);

end hier_sec_par_16_5;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_siso_gen.all;

architecture hier_sec_par_16_5 of siso_gen_DW01_add_12 is

   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INVDL
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFDL
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21M20DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M20DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n19, n20, n21, n22
      , n23, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, 
      n39, n42, n43, n44, n45, n47, n50, n51, n52, n53, n55, n56, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n70, n71, n72, n73, n75, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n102, n103, n104, n105, n107, n109, n110, n112, 
      n116, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, 
      n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, 
      n202, n203, n205, n206, n207, n208, n209 : std_logic;

begin
   
   U15 : NOR2D2 port map( A1 => B(14), A2 => A(14), Z => n23);
   U22 : AOI21D1 port map( A1 => n32, A2 => n45, B => n33, Z => n31);
   U24 : OAI21D1 port map( A1 => n34, A2 => n42, B => n35, Z => n33);
   U27 : NOR2D2 port map( A1 => B(13), A2 => A(13), Z => n34);
   U37 : NOR2D2 port map( A1 => B(12), A2 => A(12), Z => n39);
   U40 : AOI21D1 port map( A1 => n1, A2 => n44, B => n189, Z => n43);
   U46 : OAI21D1 port map( A1 => n50, A2 => n56, B => n51, Z => n45);
   U49 : NOR2D2 port map( A1 => B(11), A2 => A(11), Z => n50);
   U59 : EXOR2D1 port map( A1 => n64, A2 => n8, Z => SUM(9));
   U60 : OAI21D1 port map( A1 => n188, A2 => n58, B => n59, Z => n1);
   U62 : AOI21D1 port map( A1 => n60, A2 => n73, B => n61, Z => n59);
   U67 : NOR2D2 port map( A1 => B(9), A2 => A(9), Z => n62);
   U69 : EXOR2D1 port map( A1 => n71, A2 => n9, Z => SUM(8));
   U70 : AOI21D1 port map( A1 => n85, A2 => n65, B => n66, Z => n64);
   U79 : EXOR2D1 port map( A1 => n80, A2 => n10, Z => SUM(7));
   U86 : OAI21D1 port map( A1 => n78, A2 => n84, B => n79, Z => n73);
   U89 : NOR2D2 port map( A1 => B(7), A2 => A(7), Z => n78);
   U92 : AOI21D1 port map( A1 => n85, A2 => n81, B => n82, Z => n80);
   U99 : EXNOR2D1 port map( A1 => n91, A2 => n12, Z => SUM(5));
   U103 : OAI21D1 port map( A1 => n89, A2 => n93, B => n90, Z => n88);
   U106 : NOR2D2 port map( A1 => B(5), A2 => A(5), Z => n89);
   U108 : EXOR2D1 port map( A1 => n13, A2 => n94, Z => SUM(4));
   U112 : NOR2D2 port map( A1 => B(4), A2 => A(4), Z => n92);
   U116 : OAI21D1 port map( A1 => n98, A2 => n96, B => n97, Z => n95);
   U119 : NOR2D2 port map( A1 => B(3), A2 => A(3), Z => n96);
   U122 : AOI21D1 port map( A1 => n205, A2 => n103, B => n202, Z => n98);
   U129 : EXOR2D1 port map( A1 => n16, A2 => n107, Z => SUM(1));
   U130 : OAI21D1 port map( A1 => n104, A2 => n107, B => n105, Z => n103);
   U143 : BUFDL port map( A => n78, Z => n179);
   U144 : OA21DL port map( A1 => n89, A2 => n93, B => n90, Z => n180);
   U145 : NAN2D1 port map( A1 => B(5), A2 => A(5), Z => n90);
   U146 : EXNOR2DL port map( A1 => n85, A2 => n11, Z => SUM(6));
   U147 : NOR2M1DL port map( A1 => n72, A2 => n195, Z => n65);
   U148 : BUFDL port map( A => n72, Z => n182);
   U149 : BUFDL port map( A => B(8), Z => n181);
   U150 : NAN2D1 port map( A1 => B(7), A2 => A(7), Z => n79);
   U151 : OAI21M20DL port map( A1 => n95, A2 => n87, B => n180, Z => n85);
   U152 : OR2DL port map( A1 => B(0), A2 => A(0), Z => n183);
   U153 : NAN2D1 port map( A1 => B(10), A2 => A(10), Z => n56);
   U154 : INVD1 port map( A => A(9), Z => n187);
   U155 : OR2D1 port map( A1 => B(15), A2 => A(15), Z => n184);
   U156 : INVD1 port map( A => n186, Z => n94);
   U157 : EXNOR2DL port map( A1 => n200, A2 => n185, Z => SUM(10));
   U158 : AND2DL port map( A1 => n53, A2 => n201, Z => n185);
   U159 : INVD1 port map( A => n43, Z => n196);
   U160 : NAN2DL port map( A1 => n43, A2 => n197, Z => n198);
   U161 : NAN2D1 port map( A1 => n196, A2 => n5, Z => n199);
   U162 : AOI21DL port map( A1 => n1, A2 => n28, B => n29, Z => n27);
   U163 : NAN2D2 port map( A1 => B(4), A2 => A(4), Z => n93);
   U164 : EXOR2DL port map( A1 => n14, A2 => n98, Z => SUM(3));
   U165 : OAI21DL port map( A1 => n98, A2 => n96, B => n97, Z => n186);
   U166 : OA21M20DL port map( A1 => n206, A2 => n53, B => n201, Z => n52);
   U167 : NAN2M1DL port map( A1 => n187, A2 => B(9), Z => n63);
   U168 : NAN2D1 port map( A1 => A(13), A2 => B(13), Z => n35);
   U169 : AOI21DL port map( A1 => n95, A2 => n87, B => n88, Z => n188);
   U170 : AOI21DL port map( A1 => n95, A2 => n87, B => n88, Z => n86);
   U171 : BUFDL port map( A => n45, Z => n189);
   U172 : NOR2DL port map( A1 => A(3), A2 => B(3), Z => n190);
   U173 : NAN2D1 port map( A1 => n44, A2 => n32, Z => n30);
   U174 : INVDL port map( A => n39, Z => n191);
   U175 : INVD1 port map( A => n191, Z => n192);
   U176 : NAN2D1 port map( A1 => B(1), A2 => A(1), Z => n105);
   U177 : OAI21D1 port map( A1 => n31, A2 => n23, B => n26, Z => n22);
   U178 : NAN2D1 port map( A1 => B(6), A2 => A(6), Z => n84);
   U179 : NOR2D1 port map( A1 => B(6), A2 => A(6), Z => n83);
   U180 : NAN2D1 port map( A1 => B(8), A2 => A(8), Z => n70);
   U181 : EXNOR2DL port map( A1 => n27, A2 => n193, Z => SUM(14));
   U182 : AND2D1 port map( A1 => n109, A2 => n26, Z => n193);
   U183 : NOR2DL port map( A1 => n181, A2 => A(8), Z => n194);
   U184 : NOR2DL port map( A1 => A(8), A2 => n181, Z => n195);
   U185 : NOR2D1 port map( A1 => B(8), A2 => A(8), Z => n67);
   U186 : OAI21DL port map( A1 => n47, A2 => n192, B => n42, Z => n38);
   U187 : NAN2D1 port map( A1 => n199, A2 => n198, Z => SUM(12));
   U188 : INVDL port map( A => n5, Z => n197);
   U189 : NOR2D1 port map( A1 => n62, A2 => n67, Z => n60);
   U190 : INVDL port map( A => n206, Z => n200);
   U191 : AND2D1 port map( A1 => B(2), A2 => A(2), Z => n202);
   U192 : INVD1 port map( A => n202, Z => n102);
   U193 : NAN2D2 port map( A1 => B(0), A2 => A(0), Z => n107);
   U194 : NAN2D1 port map( A1 => n72, A2 => n60, Z => n58);
   U195 : NAN2DL port map( A1 => B(10), A2 => A(10), Z => n201);
   U196 : NOR2D2 port map( A1 => n39, A2 => n34, Z => n32);
   U197 : EXNOR2DL port map( A1 => n15, A2 => n103, Z => SUM(2));
   U198 : AOI21D1 port map( A1 => n85, A2 => n182, B => n203, Z => n71);
   U199 : INVDL port map( A => n75, Z => n203);
   U200 : NAN2D1 port map( A1 => B(11), A2 => A(11), Z => n51);
   U201 : OAI21DL port map( A1 => n94, A2 => n92, B => n93, Z => n91);
   U202 : NAN2M1DL port map( A1 => n194, A2 => n70, Z => n9);
   U203 : NAN2M1DL port map( A1 => n62, A2 => n63, Z => n8);
   U204 : INVDL port map( A => n55, Z => n53);
   U205 : NAN2M1DL port map( A1 => n89, A2 => n90, Z => n12);
   U206 : NAN2M1DL port map( A1 => n92, A2 => n93, Z => n13);
   U207 : NAN2M1DL port map( A1 => n190, A2 => n97, Z => n14);
   U208 : NAN2DL port map( A1 => n102, A2 => n205, Z => n15);
   U209 : NAN2M1DL port map( A1 => n39, A2 => n42, Z => n5);
   U210 : NAN2M1DL port map( A1 => n104, A2 => n105, Z => n16);
   U211 : NAN2D1 port map( A1 => B(14), A2 => A(14), Z => n26);
   U212 : AND2DL port map( A1 => n183, A2 => n107, Z => SUM(0));
   U213 : INVDL port map( A => n30, Z => n28);
   U214 : NOR2D1 port map( A1 => n92, A2 => n89, Z => n87);
   U215 : INVDL port map( A => n50, Z => n112);
   U216 : NOR2D1 port map( A1 => n55, A2 => n50, Z => n44);
   U217 : NAN2DL port map( A1 => n81, A2 => n84, Z => n11);
   U218 : INVDL port map( A => n83, Z => n81);
   U219 : INVDL port map( A => n84, Z => n82);
   U220 : INVDL port map( A => n23, Z => n109);
   U221 : INVDL port map( A => n34, Z => n110);
   U222 : OR2D1 port map( A1 => B(2), A2 => A(2), Z => n205);
   U223 : NOR2DL port map( A1 => n30, A2 => n23, Z => n21);
   U224 : NOR2D1 port map( A1 => B(10), A2 => A(10), Z => n55);
   U225 : NAN2D1 port map( A1 => A(3), A2 => B(3), Z => n97);
   U226 : NOR2M1DL port map( A1 => n44, A2 => n192, Z => n37);
   U227 : NOR2D1 port map( A1 => B(1), A2 => A(1), Z => n104);
   U228 : NAN2D1 port map( A1 => B(12), A2 => A(12), Z => n42);
   U229 : NAN2D1 port map( A1 => B(15), A2 => A(15), Z => n19);
   U230 : NAN2DL port map( A1 => n116, A2 => n79, Z => n10);
   U231 : INVDL port map( A => n31, Z => n29);
   U232 : OAI21DL port map( A1 => n62, A2 => n70, B => n63, Z => n61);
   U233 : AOI21DL port map( A1 => n21, A2 => n206, B => n22, Z => n20);
   U234 : AOI21DL port map( A1 => n206, A2 => n37, B => n38, Z => n36);
   U235 : NOR2D1 port map( A1 => n78, A2 => n83, Z => n72);
   U236 : INVDL port map( A => n179, Z => n116);
   U237 : OAI21DL port map( A1 => n75, A2 => n194, B => n70, Z => n66);
   U238 : INVDL port map( A => n45, Z => n47);
   U239 : INVDL port map( A => n73, Z => n75);
   U240 : OAI21D1 port map( A1 => n58, A2 => n86, B => n59, Z => n206);
   U241 : EXNOR2DL port map( A1 => n52, A2 => n207, Z => SUM(11));
   U242 : AND2DL port map( A1 => n112, A2 => n51, Z => n207);
   U243 : EXNOR2DL port map( A1 => n36, A2 => n208, Z => SUM(13));
   U244 : AND2DL port map( A1 => n110, A2 => n35, Z => n208);
   U245 : EXNOR2D1 port map( A1 => n20, A2 => n209, Z => SUM(15));
   U246 : AND2D1 port map( A1 => n184, A2 => n19, Z => n209);

end hier_sec_par_16_5;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_siso_gen.all;

architecture hier_sec_par_16_5 of siso_gen_DW01_add_11 is

   component OAI21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVDL
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFDL
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M10DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AO21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INVBD32
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n12, n13, n14, n15, n16, n27, n28, n29, n34, 
      n35, n36, n39, n42, n43, n44, n45, n50, n51, n52, n53, n54, n55, n56, n65
      , n66, n70, n71, n75, n78, n79, n80, n81, n82, n83, n84, n85, n89, n90, 
      n91, n92, n93, n94, n95, n96, n97, n98, n100, n102, n103, n104, n105, 
      n107, net9993, net11959, net12025, net12169, net12355, net12354, n88, n87
      , n73, n116, n37, n72, n67, n63, n62, n61, n60, net11588, net11559, n59, 
      n58, n38, n33, n32, n31, n30, n26, n23, n22, n21, n20, n19, n109, n1, 
      n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, 
      n191, n192, n193, n194, n195, n196, n197, n198, n199, n201 : std_logic;

begin
   
   U17 : EXOR2D1 port map( A1 => n36, A2 => n4, Z => SUM(13));
   U29 : EXOR2D1 port map( A1 => n43, A2 => n5, Z => SUM(12));
   U37 : NOR2D2 port map( A1 => B(12), A2 => A(12), Z => n39);
   U46 : OAI21D1 port map( A1 => n199, A2 => n56, B => n51, Z => n45);
   U69 : EXOR2D1 port map( A1 => n71, A2 => n9, Z => SUM(8));
   U89 : NOR2D2 port map( A1 => B(7), A2 => A(7), Z => n78);
   U99 : EXNOR2D1 port map( A1 => n91, A2 => n12, Z => SUM(5));
   U106 : NOR2D2 port map( A1 => B(5), A2 => A(5), Z => n89);
   U112 : NOR2D2 port map( A1 => B(4), A2 => A(4), Z => n92);
   U116 : OAI21D1 port map( A1 => n98, A2 => n96, B => n97, Z => n95);
   U119 : NOR2D2 port map( A1 => B(3), A2 => A(3), Z => n96);
   U122 : AOI21D1 port map( A1 => n103, A2 => n201, B => n100, Z => n98);
   U129 : EXOR2D1 port map( A1 => n16, A2 => n107, Z => SUM(1));
   U130 : OAI21D1 port map( A1 => n104, A2 => n107, B => n105, Z => n103);
   U103 : OAI21D1 port map( A1 => n89, A2 => n93, B => n90, Z => n88);
   U86 : OAI21D1 port map( A1 => n78, A2 => n84, B => n79, Z => n73);
   U67 : NOR2D2 port map( A1 => B(9), A2 => A(9), Z => n62);
   U77 : NOR2D2 port map( A1 => B(8), A2 => A(8), Z => n67);
   U62 : AOI21D1 port map( A1 => n60, A2 => n73, B => n61, Z => n59);
   U22 : AOI21D1 port map( A1 => n32, A2 => n45, B => n33, Z => n31);
   U30 : AOI21D1 port map( A1 => n1, A2 => n37, B => n38, Z => n36);
   U40 : AOI21D1 port map( A1 => n1, A2 => n44, B => n191, Z => n43);
   U60 : OAI21D1 port map( A1 => n58, A2 => n189, B => net11588, Z => n1);
   U10 : OAI21D1 port map( A1 => n31, A2 => n23, B => n26, Z => n22);
   U143 : AOI21D1 port map( A1 => n103, A2 => n201, B => n100, Z => n179);
   U144 : NAN2D1 port map( A1 => n60, A2 => n72, Z => n180);
   U145 : NOR2M1D1 port map( A1 => n181, A2 => B(11), Z => n50);
   U146 : INVBD32 port map( A => A(11), Z => n181);
   U147 : OAI21D1 port map( A1 => n179, A2 => n96, B => n97, Z => n182);
   U148 : NAN2D2 port map( A1 => B(4), A2 => A(4), Z => n93);
   U149 : NOR2D2 port map( A1 => n39, A2 => n34, Z => n32);
   U150 : INVDL port map( A => n189, Z => n85);
   U151 : EXNOR2DL port map( A1 => net9993, A2 => n7, Z => SUM(10));
   U152 : AOI21D1 port map( A1 => net9993, A2 => n53, B => n54, Z => n52);
   U153 : EXNOR2DL port map( A1 => n183, A2 => n8, Z => SUM(9));
   U154 : AO21DL port map( A1 => n85, A2 => n65, B => n66, Z => n183);
   U155 : OAI21DL port map( A1 => n78, A2 => n84, B => n79, Z => n184);
   U156 : OR2DL port map( A1 => B(0), A2 => A(0), Z => n185);
   U157 : AOI21D1 port map( A1 => n87, A2 => n95, B => n88, Z => n189);
   U158 : NAN2M1DL port map( A1 => n199, A2 => n51, Z => n6);
   U159 : INVD1 port map( A => A(2), Z => n188);
   U160 : NAN2D1 port map( A1 => B(15), A2 => A(15), Z => n19);
   U161 : EXOR2D1 port map( A1 => n198, A2 => n14, Z => SUM(3));
   U162 : NAN2M1DL port map( A1 => n96, A2 => n97, Z => n14);
   U163 : EXNOR2D1 port map( A1 => net12025, A2 => n13, Z => SUM(4));
   U164 : INVDL port map( A => net12025, Z => n94);
   U165 : EXNOR2DL port map( A1 => n85, A2 => n186, Z => SUM(6));
   U166 : NAN2D1 port map( A1 => n81, A2 => net11959, Z => n186);
   U167 : AOI21DL port map( A1 => n85, A2 => n81, B => n82, Z => n80);
   U168 : EXNOR2DL port map( A1 => n80, A2 => n187, Z => SUM(7));
   U169 : AND2DL port map( A1 => n116, A2 => n79, Z => n187);
   U170 : NAN2M1D1 port map( A1 => B(2), A2 => n188, Z => n201);
   U171 : NOR2D2 port map( A1 => B(1), A2 => A(1), Z => n104);
   U172 : NAN2D1 port map( A1 => n193, A2 => n6, Z => n196);
   U173 : INVD1 port map( A => n52, Z => n193);
   U174 : AOI21DL port map( A1 => n87, A2 => n182, B => n88, Z => n190);
   U175 : NAN2M1D1 port map( A1 => n104, A2 => n105, Z => n16);
   U176 : NAN2D1 port map( A1 => B(1), A2 => A(1), Z => n105);
   U177 : BUFDL port map( A => n45, Z => n191);
   U178 : EXNOR2DL port map( A1 => n20, A2 => net11559, Z => SUM(15));
   U179 : AND2D1 port map( A1 => n192, A2 => n19, Z => net11559);
   U180 : OR2D1 port map( A1 => B(15), A2 => A(15), Z => n192);
   U181 : AOI21DL port map( A1 => n21, A2 => n1, B => n22, Z => n20);
   U182 : NOR2DL port map( A1 => n30, A2 => n23, Z => n21);
   U183 : AOI21D1 port map( A1 => n60, A2 => n73, B => n61, Z => net11588);
   U184 : INVDL port map( A => n31, Z => n29);
   U185 : OAI21D1 port map( A1 => n42, A2 => n34, B => n35, Z => n33);
   U186 : NOR2D1 port map( A1 => B(14), A2 => A(14), Z => n23);
   U187 : INVDL port map( A => n23, Z => n109);
   U188 : NAN2DL port map( A1 => B(14), A2 => A(14), Z => n26);
   U189 : AND2D1 port map( A1 => n109, A2 => n26, Z => net12169);
   U190 : NAN2D1 port map( A1 => n44, A2 => n32, Z => n30);
   U191 : INVDL port map( A => n30, Z => n28);
   U192 : OAI21D1 port map( A1 => n180, A2 => n190, B => n59, Z => net9993);
   U193 : NAN2D1 port map( A1 => n60, A2 => n72, Z => n58);
   U194 : INVDL port map( A => n73, Z => n75);
   U195 : OAI21M10DL port map( A1 => n45, A2 => n39, B => n42, Z => n38);
   U196 : NAN2M1DL port map( A1 => n39, A2 => n42, Z => n5);
   U197 : NAN2M1DL port map( A1 => n34, A2 => n35, Z => n4);
   U198 : NOR2D2 port map( A1 => n62, A2 => n67, Z => n60);
   U199 : INVDL port map( A => n67, Z => net12354);
   U200 : OAI21D1 port map( A1 => n70, A2 => n62, B => n63, Z => n61);
   U201 : NAN2M1DL port map( A1 => n62, A2 => n63, Z => n8);
   U202 : NAN2D1 port map( A1 => B(8), A2 => A(8), Z => n70);
   U203 : NAN2DL port map( A1 => A(9), A2 => B(9), Z => n63);
   U204 : NOR2D1 port map( A1 => n78, A2 => n83, Z => n72);
   U205 : AOI21D1 port map( A1 => n85, A2 => n72, B => n184, Z => n71);
   U206 : NOR2M1DL port map( A1 => n72, A2 => net12355, Z => n65);
   U207 : INVDL port map( A => n78, Z => n116);
   U208 : INVDL port map( A => n83, Z => n81);
   U209 : NOR2M1DL port map( A1 => n44, A2 => n39, Z => n37);
   U210 : NOR2D1 port map( A1 => n92, A2 => n89, Z => n87);
   U211 : BUFDL port map( A => n182, Z => net12025);
   U212 : NAN2M1DL port map( A1 => n89, A2 => n90, Z => n12);
   U213 : OAI21DL port map( A1 => n94, A2 => n92, B => n93, Z => n91);
   U214 : NAN2M1DL port map( A1 => n92, A2 => n93, Z => n13);
   U215 : INVDL port map( A => n84, Z => n82);
   U216 : NAN2M1DL port map( A1 => net12355, A2 => n70, Z => n9);
   U217 : INVD1 port map( A => net12354, Z => net12355);
   U218 : AOI21DL port map( A1 => net9993, A2 => n28, B => n29, Z => n27);
   U219 : EXNOR2DL port map( A1 => n27, A2 => net12169, Z => SUM(14));
   U220 : NAN2DL port map( A1 => n194, A2 => n52, Z => n195);
   U221 : NAN2D1 port map( A1 => n196, A2 => n195, Z => SUM(11));
   U222 : INVDL port map( A => n6, Z => n194);
   U223 : INVDL port map( A => n100, Z => n197);
   U224 : NAN2D1 port map( A1 => B(12), A2 => A(12), Z => n42);
   U225 : BUFDL port map( A => n179, Z => n198);
   U226 : INVDL port map( A => n82, Z => net11959);
   U227 : EXNOR2DL port map( A1 => n15, A2 => n103, Z => SUM(2));
   U228 : NAN2D2 port map( A1 => B(0), A2 => A(0), Z => n107);
   U229 : NAN2D1 port map( A1 => B(6), A2 => A(6), Z => n84);
   U230 : NOR2D2 port map( A1 => n55, A2 => n50, Z => n44);
   U231 : NAN2D2 port map( A1 => B(10), A2 => A(10), Z => n56);
   U232 : NOR2D2 port map( A1 => B(11), A2 => A(11), Z => n199);
   U233 : NAN2D1 port map( A1 => B(11), A2 => A(11), Z => n51);
   U234 : NOR2D2 port map( A1 => B(13), A2 => A(13), Z => n34);
   U235 : NAN2DL port map( A1 => n53, A2 => n56, Z => n7);
   U236 : INVDL port map( A => n55, Z => n53);
   U237 : INVDL port map( A => n56, Z => n54);
   U238 : NAN2DL port map( A1 => n197, A2 => n201, Z => n15);
   U239 : NAN2DL port map( A1 => B(2), A2 => A(2), Z => n102);
   U240 : AND2DL port map( A1 => n185, A2 => n107, Z => SUM(0));
   U241 : INVD1 port map( A => n102, Z => n100);
   U242 : NOR2D1 port map( A1 => B(6), A2 => A(6), Z => n83);
   U243 : NAN2D1 port map( A1 => B(3), A2 => A(3), Z => n97);
   U244 : NAN2DL port map( A1 => B(13), A2 => A(13), Z => n35);
   U245 : NOR2D1 port map( A1 => A(10), A2 => B(10), Z => n55);
   U246 : NAN2DL port map( A1 => B(5), A2 => A(5), Z => n90);
   U247 : NAN2D1 port map( A1 => B(7), A2 => A(7), Z => n79);
   U248 : OAI21DL port map( A1 => n75, A2 => net12355, B => n70, Z => n66);

end hier_sec_par_16_5;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_siso_gen.all;

architecture hier_sec_par_16_5 of siso_gen_DW_mult_tc_10 is

   component EXNOR2D4
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVDL
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AO21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22DL
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21M20DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN3D2
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D4
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR3D2
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22D2
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD16
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADFULD2
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component ADFULDL
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component BUFDL
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD20
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN3M1D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN3M1DL
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR3DL
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M20D2
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AO21M10DL
      port( A2, A1, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M10DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OA22DL
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component ADHALFD1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component AO21D2
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   signal n6, n9, n12, n16, n18, n22, n24, n28, n30, n34, n36, n40, n42, n46, 
      n48, n52, n53, n54, n55, n57, n60, n61, n62, n64, n69, n84, n85, n86, n87
      , n92, n93, n94, n95, n96, n97, n100, n101, n102, n103, n104, n105, n106,
      n107, n108, n109, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n125, n126, n127, n128, n129, n130, n133, n134, n135, n136, n139, n140, 
      n141, n142, n146, n147, n148, n149, n150, n151, n155, n157, n158, n159, 
      n160, n161, n162, n164, n167, n168, n169, n170, n171, n188, n189, n190, 
      n195, n202, n203, n204, n207, n208, n215, n216, n220, n267, n274, n275, 
      n276, n277, n287, n288, n289, n290, n293, n296, n297, n298, n299, n315, 
      n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, 
      n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, 
      n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, 
      n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, 
      n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, 
      n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, 
      n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, 
      n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, 
      n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, 
      n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, 
      n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, 
      n448, n449, n450, n453, n454, n457, n458, n459, n460, n462, n463, n467, 
      n471, n474, n476, n479, n480, n485, n486, n487, n488, n489, n490, n491, 
      n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, 
      n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, 
      n516, n517, n518, n519, n520, n521, n522, n523, n524, n526, n527, n528, 
      n529, n530, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, 
      n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, 
      n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, 
      n566, n567, n568, n569, n570, n571, n572, n573, n574, n577, n578, n579, 
      n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n592, 
      n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n606, 
      n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, 
      n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, 
      n631, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, 
      n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, 
      n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, 
      n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, 
      n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, 
      n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, 
      n705, n706, n707, n708, n710, n711, n712, n713, n714, n715, n716, n717, 
      n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, 
      n730, n731, n732, n733, n734, n735, n736, n738, n739, n740, n741, n742, 
      n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, 
      n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, 
      n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, 
      n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, 
      n792, n793, n794, n811, n812, n814, n834, n835, n842, net9957, net9959, 
      net10919, net10923, net11021, net11247, net11339, net11524, net11523, 
      net11686, net11792, net11944, net11943, net11942, net11946, net12005, 
      net12088, net12114, net12160, net12184, net12187, net12262, net12273, 
      net12315, net12321, net12350, net11920, n737, n206, n197, n196, n194, 
      n191, n187, n186, n300, n214, n213, n212, n211, net9976, net9975, net9974
      , net9972, net9971, net9969, net9968, net9967, net11982, net11981, 
      net11961, n469, n465, n456, n455, n452, n451, n221, n219, n218, n217, 
      net12148, net11941, n475, n468, net12274, n63, n295, n294, n199, n185, 
      n184, n183, n180, n179, n178, n176, n175, n174, net11996, n767, n632, 
      n604, n576, net12275, n484, n483, n269, n268, n266, n261, n250, n248, 
      n243, n235, n233, n231, n230, net11337, n709, n633, n605, n591, n525, 
      n482, n481, n478, n477, n472, n470, n466, net11803, net11797, net11020, 
      n473, n464, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, 
      n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, 
      n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, 
      n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, 
      n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, 
      n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, 
      n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, 
      n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, 
      n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, 
      n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, 
      n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, 
      n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, 
      n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
      n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
      n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, 
      n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, 
      n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
      n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, 
      n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, 
      n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, 
      n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, 
      n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, 
      n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, 
      n1153, n1154, n1155, n1156, n1157 : std_logic;

begin
   
   U54 : EXOR2D1 port map( A1 => n85, A2 => n54, Z => product(29));
   U59 : EXOR2D1 port map( A1 => n94, A2 => n55, Z => product(28));
   U78 : AOI21D1 port map( A1 => n120, A2 => n101, B => n102, Z => n100);
   U80 : OAI21D1 port map( A1 => n113, A2 => n103, B => n104, Z => n102);
   U108 : OAI21D1 port map( A1 => n133, A2 => n125, B => n126, Z => n120);
   U111 : NOR2D2 port map( A1 => n326, A2 => n331, Z => n125);
   U140 : AOI21D1 port map( A1 => net12273, A2 => n148, B => n149, Z => n147);
   U142 : OAI21D1 port map( A1 => n171, A2 => n150, B => n151, Z => n149);
   U154 : AOI21D1 port map( A1 => n159, A2 => net12273, B => n160, Z => n158);
   U156 : OAI21D1 port map( A1 => n171, A2 => n161, B => n162, Z => n160);
   U163 : NOR2D2 port map( A1 => n354, A2 => n363, Z => n161);
   U215 : NOR2D2 port map( A1 => n412, A2 => n425, Z => n202);
   U242 : NOR2D2 port map( A1 => net11792, A2 => n463, Z => n220);
   U324 : OAI21D1 port map( A1 => n275, A2 => n277, B => n276, Z => n274);
   U330 : AOI21D1 port map( A1 => n1150, A2 => n1152, B => n1151, Z => n277);
   U344 : ADFULD1 port map( A => n532, B => n319, CI => n547, CO => n315, S => 
                           n316);
   U345 : ADFULD1 port map( A => n320, B => n533, CI => n323, CO => n317, S => 
                           n318);
   U347 : ADFULD1 port map( A => n327, B => n534, CI => n324, CO => n321, S => 
                           n322);
   U348 : ADFULD1 port map( A => n548, B => n329, CI => n563, CO => n323, S => 
                           n324);
   U349 : ADFULD1 port map( A => n328, B => n335, CI => n333, CO => n325, S => 
                           n326);
   U350 : ADFULD1 port map( A => n535, B => n549, CI => n330, CO => n327, S => 
                           n328);
   U352 : ADFULD1 port map( A => n339, B => n336, CI => n334, CO => n331, S => 
                           n332);
   U353 : ADFULD1 port map( A => n343, B => n564, CI => n341, CO => n333, S => 
                           n334);
   U354 : ADFULD1 port map( A => n550, B => n536, CI => n579, CO => n335, S => 
                           n336);
   U355 : ADFULD1 port map( A => n347, B => n342, CI => n340, CO => n337, S => 
                           n338);
   U356 : ADFULD1 port map( A => n351, B => n344, CI => n349, CO => n339, S => 
                           n340);
   U357 : ADFULD1 port map( A => n537, B => n551, CI => n565, CO => n341, S => 
                           n342);
   U359 : ADFULD1 port map( A => n348, B => n357, CI => n355, CO => n345, S => 
                           n346);
   U360 : ADFULD1 port map( A => n350, B => n359, CI => n352, CO => n347, S => 
                           n348);
   U361 : ADFULD1 port map( A => n552, B => n361, CI => n566, CO => n349, S => 
                           n350);
   U362 : ADFULD1 port map( A => n580, B => n538, CI => n595, CO => n351, S => 
                           n352);
   U363 : ADFULD1 port map( A => n365, B => n358, CI => n356, CO => n353, S => 
                           n354);
   U364 : ADFULD1 port map( A => n360, B => n369, CI => n367, CO => n355, S => 
                           n356);
   U365 : ADFULD1 port map( A => n362, B => n567, CI => n371, CO => n357, S => 
                           n358);
   U366 : ADFULD1 port map( A => n581, B => n553, CI => n539, CO => n359, S => 
                           n360);
   U368 : ADFULD1 port map( A => n375, B => n368, CI => n366, CO => n363, S => 
                           n364);
   U369 : ADFULD1 port map( A => n372, B => n370, CI => n377, CO => n365, S => 
                           n366);
   U370 : ADFULD1 port map( A => n381, B => n582, CI => n379, CO => n367, S => 
                           n368);
   U371 : ADFULD1 port map( A => n554, B => n596, CI => n568, CO => n369, S => 
                           n370);
   U375 : ADFULD1 port map( A => n393, B => n395, CI => n382, CO => n377, S => 
                           n378);
   U376 : ADFULD1 port map( A => n541, B => n555, CI => n384, CO => n379, S => 
                           n380);
   U377 : ADFULD1 port map( A => n597, B => n569, CI => n583, CO => n381, S => 
                           n382);
   U380 : ADFULD1 port map( A => n392, B => n403, CI => n401, CO => n387, S => 
                           n388);
   U383 : ADFULD1 port map( A => n612, B => n556, CI => n598, CO => n393, S => 
                           n394);
   U384 : ADFULD1 port map( A => n409, B => n542, CI => n627, CO => n395, S => 
                           n396);
   U385 : ADFULD1 port map( A => n413, B => n402, CI => n400, CO => n397, S => 
                           n398);
   U386 : ADFULD1 port map( A => n404, B => n417, CI => n415, CO => n399, S => 
                           n400);
   U388 : ADFULD1 port map( A => n423, B => n410, CI => n421, CO => n403, S => 
                           n404);
   U390 : ADFULD1 port map( A => n613, B => n571, CI => n543, CO => n407, S => 
                           n408);
   U396 : ADFULD1 port map( A => n614, B => n628, CI => n572, CO => n419, S => 
                           n420);
   U399 : OR2D1 port map( A1 => n600, A2 => n558, Z => n423);
   U401 : ADFULD1 port map( A => n432, B => n436, CI => n443, CO => n427, S => 
                           n428);
   U403 : ADFULD1 port map( A => n438, B => n629, CI => n449, CO => n431, S => 
                           n432);
   U404 : ADFULD1 port map( A => n644, B => n587, CI => n615, CO => n433, S => 
                           n434);
   U405 : ADFULD1 port map( A => n545, B => n601, CI => n573, CO => n435, S => 
                           n436);
   U406 : ADHALFD1 port map( A => n559, B => n523, CO => n437, S => n438);
   U411 : ADFULD1 port map( A => n560, B => n630, CI => n588, CO => n447, S => 
                           n448);
   U414 : ADFULD1 port map( A => n458, B => n460, CI => n467, CO => n453, S => 
                           n454);
   U416 : ADFULD1 port map( A => n561, B => n617, CI => n589, CO => n457, S => 
                           n458);
   U430 : ADFULD1 port map( A => n495, B => n497, CI => n490, CO => n485, S => 
                           n486);
   U432 : ADFULD1 port map( A => n606, B => n578, CI => n649, CO => n489, S => 
                           n490);
   U433 : ADFULD1 port map( A => n496, B => n501, CI => n494, CO => n491, S => 
                           n492);
   U434 : ADFULD1 port map( A => n498, B => n650, CI => n503, CO => n493, S => 
                           n494);
   U436 : ADHALFD1 port map( A => n607, B => n526, CO => n497, S => n498);
   U437 : ADFULD1 port map( A => n504, B => n507, CI => n502, CO => n499, S => 
                           n500);
   U438 : ADFULD1 port map( A => n608, B => n636, CI => n509, CO => n501, S => 
                           n502);
   U439 : ADFULD1 port map( A => n622, B => n594, CI => n651, CO => n503, S => 
                           n504);
   U440 : ADFULD1 port map( A => n513, B => n510, CI => n508, CO => n505, S => 
                           n506);
   U441 : ADFULD1 port map( A => n609, B => n652, CI => n637, CO => n507, S => 
                           n508);
   U443 : ADFULD1 port map( A => n517, B => n624, CI => n514, CO => n511, S => 
                           n512);
   U444 : ADFULD1 port map( A => n653, B => n610, CI => n638, CO => n513, S => 
                           n514);
   U445 : ADFULD1 port map( A => n625, B => n639, CI => n518, CO => n515, S => 
                           n516);
   U446 : ADHALFD1 port map( A => n654, B => n528, CO => n517, S => n518);
   U447 : ADFULD1 port map( A => n655, B => n626, CI => n640, CO => n519, S => 
                           n520);
   U448 : ADHALFD1 port map( A => n656, B => n529, CO => n521, S => n522);
   U449 : OAI22D1 port map( A1 => n48, A2 => n835, B1 => n675, B2 => n46, Z => 
                           n523);
   U452 : OAI22D1 port map( A1 => n662, A2 => n48, B1 => n661, B2 => n46, Z => 
                           n533);
   U453 : OAI22D1 port map( A1 => n663, A2 => n48, B1 => n662, B2 => n46, Z => 
                           n534);
   U454 : OAI22D1 port map( A1 => n664, A2 => n48, B1 => n663, B2 => n46, Z => 
                           n535);
   U456 : OAI22D1 port map( A1 => n666, A2 => n48, B1 => n665, B2 => n46, Z => 
                           n537);
   U457 : OAI22D1 port map( A1 => n667, A2 => n48, B1 => n666, B2 => n46, Z => 
                           n538);
   U458 : OAI22D1 port map( A1 => n668, A2 => n48, B1 => n667, B2 => n46, Z => 
                           n539);
   U459 : OAI22D1 port map( A1 => n669, A2 => n48, B1 => n668, B2 => n46, Z => 
                           n540);
   U460 : OAI22D1 port map( A1 => n670, A2 => n48, B1 => n669, B2 => n46, Z => 
                           n541);
   U463 : OAI22D1 port map( A1 => n673, A2 => n48, B1 => n1057, B2 => n46, Z =>
                           n544);
   U465 : NOR2M1D1 port map( A1 => b(0), A2 => n46, Z => n546);
   U467 : EXNOR2D1 port map( A1 => b(14), A2 => a(15), Z => n660);
   U468 : EXNOR2D1 port map( A1 => b(13), A2 => a(15), Z => n661);
   U469 : EXNOR2D1 port map( A1 => b(12), A2 => a(15), Z => n662);
   U470 : EXNOR2D1 port map( A1 => b(11), A2 => a(15), Z => n663);
   U473 : EXNOR2D1 port map( A1 => b(8), A2 => a(15), Z => n666);
   U475 : EXNOR2D1 port map( A1 => b(6), A2 => a(15), Z => n668);
   U477 : EXNOR2D1 port map( A1 => b(4), A2 => a(15), Z => n670);
   U478 : EXNOR2D1 port map( A1 => b(3), A2 => a(15), Z => n671);
   U482 : NAN2M1D1 port map( A1 => b(0), A2 => a(15), Z => n675);
   U485 : OAI22D1 port map( A1 => n677, A2 => n42, B1 => n676, B2 => n40, Z => 
                           n319);
   U486 : OAI22D1 port map( A1 => n678, A2 => n42, B1 => n677, B2 => n40, Z => 
                           n548);
   U487 : OAI22D1 port map( A1 => n679, A2 => n42, B1 => n678, B2 => n40, Z => 
                           n549);
   U488 : OAI22D1 port map( A1 => n680, A2 => n42, B1 => n679, B2 => n40, Z => 
                           n550);
   U489 : OAI22D1 port map( A1 => n681, A2 => n42, B1 => n680, B2 => n40, Z => 
                           n551);
   U490 : OAI22D1 port map( A1 => n682, A2 => n42, B1 => n681, B2 => n40, Z => 
                           n552);
   U491 : OAI22D1 port map( A1 => n683, A2 => n42, B1 => n682, B2 => n40, Z => 
                           n553);
   U492 : OAI22D1 port map( A1 => n684, A2 => n42, B1 => n683, B2 => n40, Z => 
                           n554);
   U493 : OAI22D1 port map( A1 => n685, A2 => n42, B1 => n684, B2 => n40, Z => 
                           n555);
   U494 : OAI22D1 port map( A1 => n686, A2 => n42, B1 => n685, B2 => n40, Z => 
                           n556);
   U496 : OAI22D1 port map( A1 => n688, A2 => n42, B1 => n687, B2 => n40, Z => 
                           n558);
   U497 : OAI22D1 port map( A1 => n689, A2 => n42, B1 => n688, B2 => n40, Z => 
                           n559);
   U499 : OAI22D1 port map( A1 => n691, A2 => n42, B1 => n690, B2 => n40, Z => 
                           n561);
   U500 : NOR2M1D1 port map( A1 => b(0), A2 => n40, Z => n562);
   U501 : EXNOR2D1 port map( A1 => b(15), A2 => a(13), Z => n676);
   U502 : EXNOR2D1 port map( A1 => b(14), A2 => a(13), Z => n677);
   U503 : EXNOR2D1 port map( A1 => b(13), A2 => a(13), Z => n678);
   U504 : EXNOR2D1 port map( A1 => b(12), A2 => a(13), Z => n679);
   U505 : EXNOR2D1 port map( A1 => b(11), A2 => a(13), Z => n680);
   U506 : EXNOR2D1 port map( A1 => b(10), A2 => a(13), Z => n681);
   U507 : EXNOR2D1 port map( A1 => b(9), A2 => a(13), Z => n682);
   U508 : EXNOR2D1 port map( A1 => b(8), A2 => a(13), Z => n683);
   U510 : EXNOR2D1 port map( A1 => b(6), A2 => a(13), Z => n685);
   U512 : EXNOR2D1 port map( A1 => b(4), A2 => a(13), Z => n687);
   U514 : EXNOR2D1 port map( A1 => b(2), A2 => a(13), Z => n689);
   U520 : OAI22D1 port map( A1 => n694, A2 => n36, B1 => n693, B2 => n34, Z => 
                           n329);
   U521 : OAI22D1 port map( A1 => n695, A2 => n36, B1 => n694, B2 => n34, Z => 
                           n564);
   U522 : OAI22D1 port map( A1 => n696, A2 => n36, B1 => n695, B2 => n34, Z => 
                           n565);
   U523 : OAI22D1 port map( A1 => n697, A2 => n36, B1 => n696, B2 => n34, Z => 
                           n566);
   U525 : OAI22D1 port map( A1 => n699, A2 => n36, B1 => n698, B2 => n34, Z => 
                           n568);
   U526 : OAI22D1 port map( A1 => n700, A2 => n36, B1 => n699, B2 => n34, Z => 
                           n569);
   U529 : OAI22D1 port map( A1 => n703, A2 => n36, B1 => n702, B2 => n34, Z => 
                           n572);
   U535 : NOR2M1D1 port map( A1 => b(0), A2 => n34, Z => n578);
   U536 : EXNOR2D1 port map( A1 => b(15), A2 => a(11), Z => n693);
   U537 : EXNOR2D1 port map( A1 => b(14), A2 => a(11), Z => n694);
   U538 : EXNOR2D1 port map( A1 => b(13), A2 => a(11), Z => n695);
   U539 : EXNOR2D1 port map( A1 => b(12), A2 => a(11), Z => n696);
   U540 : EXNOR2D1 port map( A1 => b(11), A2 => a(11), Z => n697);
   U542 : EXNOR2D1 port map( A1 => b(9), A2 => a(11), Z => n699);
   U543 : EXNOR2D1 port map( A1 => b(8), A2 => a(11), Z => n700);
   U545 : EXNOR2D1 port map( A1 => b(6), A2 => a(11), Z => n702);
   U546 : EXNOR2D1 port map( A1 => b(5), A2 => a(11), Z => n703);
   U551 : EXNOR2D1 port map( A1 => b(0), A2 => a(11), Z => n708);
   U553 : OAI22D1 port map( A1 => n30, A2 => n1056, B1 => n726, B2 => n28, Z =>
                           n526);
   U555 : OAI22D1 port map( A1 => n711, A2 => n30, B1 => n710, B2 => n28, Z => 
                           n343);
   U556 : OAI22D1 port map( A1 => n712, A2 => n30, B1 => n711, B2 => n28, Z => 
                           n580);
   U557 : OAI22D1 port map( A1 => n713, A2 => n30, B1 => n712, B2 => n28, Z => 
                           n581);
   U558 : OAI22D1 port map( A1 => n714, A2 => n30, B1 => n713, B2 => n28, Z => 
                           n582);
   U559 : OAI22D1 port map( A1 => n715, A2 => n30, B1 => n714, B2 => n28, Z => 
                           n583);
   U562 : OAI22D1 port map( A1 => n718, A2 => n30, B1 => n717, B2 => n28, Z => 
                           n586);
   U565 : OAI22D1 port map( A1 => n1106, A2 => n30, B1 => n720, B2 => n28, Z =>
                           n589);
   U566 : OAI22D1 port map( A1 => n722, A2 => n30, B1 => n721, B2 => n28, Z => 
                           n590);
   U569 : OAI22D1 port map( A1 => n725, A2 => n30, B1 => n724, B2 => n28, Z => 
                           n593);
   U570 : NOR2M1D1 port map( A1 => b(0), A2 => n28, Z => n594);
   U571 : EXNOR2D1 port map( A1 => b(15), A2 => a(9), Z => n710);
   U572 : EXNOR2D1 port map( A1 => b(14), A2 => a(9), Z => n711);
   U573 : EXNOR2D1 port map( A1 => b(13), A2 => a(9), Z => n712);
   U574 : EXNOR2D1 port map( A1 => b(12), A2 => a(9), Z => n713);
   U575 : EXNOR2D1 port map( A1 => b(11), A2 => a(9), Z => n714);
   U576 : EXNOR2D1 port map( A1 => b(10), A2 => a(9), Z => n715);
   U586 : EXNOR2D1 port map( A1 => b(0), A2 => a(9), Z => n725);
   U587 : NAN2M1D1 port map( A1 => b(0), A2 => a(9), Z => n726);
   U588 : OAI22D1 port map( A1 => n24, A2 => net11920, B1 => n743, B2 => n22, Z
                           => n527);
   U590 : OAI22D1 port map( A1 => n728, A2 => n24, B1 => n727, B2 => n22, Z => 
                           n361);
   U591 : OAI22D1 port map( A1 => n729, A2 => n24, B1 => n728, B2 => n22, Z => 
                           n596);
   U592 : OAI22D1 port map( A1 => n730, A2 => n24, B1 => n729, B2 => n22, Z => 
                           n597);
   U593 : OAI22D1 port map( A1 => n731, A2 => n24, B1 => n730, B2 => n22, Z => 
                           n598);
   U594 : OAI22D1 port map( A1 => n732, A2 => n24, B1 => n731, B2 => n22, Z => 
                           n599);
   U595 : OAI22D1 port map( A1 => n733, A2 => n24, B1 => n732, B2 => n22, Z => 
                           n600);
   U596 : OAI22D1 port map( A1 => n734, A2 => n24, B1 => n733, B2 => n22, Z => 
                           n601);
   U597 : OAI22D1 port map( A1 => n735, A2 => n24, B1 => n734, B2 => n22, Z => 
                           n602);
   U598 : OAI22D1 port map( A1 => n736, A2 => n24, B1 => n735, B2 => n22, Z => 
                           n603);
   U601 : OAI22D1 port map( A1 => n739, A2 => n24, B1 => n738, B2 => n22, Z => 
                           n606);
   U603 : OAI22D1 port map( A1 => n741, A2 => n24, B1 => n740, B2 => n22, Z => 
                           n608);
   U604 : OAI22D1 port map( A1 => n742, A2 => n24, B1 => n741, B2 => n22, Z => 
                           n609);
   U605 : NOR2M1D1 port map( A1 => b(0), A2 => n22, Z => n610);
   U606 : EXNOR2D1 port map( A1 => b(15), A2 => a(7), Z => n727);
   U607 : EXNOR2D1 port map( A1 => b(14), A2 => a(7), Z => n728);
   U608 : EXNOR2D1 port map( A1 => b(13), A2 => a(7), Z => n729);
   U609 : EXNOR2D1 port map( A1 => b(12), A2 => a(7), Z => n730);
   U610 : EXNOR2D1 port map( A1 => b(11), A2 => a(7), Z => n731);
   U613 : EXNOR2D1 port map( A1 => b(8), A2 => a(7), Z => n734);
   U617 : EXNOR2D1 port map( A1 => b(4), A2 => a(7), Z => n738);
   U618 : EXNOR2D1 port map( A1 => b(3), A2 => a(7), Z => n739);
   U619 : EXNOR2D1 port map( A1 => b(2), A2 => a(7), Z => n740);
   U620 : EXNOR2D1 port map( A1 => b(1), A2 => a(7), Z => n741);
   U621 : EXNOR2D1 port map( A1 => b(0), A2 => a(7), Z => n742);
   U622 : NAN2M1D1 port map( A1 => b(0), A2 => a(7), Z => n743);
   U623 : OAI22D1 port map( A1 => n18, A2 => net12088, B1 => n760, B2 => n16, Z
                           => n528);
   U625 : OAI22D1 port map( A1 => n745, A2 => n18, B1 => n744, B2 => n16, Z => 
                           n383);
   U626 : OAI22D1 port map( A1 => n746, A2 => n18, B1 => n745, B2 => n16, Z => 
                           n612);
   U627 : OAI22D1 port map( A1 => n747, A2 => n18, B1 => n746, B2 => n16, Z => 
                           n613);
   U628 : OAI22D1 port map( A1 => n748, A2 => n18, B1 => n747, B2 => n16, Z => 
                           n614);
   U629 : OAI22D1 port map( A1 => n749, A2 => n18, B1 => n1090, B2 => n16, Z =>
                           n615);
   U631 : OAI22D1 port map( A1 => n751, A2 => n18, B1 => n750, B2 => n16, Z => 
                           n617);
   U635 : OAI22D1 port map( A1 => n755, A2 => n18, B1 => n754, B2 => n16, Z => 
                           n621);
   U636 : OAI22D1 port map( A1 => n756, A2 => n18, B1 => n755, B2 => n16, Z => 
                           n622);
   U637 : OAI22D1 port map( A1 => n757, A2 => n18, B1 => n756, B2 => n16, Z => 
                           n623);
   U639 : OAI22D1 port map( A1 => n759, A2 => n18, B1 => n758, B2 => n16, Z => 
                           n625);
   U640 : NOR2M1D1 port map( A1 => b(0), A2 => n16, Z => n626);
   U641 : EXNOR2D1 port map( A1 => b(15), A2 => a(5), Z => n744);
   U642 : EXNOR2D1 port map( A1 => b(14), A2 => a(5), Z => n745);
   U643 : EXNOR2D1 port map( A1 => b(13), A2 => a(5), Z => n746);
   U653 : EXNOR2D1 port map( A1 => b(3), A2 => a(5), Z => n756);
   U656 : EXNOR2D1 port map( A1 => b(0), A2 => a(5), Z => n759);
   U657 : NAN2M1D1 port map( A1 => b(0), A2 => a(5), Z => n760);
   U658 : OAI22D1 port map( A1 => n12, A2 => net12160, B1 => n777, B2 => n9, Z 
                           => n529);
   U660 : OAI22D1 port map( A1 => n762, A2 => n12, B1 => n761, B2 => n9, Z => 
                           n409);
   U661 : OAI22D1 port map( A1 => n763, A2 => n12, B1 => n762, B2 => n9, Z => 
                           n628);
   U664 : OAI22D1 port map( A1 => n766, A2 => n12, B1 => n765, B2 => n9, Z => 
                           n631);
   U667 : OAI22D1 port map( A1 => n769, A2 => n12, B1 => n768, B2 => n9, Z => 
                           n634);
   U668 : OAI22D1 port map( A1 => n770, A2 => n12, B1 => n769, B2 => n9, Z => 
                           n635);
   U669 : OAI22D1 port map( A1 => n771, A2 => n12, B1 => n770, B2 => n9, Z => 
                           n636);
   U670 : OAI22D1 port map( A1 => n772, A2 => n12, B1 => n771, B2 => n9, Z => 
                           n637);
   U671 : OAI22D1 port map( A1 => n773, A2 => n12, B1 => n772, B2 => n9, Z => 
                           n638);
   U672 : OAI22D1 port map( A1 => n774, A2 => n12, B1 => n773, B2 => n9, Z => 
                           n639);
   U673 : OAI22D1 port map( A1 => n775, A2 => n12, B1 => n774, B2 => n9, Z => 
                           n640);
   U674 : OAI22D1 port map( A1 => n776, A2 => n12, B1 => n775, B2 => n9, Z => 
                           n641);
   U675 : NOR2M1D1 port map( A1 => b(0), A2 => n9, Z => n642);
   U676 : EXNOR2D1 port map( A1 => b(15), A2 => a(3), Z => n761);
   U679 : EXNOR2D1 port map( A1 => b(12), A2 => a(3), Z => n764);
   U683 : EXNOR2D1 port map( A1 => b(8), A2 => a(3), Z => n768);
   U685 : EXNOR2D1 port map( A1 => b(6), A2 => a(3), Z => n770);
   U686 : EXNOR2D1 port map( A1 => b(5), A2 => a(3), Z => n771);
   U687 : EXNOR2D1 port map( A1 => b(4), A2 => a(3), Z => n772);
   U688 : EXNOR2D1 port map( A1 => b(3), A2 => a(3), Z => n773);
   U689 : EXNOR2D1 port map( A1 => b(2), A2 => a(3), Z => n774);
   U690 : EXNOR2D1 port map( A1 => b(1), A2 => a(3), Z => n775);
   U691 : EXNOR2D1 port map( A1 => b(0), A2 => a(3), Z => n776);
   U692 : NAN2M1D1 port map( A1 => b(0), A2 => a(3), Z => n777);
   U693 : OAI22D1 port map( A1 => n6, A2 => n842, B1 => n794, B2 => n834, Z => 
                           n530);
   U694 : AO21D2 port map( A1 => n6, A2 => n834, B => n778, Z => n643);
   U695 : OAI22D1 port map( A1 => n779, A2 => n6, B1 => n931, B2 => n834, Z => 
                           n644);
   U696 : OAI22D1 port map( A1 => n780, A2 => n6, B1 => n1082, B2 => n834, Z =>
                           n645);
   U698 : OAI22D1 port map( A1 => n1107, A2 => n6, B1 => n781, B2 => n834, Z =>
                           n647);
   U699 : OAI22D1 port map( A1 => n783, A2 => n6, B1 => n782, B2 => n834, Z => 
                           n648);
   U702 : OAI22D1 port map( A1 => n786, A2 => n6, B1 => n785, B2 => n834, Z => 
                           n651);
   U703 : OAI22D1 port map( A1 => n787, A2 => n6, B1 => n786, B2 => n834, Z => 
                           n652);
   U704 : OAI22D1 port map( A1 => n788, A2 => n6, B1 => n787, B2 => n834, Z => 
                           n653);
   U706 : OAI22D1 port map( A1 => n790, A2 => n6, B1 => n789, B2 => n834, Z => 
                           n655);
   U708 : OAI22D1 port map( A1 => n792, A2 => n6, B1 => n791, B2 => n834, Z => 
                           n657);
   U711 : EXNOR2D1 port map( A1 => b(15), A2 => a(1), Z => n778);
   U713 : EXNOR2D1 port map( A1 => b(13), A2 => a(1), Z => n780);
   U718 : EXNOR2D1 port map( A1 => b(8), A2 => a(1), Z => n785);
   U720 : EXNOR2D1 port map( A1 => b(6), A2 => a(1), Z => n787);
   U721 : EXNOR2D1 port map( A1 => b(5), A2 => a(1), Z => n788);
   U722 : EXNOR2D1 port map( A1 => b(4), A2 => a(1), Z => n789);
   U723 : EXNOR2D1 port map( A1 => b(3), A2 => a(1), Z => n790);
   U724 : EXNOR2D1 port map( A1 => b(2), A2 => a(1), Z => n791);
   U725 : EXNOR2D1 port map( A1 => b(1), A2 => a(1), Z => n792);
   U726 : EXNOR2D1 port map( A1 => b(0), A2 => a(1), Z => n793);
   U727 : NAN2M1D1 port map( A1 => b(0), A2 => a(1), Z => n794);
   U752 : EXOR2D1 port map( A1 => a(14), A2 => a(15), Z => n811);
   U755 : EXOR2D1 port map( A1 => a(13), A2 => a(12), Z => n812);
   U761 : EXOR2D1 port map( A1 => a(9), A2 => a(8), Z => n814);
   U203 : NOR2D2 port map( A1 => n398, A2 => n411, Z => n191);
   U212 : OAI21D1 port map( A1 => n208, A2 => n202, B => n203, Z => n197);
   U415 : ADFULD1 port map( A => n462, B => n471, CI => n469, CO => n455, S => 
                           n456);
   U232 : NOR2D2 port map( A1 => n440, A2 => n451, Z => n213);
   U188 : AOI21D1 port map( A1 => n197, A2 => n1033, B => n185, Z => n183);
   U172 : OAI21D1 port map( A1 => n174, A2 => n180, B => n175, Z => n169);
   U534 : OAI22D1 port map( A1 => n708, A2 => n36, B1 => n707, B2 => n34, Z => 
                           n577);
   U665 : OAI22D1 port map( A1 => n767, A2 => n12, B1 => n1030, B2 => n9, Z => 
                           n632);
   U316 : AOI21D1 port map( A1 => net10919, A2 => n274, B => n1018, Z => n269);
   U310 : OAI21D1 port map( A1 => n267, A2 => n269, B => n268, Z => n266);
   U302 : AOI21D1 port map( A1 => net10923, A2 => n266, B => n1019, Z => n261);
   U285 : AOI21D1 port map( A1 => net11021, A2 => n1024, B => n1022, Z => n250)
                           ;
   U275 : AOI21D1 port map( A1 => n248, A2 => n1021, B => n1020, Z => n243);
   U263 : NOR2D2 port map( A1 => n474, A2 => n483, Z => n235);
   U429 : ADFULD1 port map( A => n493, B => n488, CI => n486, CO => n483, S => 
                           n484);
   U218 : AOI21D1 port map( A1 => n299, A2 => net12275, B => n206, Z => n204);
   U552 : NAN2M1D1 port map( A1 => b(0), A2 => a(11), Z => n709);
   U518 : OAI22D1 port map( A1 => n36, A2 => net11946, B1 => n709, B2 => n34, Z
                           => n525);
   U428 : ADHALFD1 port map( A => n525, B => n591, CO => n481, S => n482);
   U426 : ADFULD1 port map( A => n605, B => n633, CI => n482, CO => n477, S => 
                           n478);
   U599 : OAI22D1 port map( A1 => n737, A2 => n24, B1 => n1016, B2 => n22, Z =>
                           n604);
   U237 : AOI21D1 port map( A1 => n218, A2 => net12350, B => n219, Z => n217);
   U777 : INVDL port map( A => n485, Z => n910);
   U778 : INVDL port map( A => n910, Z => n911);
   U779 : NAN2DL port map( A1 => n472, A2 => n477, Z => net9969);
   U780 : EXOR3D2 port map( A1 => n437, A2 => n424, A3 => n435, Z => n418);
   U781 : NAN2D1 port map( A1 => n427, A2 => n416, Z => n914);
   U782 : NAN2D2 port map( A1 => n912, A2 => n913, Z => n915);
   U783 : NAN2D2 port map( A1 => n914, A2 => n915, Z => n1081);
   U784 : INVD1 port map( A => n427, Z => n912);
   U785 : INVDL port map( A => n416, Z => n913);
   U786 : EXOR3D2 port map( A1 => n433, A2 => n422, A3 => n420, Z => n416);
   U787 : EXOR3D2 port map( A1 => n465, A2 => n456, A3 => n454, Z => net11792);
   U788 : NAN2D2 port map( A1 => n1073, A2 => n1074, Z => n751);
   U789 : EXNOR2DL port map( A1 => b(6), A2 => a(7), Z => n916);
   U790 : EXNOR2D1 port map( A1 => b(2), A2 => a(9), Z => n917);
   U791 : NAN2D1 port map( A1 => n424, A2 => n435, Z => n1048);
   U792 : NAN2D1 port map( A1 => b(3), A2 => a(13), Z => n920);
   U793 : NAN2D2 port map( A1 => n918, A2 => n919, Z => n921);
   U794 : NAN2D2 port map( A1 => n920, A2 => n921, Z => n688);
   U795 : INVD2 port map( A => b(3), Z => n918);
   U796 : INVDL port map( A => a(13), Z => n919);
   U797 : EXNOR2D1 port map( A1 => b(10), A2 => a(3), Z => n1030);
   U798 : NAN2D1 port map( A1 => n1113, A2 => n923, Z => n924);
   U799 : NAN2D1 port map( A1 => n922, A2 => n428, Z => n925);
   U800 : NAN2D2 port map( A1 => n924, A2 => n925, Z => n426);
   U801 : INVD2 port map( A => n1113, Z => n922);
   U802 : INVDL port map( A => n428, Z => n923);
   U803 : NAN2D1 port map( A1 => n426, A2 => n439, Z => n954);
   U804 : NOR2D1 port map( A1 => n426, A2 => n439, Z => n207);
   U805 : INVD1 port map( A => n199, Z => n926);
   U806 : INVD1 port map( A => n197, Z => n199);
   U807 : NAN2DL port map( A1 => b(6), A2 => a(7), Z => n929);
   U808 : NAN2D1 port map( A1 => n927, A2 => n928, Z => n930);
   U809 : NAN2D1 port map( A1 => n929, A2 => n930, Z => n1016);
   U810 : INVD1 port map( A => b(6), Z => n927);
   U811 : INVDL port map( A => a(7), Z => n928);
   U812 : INVD1 port map( A => n221, Z => n219);
   U813 : EXNOR2DL port map( A1 => b(15), A2 => a(1), Z => n931);
   U814 : AND2D1 port map( A1 => n464, A2 => n473, Z => net12350);
   U815 : AOI21D1 port map( A1 => n169, A2 => n139, B => n140, Z => n1064);
   U816 : INVDL port map( A => net12187, Z => n1002);
   U817 : EXOR3D1 port map( A1 => n399, A2 => n390, A3 => n388, Z => n386);
   U818 : NAN2DL port map( A1 => n399, A2 => n388, Z => n932);
   U819 : NAN2DL port map( A1 => n399, A2 => n390, Z => n933);
   U820 : NAN2DL port map( A1 => n388, A2 => n390, Z => n934);
   U821 : NAN3D1 port map( A1 => n932, A2 => n934, A3 => n933, Z => n385);
   U822 : EXOR3D1 port map( A1 => n405, A2 => n394, A3 => n396, Z => n390);
   U823 : NOR2D1 port map( A1 => n386, A2 => n397, Z => n186);
   U824 : INVD2 port map( A => n430, Z => n1077);
   U825 : OAI21D1 port map( A1 => n141, A2 => n162, B => n142, Z => n140);
   U826 : INVD2 port map( A => b(9), Z => net11996);
   U827 : NAN2D1 port map( A1 => b(10), A2 => n1075, Z => n937);
   U828 : NAN2D1 port map( A1 => n935, A2 => n936, Z => n938);
   U829 : NAN2D1 port map( A1 => n937, A2 => n938, Z => n783);
   U830 : INVD1 port map( A => b(10), Z => n935);
   U831 : INVD1 port map( A => n1075, Z => n936);
   U832 : EXNOR2DL port map( A1 => b(10), A2 => a(15), Z => n664);
   U833 : EXNOR2DL port map( A1 => b(10), A2 => a(5), Z => n749);
   U834 : INVD16 port map( A => b(10), Z => n986);
   U835 : NAN2D2 port map( A1 => n1078, A2 => n1079, Z => n1113);
   U836 : NOR2DL port map( A1 => n170, A2 => n161, Z => n159);
   U837 : INVDL port map( A => n125, Z => n289);
   U838 : EXOR2D1 port map( A1 => n57, A2 => n114, Z => product(26));
   U839 : NAN2DL port map( A1 => b(11), A2 => a(5), Z => n994);
   U840 : INVD1 port map( A => n842, Z => n1075);
   U841 : OR2D1 port map( A1 => n752, A2 => n16, Z => n1141);
   U842 : NAN2D1 port map( A1 => n1087, A2 => n1088, Z => n752);
   U843 : INVD16 port map( A => b(3), Z => n1110);
   U844 : NAN3D1 port map( A1 => n1096, A2 => n1098, A3 => n1097, Z => n405);
   U845 : INVD1 port map( A => a(0), Z => n834);
   U846 : OAI22D1 port map( A1 => n1108, A2 => n18, B1 => n1105, B2 => n16, Z 
                           => n618);
   U847 : OAI22DL port map( A1 => n754, A2 => n18, B1 => n1104, B2 => n16, Z =>
                           n620);
   U848 : NOR2D1 port map( A1 => n332, A2 => n337, Z => n130);
   U849 : NAN2DL port map( A1 => n294, A2 => n175, Z => n63);
   U850 : INVD1 port map( A => a(5), Z => net12088);
   U851 : INVD1 port map( A => a(9), Z => n1056);
   U852 : INVDL port map( A => a(11), Z => net11946);
   U853 : INVDL port map( A => a(3), Z => net12160);
   U854 : AND2D1 port map( A1 => n943, A2 => n524, Z => n939);
   U855 : AND2DL port map( A1 => n911, A2 => n478, Z => n940);
   U856 : AND2DL port map( A1 => n290, A2 => n133, Z => n941);
   U857 : OA22DL port map( A1 => n660, A2 => n48, B1 => n659, B2 => n46, Z => 
                           n942);
   U858 : EXNOR2D1 port map( A1 => b(12), A2 => a(1), Z => n781);
   U859 : EXOR2D1 port map( A1 => n623, A2 => n527, Z => n510);
   U860 : OAI22D1 port map( A1 => n706, A2 => n36, B1 => n1080, B2 => n34, Z =>
                           n943);
   U861 : EXNOR2D1 port map( A1 => b(8), A2 => a(9), Z => n1092);
   U862 : OAI22DL port map( A1 => n704, A2 => n36, B1 => n703, B2 => n34, Z => 
                           n573);
   U863 : EXNOR2D1 port map( A1 => b(4), A2 => a(11), Z => n704);
   U864 : EXOR2D1 port map( A1 => n947, A2 => n450, Z => n444);
   U865 : NAN2D2 port map( A1 => n1072, A2 => net12088, Z => n1074);
   U866 : NAN2DL port map( A1 => n422, A2 => n420, Z => n944);
   U867 : NAN2DL port map( A1 => n422, A2 => n433, Z => n945);
   U868 : NAN2D1 port map( A1 => n420, A2 => n433, Z => n946);
   U869 : NAN3D1 port map( A1 => n944, A2 => n946, A3 => n945, Z => n415);
   U870 : EXOR3D1 port map( A1 => n643, A2 => n544, A3 => n586, Z => n422);
   U871 : EXOR3D2 port map( A1 => n574, A2 => n546, A3 => n645, Z => n450);
   U872 : EXOR2D1 port map( A1 => n457, A2 => n459, Z => n947);
   U873 : NAN2D1 port map( A1 => n574, A2 => n546, Z => n948);
   U874 : NAN2D1 port map( A1 => n574, A2 => n645, Z => n949);
   U875 : NAN2D1 port map( A1 => n546, A2 => n645, Z => n950);
   U876 : NAN3D2 port map( A1 => n948, A2 => n949, A3 => n950, Z => n449);
   U877 : NAN2DL port map( A1 => n457, A2 => n459, Z => n951);
   U878 : NAN2D1 port map( A1 => n457, A2 => n450, Z => n952);
   U879 : NAN2D1 port map( A1 => n459, A2 => n450, Z => n953);
   U880 : NAN3D2 port map( A1 => n951, A2 => n952, A3 => n953, Z => n443);
   U881 : NAN2D1 port map( A1 => n1043, A2 => n1044, Z => n737);
   U882 : NAN2DL port map( A1 => n426, A2 => n439, Z => n208);
   U883 : INVDL port map( A => n999, Z => n1028);
   U884 : INVD2 port map( A => n1001, Z => n509);
   U885 : NOR2DL port map( A1 => n202, A2 => n207, Z => n955);
   U886 : NOR2DL port map( A1 => n202, A2 => n207, Z => n956);
   U887 : NOR2DL port map( A1 => n202, A2 => n207, Z => n196);
   U888 : NAN2D1 port map( A1 => b(1), A2 => a(13), Z => n958);
   U889 : NAN2D2 port map( A1 => n957, A2 => n1061, Z => n959);
   U890 : NAN2D2 port map( A1 => n958, A2 => n959, Z => n690);
   U891 : INVD4 port map( A => b(1), Z => n957);
   U892 : NAN2D2 port map( A1 => n1067, A2 => net12160, Z => n1068);
   U893 : NAN2D2 port map( A1 => n1111, A2 => n1112, Z => n722);
   U894 : OAI22D1 port map( A1 => n672, A2 => n48, B1 => n671, B2 => n46, Z => 
                           n543);
   U895 : EXNOR2DL port map( A1 => b(2), A2 => a(15), Z => n672);
   U896 : NAN2D1 port map( A1 => b(11), A2 => a(3), Z => n960);
   U897 : NAN2D2 port map( A1 => n993, A2 => net12160, Z => n961);
   U898 : NAN2D2 port map( A1 => n960, A2 => n961, Z => n765);
   U899 : OAI22DL port map( A1 => n765, A2 => n12, B1 => n764, B2 => n9, Z => 
                           n630);
   U900 : NAN2D1 port map( A1 => b(9), A2 => a(9), Z => n963);
   U901 : NAN2D2 port map( A1 => n962, A2 => n1056, Z => n964);
   U902 : NAN2D1 port map( A1 => n963, A2 => n964, Z => n716);
   U903 : INVD2 port map( A => b(9), Z => n962);
   U904 : OAI22D1 port map( A1 => n716, A2 => n30, B1 => n715, B2 => n28, Z => 
                           n584);
   U905 : NAN3D2 port map( A1 => n1048, A2 => n1050, A3 => n1049, Z => n417);
   U906 : NAN2D1 port map( A1 => n374, A2 => n385, Z => n180);
   U907 : NAN2D2 port map( A1 => n993, A2 => net12088, Z => n995);
   U908 : INVD20 port map( A => b(11), Z => n993);
   U909 : NAN2D1 port map( A1 => n1081, A2 => n414, Z => n967);
   U910 : NAN2D2 port map( A1 => n965, A2 => n966, Z => n968);
   U911 : NAN2D2 port map( A1 => n967, A2 => n968, Z => n412);
   U912 : INVD2 port map( A => n1081, Z => n965);
   U913 : INVD2 port map( A => n414, Z => n966);
   U914 : NAN2D1 port map( A1 => n429, A2 => n431, Z => n1120);
   U915 : NAN2D1 port map( A1 => n394, A2 => n396, Z => n969);
   U916 : NAN2D1 port map( A1 => n394, A2 => n405, Z => n970);
   U917 : NAN2D1 port map( A1 => n396, A2 => n405, Z => n971);
   U918 : NAN3D2 port map( A1 => n969, A2 => n971, A3 => n970, Z => n389);
   U919 : EXOR3D1 port map( A1 => n391, A2 => n380, A3 => n389, Z => n376);
   U920 : EXOR2D2 port map( A1 => n387, A2 => n378, Z => n972);
   U921 : EXOR2D1 port map( A1 => n972, A2 => n376, Z => n374);
   U922 : NAN2DL port map( A1 => n391, A2 => n380, Z => n973);
   U923 : NAN2D1 port map( A1 => n391, A2 => n389, Z => n974);
   U924 : NAN2D1 port map( A1 => n380, A2 => n389, Z => n975);
   U925 : NAN3D2 port map( A1 => n973, A2 => n974, A3 => n975, Z => n375);
   U926 : NAN2DL port map( A1 => n387, A2 => n378, Z => n976);
   U927 : NAN2DL port map( A1 => n387, A2 => n376, Z => n977);
   U928 : NAN2DL port map( A1 => n378, A2 => n376, Z => n978);
   U929 : NAN3D1 port map( A1 => n976, A2 => n977, A3 => n978, Z => n373);
   U930 : INVD16 port map( A => b(5), Z => n1042);
   U931 : INVDL port map( A => n604, Z => net11981);
   U932 : EXNOR2DL port map( A1 => b(9), A2 => a(5), Z => n979);
   U933 : NAN2D1 port map( A1 => n994, A2 => n995, Z => n748);
   U934 : AND2D1 port map( A1 => n297, A2 => n1010, Z => net9957);
   U935 : NAN2D1 port map( A1 => b(12), A2 => a(5), Z => n981);
   U936 : NAN2D2 port map( A1 => n980, A2 => net12088, Z => n982);
   U937 : NAN2D2 port map( A1 => n981, A2 => n982, Z => n747);
   U938 : INVD2 port map( A => b(12), Z => n980);
   U939 : EXOR3D1 port map( A1 => n602, A2 => n616, A3 => n939, Z => n446);
   U940 : NAN2DL port map( A1 => n616, A2 => n939, Z => n983);
   U941 : NAN2DL port map( A1 => n616, A2 => n602, Z => n984);
   U942 : NAN2D1 port map( A1 => n939, A2 => n602, Z => n985);
   U943 : NAN3D1 port map( A1 => n983, A2 => n985, A3 => n984, Z => n445);
   U944 : OAI22D1 port map( A1 => n28, A2 => n718, B1 => n719, B2 => n30, Z => 
                           n587);
   U945 : NAN2D1 port map( A1 => b(10), A2 => a(7), Z => n987);
   U946 : NAN2D2 port map( A1 => n986, A2 => net11920, Z => n988);
   U947 : NAN2D2 port map( A1 => n987, A2 => n988, Z => n732);
   U948 : EXNOR2D2 port map( A1 => n989, A2 => n442, Z => n440);
   U949 : EXNOR2D1 port map( A1 => n453, A2 => n444, Z => n989);
   U950 : EXNOR2D2 port map( A1 => b(6), A2 => a(9), Z => n719);
   U951 : OAI21DL port map( A1 => n52, A2 => n130, B => n133, Z => n129);
   U952 : EXOR2D1 port map( A1 => n485, A2 => n478, Z => net11797);
   U953 : NAN2DL port map( A1 => n544, A2 => n586, Z => n990);
   U954 : NAN2DL port map( A1 => n544, A2 => n643, Z => n991);
   U955 : NAN2DL port map( A1 => n586, A2 => n643, Z => n992);
   U956 : NAN3D1 port map( A1 => n992, A2 => n990, A3 => n991, Z => n421);
   U957 : OAI22DL port map( A1 => n979, A2 => n18, B1 => n749, B2 => n16, Z => 
                           n616);
   U958 : EXNOR2D1 port map( A1 => b(2), A2 => a(15), Z => n1057);
   U959 : NAN2DL port map( A1 => n428, A2 => n441, Z => n1115);
   U960 : NAN3D2 port map( A1 => n1123, A2 => n1124, A3 => n1125, Z => n411);
   U961 : OAI22DL port map( A1 => n42, A2 => n1061, B1 => n692, B2 => n40, Z =>
                           n524);
   U962 : EXOR3D2 port map( A1 => n429, A2 => n431, A3 => n418, Z => n414);
   U963 : OAI21D1 port map( A1 => n1067, A2 => net12160, B => n1068, Z => n763)
                           ;
   U964 : INVD20 port map( A => b(13), Z => n1067);
   U965 : OAI22D1 port map( A1 => n716, A2 => n28, B1 => n30, B2 => n1092, Z =>
                           n585);
   U966 : OAI21M20D2 port map( A1 => n230, A2 => n211, B => n996, Z => net12275
                           );
   U967 : INVD1 port map( A => n212, Z => n996);
   U968 : EXOR3D1 port map( A1 => n599, A2 => n585, A3 => n557, Z => n406);
   U969 : OAI21M20D1 port map( A1 => n997, A2 => n998, B => n218, Z => n216);
   U970 : INVDL port map( A => n464, Z => n997);
   U971 : INVDL port map( A => n473, Z => n998);
   U972 : OAI22D1 port map( A1 => n36, A2 => n705, B1 => n704, B2 => n34, Z => 
                           n574);
   U973 : OAI21D1 port map( A1 => n235, A2 => n1025, B => n1027, Z => n999);
   U974 : OAI21M10DL port map( A1 => n119, A2 => n52, B => n118, Z => n116);
   U975 : NAN2M1D1 port map( A1 => n1000, A2 => n623, Z => n1001);
   U976 : INVDL port map( A => n527, Z => n1000);
   U977 : NAN3M1D1 port map( A1 => n940, A2 => n1015, A3 => net11803, Z => n473
                           );
   U978 : AO21M10DL port map( A2 => n230, A1 => n216, B => n1002, Z => n215);
   U979 : EXNOR2D1 port map( A1 => b(2), A2 => a(9), Z => n723);
   U980 : NAN2D1 port map( A1 => b(7), A2 => a(11), Z => n1004);
   U981 : NAN2D2 port map( A1 => n1003, A2 => net11946, Z => n1005);
   U982 : NAN2D2 port map( A1 => n1004, A2 => n1005, Z => n701);
   U983 : INVD4 port map( A => b(7), Z => n1003);
   U984 : NOR2DL port map( A1 => n397, A2 => n386, Z => n1006);
   U985 : OAI22D1 port map( A1 => n701, A2 => n36, B1 => n700, B2 => n34, Z => 
                           n570);
   U986 : NAN2DL port map( A1 => b(6), A2 => a(5), Z => n1008);
   U987 : NAN2D1 port map( A1 => n1007, A2 => net12088, Z => n1009);
   U988 : NAN2D1 port map( A1 => n1008, A2 => n1009, Z => n753);
   U989 : INVD2 port map( A => b(6), Z => n1007);
   U990 : OR2D1 port map( A1 => n753, A2 => n18, Z => n1140);
   U991 : INVD2 port map( A => n220, Z => n218);
   U992 : NAN2DL port map( A1 => n1038, A2 => n411, Z => n1010);
   U993 : NAN2DL port map( A1 => n1038, A2 => n411, Z => n194);
   U994 : NAN2D2 port map( A1 => n1042, A2 => net11920, Z => n1044);
   U995 : NAN2DL port map( A1 => net11020, A2 => n466, Z => n1013);
   U996 : NAN2D1 port map( A1 => n1011, A2 => n1012, Z => n1014);
   U997 : NAN2D1 port map( A1 => n1013, A2 => n1014, Z => n464);
   U998 : INVD1 port map( A => net11020, Z => n1011);
   U999 : INVDL port map( A => n466, Z => n1012);
   U1000 : EXOR3D1 port map( A1 => n470, A2 => n472, A3 => n477, Z => n466);
   U1001 : EXNOR2D1 port map( A1 => n468, A2 => n475, Z => net11020);
   U1002 : NAN2DL port map( A1 => n478, A2 => n476, Z => net11803);
   U1003 : NAN2DL port map( A1 => n476, A2 => n911, Z => n1015);
   U1004 : NAN2DL port map( A1 => n468, A2 => n466, Z => net9971);
   U1005 : NAN2DL port map( A1 => n475, A2 => n466, Z => net9972);
   U1006 : AND2DL port map( A1 => n468, A2 => n475, Z => net11961);
   U1007 : EXOR2D1 port map( A1 => net11797, A2 => n476, Z => n474);
   U1008 : EXOR2D2 port map( A1 => net11337, A2 => n576, Z => n470);
   U1009 : NAN2DL port map( A1 => n470, A2 => n472, Z => net9967);
   U1010 : NAN2DL port map( A1 => n477, A2 => n470, Z => net9968);
   U1011 : EXOR2D1 port map( A1 => n632, A2 => n604, Z => net11337);
   U1012 : EXOR3D1 port map( A1 => n562, A2 => n590, A3 => n647, Z => n472);
   U1013 : NAN2D1 port map( A1 => n479, A2 => n481, Z => net11942);
   U1014 : NAN2DL port map( A1 => n481, A2 => n618, Z => net11944);
   U1015 : EXOR2DL port map( A1 => n618, A2 => n481, Z => net11941);
   U1016 : OAI22D1 port map( A1 => n28, A2 => n722, B1 => n723, B2 => n30, Z =>
                           n591);
   U1017 : OAI22DL port map( A1 => n768, A2 => n12, B1 => n1017, B2 => n9, Z =>
                           n633);
   U1018 : EXNOR2DL port map( A1 => b(9), A2 => a(3), Z => n1017);
   U1019 : OAI22DL port map( A1 => n738, A2 => n24, B1 => n737, B2 => n22, Z =>
                           n605);
   U1020 : NAN2DL port map( A1 => net11982, A2 => n576, Z => net9975);
   U1021 : NAN2DL port map( A1 => n576, A2 => n632, Z => net9974);
   U1022 : NAN2DL port map( A1 => net11982, A2 => n632, Z => net9976);
   U1023 : NAN2D1 port map( A1 => n647, A2 => n562, Z => net12114);
   U1024 : AOI21DL port map( A1 => net12275, A2 => n956, B => n926, Z => n195);
   U1025 : OAI21M20D2 port map( A1 => net12274, A2 => net12275, B => n183, Z =>
                           net12273);
   U1026 : BUFDL port map( A => net12275, Z => net11686);
   U1027 : OAI21D1 port map( A1 => n243, A2 => n231, B => n1028, Z => n230);
   U1028 : AO21D1 port map( A1 => n230, A2 => n211, B => n212, Z => net12315);
   U1029 : NAN2DL port map( A1 => n474, A2 => n483, Z => n1027);
   U1030 : NAN2D1 port map( A1 => n484, A2 => n491, Z => n1025);
   U1031 : NAN2D1 port map( A1 => n233, A2 => n1023, Z => n231);
   U1032 : OR2D1 port map( A1 => n1026, A2 => n491, Z => n1023);
   U1033 : EXOR3DL port map( A1 => n493, A2 => n488, A3 => n486, Z => n1026);
   U1034 : INVDL port map( A => n235, Z => n233);
   U1035 : AND2D1 port map( A1 => n492, A2 => n499, Z => n1020);
   U1036 : OR2D1 port map( A1 => n492, A2 => n499, Z => n1021);
   U1037 : OAI21D1 port map( A1 => net11339, A2 => n261, B => n250, Z => n248);
   U1038 : AND2DL port map( A1 => n500, A2 => n505, Z => n1022);
   U1039 : AND2DL port map( A1 => n506, A2 => n511, Z => n1024);
   U1040 : AND2DL port map( A1 => n512, A2 => n515, Z => n1019);
   U1041 : NAN2DL port map( A1 => n516, A2 => n519, Z => n268);
   U1042 : AND2D1 port map( A1 => n520, A2 => n521, Z => n1018);
   U1043 : OAI22D1 port map( A1 => n707, A2 => n36, B1 => n1029, B2 => n34, Z 
                           => n576);
   U1044 : EXNOR2DL port map( A1 => a(11), A2 => b(2), Z => n1029);
   U1045 : NAN2D1 port map( A1 => n1031, A2 => n1032, Z => n767);
   U1046 : NAN2D1 port map( A1 => net11996, A2 => net12160, Z => n1032);
   U1047 : NAN2DL port map( A1 => b(9), A2 => a(3), Z => n1031);
   U1048 : EXOR2D2 port map( A1 => n176, A2 => n63, Z => product(20));
   U1049 : INVDL port map( A => n174, Z => n294);
   U1050 : AOI21D1 port map( A1 => net12273, A2 => n295, B => n178, Z => n176);
   U1051 : INVDL port map( A => n180, Z => n178);
   U1052 : INVDL port map( A => n179, Z => n295);
   U1053 : NAN2DL port map( A1 => n295, A2 => n180, Z => n64);
   U1054 : NAN2D1 port map( A1 => n364, A2 => n373, Z => n175);
   U1055 : NOR2D2 port map( A1 => n364, A2 => n373, Z => n174);
   U1056 : NOR2D1 port map( A1 => n179, A2 => n174, Z => n168);
   U1057 : OAI21DL port map( A1 => n194, A2 => n186, B => n187, Z => n185);
   U1058 : NOR2DL port map( A1 => n191, A2 => n186, Z => n1033);
   U1059 : AND2D1 port map( A1 => n184, A2 => n196, Z => net12274);
   U1060 : NOR2D1 port map( A1 => n191, A2 => n186, Z => n184);
   U1061 : NOR2D1 port map( A1 => n374, A2 => n385, Z => n179);
   U1062 : OAI21DL port map( A1 => n199, A2 => net12005, B => n1010, Z => n190)
                           ;
   U1063 : AND2DL port map( A1 => n296, A2 => n187, Z => net11247);
   U1064 : NOR2M1DL port map( A1 => n955, A2 => net12005, Z => n189);
   U1065 : EXOR2D1 port map( A1 => net11941, A2 => net12148, Z => n468);
   U1066 : BUFDL port map( A => n479, Z => net12148);
   U1067 : NAN3D2 port map( A1 => n1034, A2 => n1035, A3 => n1036, Z => n475);
   U1068 : NAN2D1 port map( A1 => n489, A2 => n480, Z => n1036);
   U1069 : NAN2D1 port map( A1 => n487, A2 => n480, Z => n1035);
   U1070 : NAN2D1 port map( A1 => n487, A2 => n489, Z => n1034);
   U1071 : NAN2D1 port map( A1 => n479, A2 => n618, Z => net11943);
   U1072 : EXOR3D1 port map( A1 => n487, A2 => n489, A3 => n480, Z => n476);
   U1073 : OAI21D1 port map( A1 => n217, A2 => n213, B => n214, Z => n212);
   U1074 : AOI21DL port map( A1 => net12350, A2 => n218, B => n219, Z => 
                           net12187);
   U1075 : NAN2D1 port map( A1 => n452, A2 => n1037, Z => n221);
   U1076 : NAN3M1DL port map( A1 => net11961, A2 => net9971, A3 => net9972, Z 
                           => n1037);
   U1077 : ADFULDL port map( A => n465, B => n456, CI => n454, CO => n451, S =>
                           n452);
   U1078 : NAN2D1 port map( A1 => n440, A2 => n451, Z => n214);
   U1079 : NAN3M1D1 port map( A1 => net11961, A2 => net9971, A3 => net9972, Z 
                           => n463);
   U1080 : NAN3D2 port map( A1 => net9968, A2 => net9967, A3 => net9969, Z => 
                           n465);
   U1081 : EXOR3D1 port map( A1 => n446, A2 => n448, A3 => n455, Z => n442);
   U1082 : NAN2DL port map( A1 => n448, A2 => n455, Z => net11524);
   U1083 : NAN2DL port map( A1 => n446, A2 => n455, Z => net11523);
   U1084 : NAN3D1 port map( A1 => net9976, A2 => net9974, A3 => net9975, Z => 
                           n469);
   U1085 : INVDL port map( A => net11981, Z => net11982);
   U1086 : NOR2D1 port map( A1 => n213, A2 => n216, Z => n211);
   U1087 : INVDL port map( A => n213, Z => n300);
   U1088 : NAN2D1 port map( A1 => n300, A2 => n214, Z => n69);
   U1089 : EXOR3D1 port map( A1 => n413, A2 => n402, A3 => n1040, Z => n1038);
   U1090 : INVD1 port map( A => n1039, Z => n1040);
   U1091 : INVDL port map( A => n400, Z => n1039);
   U1092 : NAN2DL port map( A1 => n386, A2 => n397, Z => n187);
   U1093 : AND2D1 port map( A1 => n299, A2 => n954, Z => net9959);
   U1094 : INVDL port map( A => n954, Z => n206);
   U1095 : INVDL port map( A => n202, Z => n298);
   U1096 : INVDL port map( A => a(7), Z => net11920);
   U1097 : NAN2D1 port map( A1 => b(5), A2 => a(7), Z => n1043);
   U1098 : NAN2D2 port map( A1 => n1041, A2 => n22, Z => n24);
   U1099 : EXOR2DL port map( A1 => a(7), A2 => a(6), Z => n1041);
   U1100 : EXNOR2D4 port map( A1 => a(5), A2 => a(6), Z => n22);
   U1101 : NAN2D1 port map( A1 => b(8), A2 => a(5), Z => n1073);
   U1102 : EXNOR2D1 port map( A1 => net12273, A2 => n64, Z => product(19));
   U1103 : EXNOR2DL port map( A1 => b(2), A2 => a(13), Z => n1045);
   U1104 : OAI22D1 port map( A1 => n34, A2 => n701, B1 => n702, B2 => n36, Z =>
                           n571);
   U1105 : EXNOR2D4 port map( A1 => a(9), A2 => a(10), Z => n34);
   U1106 : NAN2D1 port map( A1 => b(0), A2 => a(15), Z => n1046);
   U1107 : NAN2D2 port map( A1 => net12321, A2 => n835, Z => n1047);
   U1108 : NAN2D1 port map( A1 => n1046, A2 => n1047, Z => n674);
   U1109 : INVD16 port map( A => b(0), Z => net12321);
   U1110 : NAN2DL port map( A1 => n424, A2 => n437, Z => n1049);
   U1111 : NAN2D1 port map( A1 => n435, A2 => n437, Z => n1050);
   U1112 : INVDL port map( A => n406, Z => n1051);
   U1113 : INVD1 port map( A => n1051, Z => n1052);
   U1114 : INVDL port map( A => n207, Z => n299);
   U1115 : EXNOR2DL port map( A1 => b(10), A2 => a(11), Z => n698);
   U1116 : AOI21D1 port map( A1 => net12184, A2 => n95, B => n96, Z => n94);
   U1117 : NAN2D1 port map( A1 => b(14), A2 => a(3), Z => n1054);
   U1118 : NAN2D2 port map( A1 => n1053, A2 => net12160, Z => n1055);
   U1119 : NAN2D2 port map( A1 => n1054, A2 => n1055, Z => n762);
   U1120 : INVD4 port map( A => b(14), Z => n1053);
   U1121 : NOR2DL port map( A1 => n398, A2 => n411, Z => net12262);
   U1122 : EXOR2D1 port map( A1 => b(8), A2 => n1056, Z => n717);
   U1123 : NAN3D1 port map( A1 => n1133, A2 => net11523, A3 => net11524, Z => 
                           n441);
   U1124 : EXOR2D1 port map( A1 => n158, A2 => n61, Z => product(22));
   U1125 : NAN2D1 port map( A1 => b(1), A2 => n1058, Z => n1059);
   U1126 : NAN2D1 port map( A1 => n957, A2 => n835, Z => n1060);
   U1127 : NAN2D1 port map( A1 => n1059, A2 => n1060, Z => n673);
   U1128 : INVD1 port map( A => n835, Z => n1058);
   U1129 : NAN2DL port map( A1 => b(0), A2 => a(13), Z => n1062);
   U1130 : NAN2D1 port map( A1 => net12321, A2 => n1061, Z => n1063);
   U1131 : NAN2D1 port map( A1 => n1062, A2 => n1063, Z => n691);
   U1132 : INVDL port map( A => a(13), Z => n1061);
   U1133 : AOI21DL port map( A1 => n169, A2 => n139, B => n140, Z => n52);
   U1134 : NAN2D1 port map( A1 => n590, A2 => n647, Z => n1070);
   U1135 : ADFULD2 port map( A => n593, B => n621, CI => n635, CO => n495, S =>
                           n496);
   U1136 : OAI22D1 port map( A1 => n740, A2 => n24, B1 => n1069, B2 => n22, Z 
                           => n607);
   U1137 : BUFDL port map( A => net12273, Z => net12184);
   U1138 : OAI22D2 port map( A1 => n674, A2 => n48, B1 => n1089, B2 => n46, Z 
                           => n545);
   U1139 : OAI22DL port map( A1 => n916, A2 => n24, B1 => n735, B2 => n22, Z =>
                           n1065);
   U1140 : EXNOR2DL port map( A1 => b(10), A2 => a(3), Z => n1066);
   U1141 : EXNOR2D1 port map( A1 => b(2), A2 => a(5), Z => n757);
   U1142 : NAN2M1D1 port map( A1 => b(0), A2 => a(13), Z => n692);
   U1143 : INVD20 port map( A => b(3), Z => n1084);
   U1144 : OAI22DL port map( A1 => n758, A2 => n18, B1 => n757, B2 => n16, Z =>
                           n624);
   U1145 : OAI22D1 port map( A1 => n781, A2 => n6, B1 => n780, B2 => n834, Z =>
                           n646);
   U1146 : EXNOR2D2 port map( A1 => b(4), A2 => a(5), Z => n755);
   U1147 : EXNOR2DL port map( A1 => b(3), A2 => a(7), Z => n1069);
   U1148 : EXNOR2D2 port map( A1 => b(1), A2 => a(11), Z => n707);
   U1149 : EXNOR2D1 port map( A1 => b(10), A2 => a(3), Z => n766);
   U1150 : EXNOR2D1 port map( A1 => b(5), A2 => a(13), Z => n686);
   U1151 : NAN2DL port map( A1 => n590, A2 => n562, Z => n1071);
   U1152 : NAN3D2 port map( A1 => n1070, A2 => net12114, A3 => n1071, Z => n471
                           );
   U1153 : EXNOR2D1 port map( A1 => b(4), A2 => a(9), Z => n721);
   U1154 : NAN2D1 port map( A1 => net11021, A2 => n1149, Z => net11339);
   U1155 : INVD2 port map( A => b(8), Z => n1072);
   U1156 : NAN2D1 port map( A1 => n1077, A2 => n441, Z => n1078);
   U1157 : NAN2D1 port map( A1 => n1076, A2 => n430, Z => n1079);
   U1158 : INVDL port map( A => n441, Z => n1076);
   U1159 : NAN2D1 port map( A1 => n1085, A2 => n1086, Z => n1080);
   U1160 : NAN2D2 port map( A1 => n1084, A2 => net11946, Z => n1086);
   U1161 : AOI21D1 port map( A1 => net11686, A2 => n189, B => n190, Z => n188);
   U1162 : BUFDL port map( A => net12262, Z => net12005);
   U1163 : EXNOR2D1 port map( A1 => b(7), A2 => a(7), Z => n735);
   U1164 : ADFULDL port map( A => n383, B => n540, CI => n611, CO => n371, S =>
                           n372);
   U1165 : EXNOR2DL port map( A1 => b(9), A2 => a(15), Z => n665);
   U1166 : EXNOR2D2 port map( A1 => b(9), A2 => a(7), Z => n733);
   U1167 : EXNOR2D1 port map( A1 => b(9), A2 => a(1), Z => n784);
   U1168 : EXOR2D1 port map( A1 => b(1), A2 => n1056, Z => n724);
   U1169 : NAN2D1 port map( A1 => b(3), A2 => a(11), Z => n1085);
   U1170 : EXNOR2DL port map( A1 => b(14), A2 => a(1), Z => n1082);
   U1171 : EXNOR2DL port map( A1 => b(14), A2 => a(1), Z => n779);
   U1172 : EXNOR2D1 port map( A1 => b(9), A2 => a(5), Z => n750);
   U1173 : OAI22DL port map( A1 => n1066, A2 => n12, B1 => n765, B2 => n9, Z =>
                           n1083);
   U1174 : NAN2D2 port map( A1 => n1110, A2 => n1056, Z => n1112);
   U1175 : ADFULD2 port map( A => n592, B => n634, CI => n620, CO => n487, S =>
                           n488);
   U1176 : OAI22D2 port map( A1 => n724, A2 => n30, B1 => n917, B2 => n28, Z =>
                           n592);
   U1177 : OAI22D2 port map( A1 => n690, A2 => n42, B1 => n1045, B2 => n40, Z 
                           => n560);
   U1178 : NAN3D2 port map( A1 => net11942, A2 => net11943, A3 => net11944, Z 
                           => n467);
   U1179 : NAN2D1 port map( A1 => n1085, A2 => n1086, Z => n705);
   U1180 : EXOR2D1 port map( A1 => b(2), A2 => net11946, Z => n706);
   U1181 : EXNOR2D1 port map( A1 => b(6), A2 => a(7), Z => n736);
   U1182 : NAN2D1 port map( A1 => b(7), A2 => a(5), Z => n1087);
   U1183 : NAN2D2 port map( A1 => n1126, A2 => net12088, Z => n1088);
   U1184 : EXOR2D1 port map( A1 => b(1), A2 => n835, Z => n1089);
   U1185 : OAI22DL port map( A1 => n720, A2 => n30, B1 => n719, B2 => n28, Z =>
                           n588);
   U1186 : EXOR3D2 port map( A1 => n434, A2 => n447, A3 => n445, Z => n430);
   U1187 : EXNOR2DL port map( A1 => b(11), A2 => a(5), Z => n1090);
   U1188 : EXOR3D1 port map( A1 => n419, A2 => n1052, A3 => n408, Z => n402);
   U1189 : NAN2DL port map( A1 => n408, A2 => n419, Z => n1095);
   U1190 : EXNOR2DL port map( A1 => b(5), A2 => a(15), Z => n669);
   U1191 : EXNOR2DL port map( A1 => b(5), A2 => a(5), Z => n754);
   U1192 : EXNOR2DL port map( A1 => b(5), A2 => a(9), Z => n720);
   U1193 : NAN2D2 port map( A1 => n1126, A2 => n1056, Z => n1128);
   U1194 : INVD16 port map( A => b(7), Z => n1126);
   U1195 : EXNOR2DL port map( A1 => b(13), A2 => a(3), Z => n1091);
   U1196 : NAN2DL port map( A1 => n406, A2 => n408, Z => n1093);
   U1197 : NAN2DL port map( A1 => n406, A2 => n419, Z => n1094);
   U1198 : NAN3D1 port map( A1 => n1094, A2 => n1095, A3 => n1093, Z => n401);
   U1199 : NAN2DL port map( A1 => n599, A2 => n557, Z => n1096);
   U1200 : NAN2DL port map( A1 => n599, A2 => n585, Z => n1097);
   U1201 : NAN2DL port map( A1 => n557, A2 => n585, Z => n1098);
   U1202 : OAI22DL port map( A1 => n687, A2 => n42, B1 => n686, B2 => n40, Z =>
                           n557);
   U1203 : EXOR2DL port map( A1 => n570, A2 => n584, Z => n1129);
   U1204 : NAN2DL port map( A1 => n584, A2 => n570, Z => n1132);
   U1205 : NAN2DL port map( A1 => n407, A2 => n570, Z => n1131);
   U1206 : NAN2D2 port map( A1 => n1127, A2 => n1128, Z => n718);
   U1207 : EXOR3D2 port map( A1 => n603, A2 => n631, A3 => n646, Z => n460);
   U1208 : NAN2DL port map( A1 => n1065, A2 => n646, Z => n1099);
   U1209 : NAN2DL port map( A1 => n1065, A2 => n1083, Z => n1100);
   U1210 : NAN2DL port map( A1 => n646, A2 => n1083, Z => n1101);
   U1211 : NAN3D1 port map( A1 => n1099, A2 => n1101, A3 => n1100, Z => n459);
   U1212 : OAI22D2 port map( A1 => n764, A2 => n12, B1 => n1091, B2 => n9, Z =>
                           n629);
   U1213 : INVDL port map( A => n427, Z => n1102);
   U1214 : INVDL port map( A => n1102, Z => n1103);
   U1215 : EXNOR2DL port map( A1 => b(6), A2 => a(5), Z => n1104);
   U1216 : EXOR2D1 port map( A1 => n147, A2 => n60, Z => product(23));
   U1217 : OAI22D1 port map( A1 => n784, A2 => n6, B1 => n1109, B2 => n834, Z 
                           => n649);
   U1218 : OAI22DL port map( A1 => n785, A2 => n6, B1 => n784, B2 => n834, Z =>
                           n650);
   U1219 : EXNOR2DL port map( A1 => b(8), A2 => a(5), Z => n1105);
   U1220 : EXNOR2DL port map( A1 => b(4), A2 => a(9), Z => n1106);
   U1221 : EXNOR2DL port map( A1 => b(11), A2 => a(1), Z => n1107);
   U1222 : EXNOR2DL port map( A1 => b(11), A2 => a(1), Z => n782);
   U1223 : EXNOR2DL port map( A1 => b(7), A2 => a(5), Z => n1108);
   U1224 : NAN2D1 port map( A1 => b(3), A2 => a(9), Z => n1111);
   U1225 : EXNOR2DL port map( A1 => b(10), A2 => a(1), Z => n1109);
   U1226 : OAI22D1 port map( A1 => n671, A2 => n48, B1 => n670, B2 => n46, Z =>
                           n542);
   U1227 : NAN2D1 port map( A1 => b(7), A2 => a(9), Z => n1127);
   U1228 : NAN2DL port map( A1 => n428, A2 => n430, Z => n1114);
   U1229 : NAN2DL port map( A1 => n430, A2 => n441, Z => n1116);
   U1230 : NAN3D1 port map( A1 => n1114, A2 => n1116, A3 => n1115, Z => n425);
   U1231 : AOI21DL port map( A1 => n115, A2 => net12273, B => n116, Z => n114);
   U1232 : NAN2D1 port map( A1 => n434, A2 => n445, Z => n1117);
   U1233 : NAN2D1 port map( A1 => n434, A2 => n447, Z => n1118);
   U1234 : NAN2D1 port map( A1 => n445, A2 => n447, Z => n1119);
   U1235 : NAN3D2 port map( A1 => n1117, A2 => n1119, A3 => n1118, Z => n429);
   U1236 : NAN2D1 port map( A1 => n429, A2 => n418, Z => n1121);
   U1237 : NAN2D1 port map( A1 => n431, A2 => n418, Z => n1122);
   U1238 : NAN3D2 port map( A1 => n1120, A2 => n1121, A3 => n1122, Z => n413);
   U1239 : NAN2DL port map( A1 => n1103, A2 => n416, Z => n1123);
   U1240 : NAN2DL port map( A1 => n1103, A2 => n414, Z => n1124);
   U1241 : NAN2DL port map( A1 => n416, A2 => n414, Z => n1125);
   U1242 : EXNOR2DL port map( A1 => b(7), A2 => a(13), Z => n684);
   U1243 : EXNOR2DL port map( A1 => b(7), A2 => a(3), Z => n769);
   U1244 : EXNOR2DL port map( A1 => b(7), A2 => a(15), Z => n667);
   U1245 : EXNOR2DL port map( A1 => b(7), A2 => a(1), Z => n786);
   U1246 : EXOR2D1 port map( A1 => n1129, A2 => n407, Z => n392);
   U1247 : NAN2D1 port map( A1 => n407, A2 => n584, Z => n1130);
   U1248 : NAN3D1 port map( A1 => n1130, A2 => n1132, A3 => n1131, Z => n391);
   U1249 : INVDL port map( A => n1006, Z => n296);
   U1250 : EXOR3D2 port map( A1 => n619, A2 => n648, A3 => n577, Z => n480);
   U1251 : NAN2DL port map( A1 => n446, A2 => n448, Z => n1133);
   U1252 : NAN2DL port map( A1 => n453, A2 => n444, Z => n1134);
   U1253 : NAN2DL port map( A1 => n453, A2 => n442, Z => n1135);
   U1254 : NAN2DL port map( A1 => n444, A2 => n442, Z => n1136);
   U1255 : NAN3D1 port map( A1 => n1134, A2 => n1135, A3 => n1136, Z => n439);
   U1256 : EXOR2D4 port map( A1 => n943, A2 => n524, Z => n462);
   U1257 : EXOR2D2 port map( A1 => n167, A2 => n62, Z => product(21));
   U1258 : AOI21D1 port map( A1 => net12273, A2 => n168, B => n169, Z => n167);
   U1259 : NOR2DL port map( A1 => n112, A2 => n103, Z => n101);
   U1260 : NAN2D1 port map( A1 => n619, A2 => n577, Z => n1137);
   U1261 : NAN2D1 port map( A1 => n619, A2 => n648, Z => n1138);
   U1262 : NAN2D1 port map( A1 => n577, A2 => n648, Z => n1139);
   U1263 : NAN3D2 port map( A1 => n1137, A2 => n1139, A3 => n1138, Z => n479);
   U1264 : NAN2D2 port map( A1 => n1140, A2 => n1141, Z => n619);
   U1265 : EXNOR2D4 port map( A1 => a(3), A2 => a(4), Z => n16);
   U1266 : INVDL port map( A => n162, Z => n164);
   U1267 : EXNOR2DL port map( A1 => n215, A2 => n69, Z => product(14));
   U1268 : INVDL port map( A => n53, Z => n135);
   U1269 : EXNOR2D2 port map( A1 => n188, A2 => net11247, Z => product(18));
   U1270 : INVDL port map( A => n120, Z => n118);
   U1271 : INVDL port map( A => n119, Z => n117);
   U1272 : NAN2DL port map( A1 => n1146, A2 => n146, Z => n60);
   U1273 : NAN2DL port map( A1 => n293, A2 => n162, Z => n62);
   U1274 : NAN2DL port map( A1 => n1145, A2 => n157, Z => n61);
   U1275 : EXNOR2D2 port map( A1 => n134, A2 => n941, Z => product(24));
   U1276 : AND2DL port map( A1 => n289, A2 => n126, Z => n1144);
   U1277 : EXNOR2D2 port map( A1 => n127, A2 => n1144, Z => product(25));
   U1278 : AOI21DL port map( A1 => n164, A2 => n1145, B => n155, Z => n151);
   U1279 : OA21M20DL port map( A1 => n155, A2 => n1146, B => n146, Z => n142);
   U1280 : NAN2DL port map( A1 => n293, A2 => n1145, Z => n150);
   U1281 : NOR2DL port map( A1 => n53, A2 => n130, Z => n128);
   U1282 : EXNOR2D2 port map( A1 => n105, A2 => n1142, Z => product(27));
   U1283 : AND2DL port map( A1 => n287, A2 => n104, Z => n1142);
   U1284 : NAN2DL port map( A1 => n288, A2 => n113, Z => n57);
   U1285 : OA21M20DL port map( A1 => n120, A2 => n288, B => n113, Z => n109);
   U1286 : NAN2DL port map( A1 => n346, A2 => n353, Z => n157);
   U1287 : NAN2M1DL port map( A1 => n92, A2 => n93, Z => n55);
   U1288 : OR2DL port map( A1 => n97, A2 => n92, Z => n1148);
   U1289 : NOR2D1 port map( A1 => n516, A2 => n519, Z => n267);
   U1290 : NOR2D1 port map( A1 => n522, A2 => n641, Z => n275);
   U1291 : AND2DL port map( A1 => n657, A2 => n642, Z => n1151);
   U1292 : OAI22DL port map( A1 => n793, A2 => n6, B1 => n792, B2 => n834, Z =>
                           n658);
   U1293 : OAI22DL port map( A1 => n698, A2 => n36, B1 => n697, B2 => n34, Z =>
                           n567);
   U1294 : NAN2DL port map( A1 => n315, A2 => n942, Z => n84);
   U1295 : OAI22DL port map( A1 => n665, A2 => n48, B1 => n664, B2 => n46, Z =>
                           n536);
   U1296 : OAI22DL port map( A1 => n661, A2 => n48, B1 => n660, B2 => n46, Z =>
                           n532);
   U1297 : OAI22DL port map( A1 => n789, A2 => n6, B1 => n788, B2 => n834, Z =>
                           n654);
   U1298 : OAI22DL port map( A1 => n791, A2 => n6, B1 => n790, B2 => n834, Z =>
                           n656);
   U1299 : NAN2D2 port map( A1 => n1143, A2 => n16, Z => n18);
   U1300 : EXOR2DL port map( A1 => a(5), A2 => a(4), Z => n1143);
   U1301 : EXNOR2DL port map( A1 => b(15), A2 => a(15), Z => n659);
   U1302 : EXNOR2DL port map( A1 => a(3), A2 => a(2), Z => n1155);
   U1303 : EXNOR2DL port map( A1 => a(1), A2 => a(0), Z => n1156);
   U1304 : INVDL port map( A => net12262, Z => n297);
   U1305 : INVDL port map( A => n1064, Z => n136);
   U1306 : NAN2D1 port map( A1 => n168, A2 => n139, Z => n53);
   U1307 : NOR2DL port map( A1 => n53, A2 => n108, Z => n106);
   U1308 : INVD1 port map( A => n168, Z => n170);
   U1309 : NOR2DL port map( A1 => n53, A2 => n97, Z => n95);
   U1310 : NOR2D1 port map( A1 => n170, A2 => n150, Z => n148);
   U1311 : INVDL port map( A => n130, Z => n290);
   U1312 : NOR2D1 port map( A1 => n141, A2 => n161, Z => n139);
   U1313 : NAN2D1 port map( A1 => n1145, A2 => n1146, Z => n141);
   U1314 : INVD1 port map( A => n157, Z => n155);
   U1315 : INVDL port map( A => n161, Z => n293);
   U1316 : NOR2D1 port map( A1 => n130, A2 => n125, Z => n119);
   U1317 : NAN2D1 port map( A1 => n119, A2 => n288, Z => n108);
   U1318 : NOR2DL port map( A1 => n53, A2 => n1148, Z => n86);
   U1319 : NAN2DL port map( A1 => n119, A2 => n101, Z => n97);
   U1320 : NOR2DL port map( A1 => n53, A2 => n117, Z => n115);
   U1321 : INVD1 port map( A => n103, Z => n287);
   U1322 : OR2D1 port map( A1 => n346, A2 => n353, Z => n1145);
   U1323 : NAN2D1 port map( A1 => n354, A2 => n363, Z => n162);
   U1324 : OR2D1 port map( A1 => n338, A2 => n345, Z => n1146);
   U1325 : NAN2D1 port map( A1 => n338, A2 => n345, Z => n146);
   U1326 : OA21DL port map( A1 => n100, A2 => n92, B => n93, Z => n1147);
   U1327 : NAN2D1 port map( A1 => n332, A2 => n337, Z => n133);
   U1328 : NAN2DL port map( A1 => n326, A2 => n331, Z => n126);
   U1329 : INVD1 port map( A => n112, Z => n288);
   U1330 : INVDL port map( A => n409, Z => n410);
   U1331 : OR2D1 port map( A1 => n500, A2 => n505, Z => net11021);
   U1332 : OR2D1 port map( A1 => n506, A2 => n511, Z => n1149);
   U1333 : INVD2 port map( A => n343, Z => n344);
   U1334 : NOR2D1 port map( A1 => n325, A2 => n322, Z => n112);
   U1335 : NAN2D1 port map( A1 => n325, A2 => n322, Z => n113);
   U1336 : NOR2D1 port map( A1 => n318, A2 => n321, Z => n103);
   U1337 : NAN2DL port map( A1 => n318, A2 => n321, Z => n104);
   U1338 : NOR2D1 port map( A1 => n317, A2 => n316, Z => n92);
   U1339 : NAN2DL port map( A1 => n317, A2 => n316, Z => n93);
   U1340 : INVDL port map( A => n383, Z => n384);
   U1341 : AO21D1 port map( A1 => n12, A2 => n9, B => n761, Z => n627);
   U1342 : EXNOR2D1 port map( A1 => n600, A2 => n558, Z => n424);
   U1343 : OR2D1 port map( A1 => n512, A2 => n515, Z => net10923);
   U1344 : AO21D1 port map( A1 => n18, A2 => n16, B => n744, Z => n611);
   U1345 : AO21D1 port map( A1 => n24, A2 => n22, B => n727, Z => n595);
   U1346 : OR2D1 port map( A1 => n520, A2 => n521, Z => net10919);
   U1347 : INVDL port map( A => n361, Z => n362);
   U1348 : NAN2DL port map( A1 => n522, A2 => n641, Z => n276);
   U1349 : NAN2D1 port map( A1 => n1153, A2 => n84, Z => n54);
   U1350 : OR2D1 port map( A1 => n657, A2 => n642, Z => n1150);
   U1351 : AND2D1 port map( A1 => n658, A2 => n530, Z => n1152);
   U1352 : INVD1 port map( A => n329, Z => n330);
   U1353 : AO21D1 port map( A1 => n30, A2 => n28, B => n710, Z => n579);
   U1354 : AO21D1 port map( A1 => n36, A2 => n34, B => n693, Z => n563);
   U1355 : INVDL port map( A => n319, Z => n320);
   U1356 : AO21D1 port map( A1 => n42, A2 => n40, B => n676, Z => n547);
   U1357 : OR2D1 port map( A1 => n315, A2 => n942, Z => n1153);
   U1358 : INVDL port map( A => a(15), Z => n835);
   U1359 : NAN2D2 port map( A1 => n812, A2 => n40, Z => n42);
   U1360 : NAN2D2 port map( A1 => n814, A2 => n28, Z => n30);
   U1361 : NAN2M1D2 port map( A1 => n1154, A2 => n34, Z => n36);
   U1362 : EXNOR2DL port map( A1 => a(11), A2 => a(10), Z => n1154);
   U1363 : NAN2M1D2 port map( A1 => n1155, A2 => n9, Z => n12);
   U1364 : EXNOR2D2 port map( A1 => a(13), A2 => a(14), Z => n46);
   U1365 : NAN2D2 port map( A1 => n811, A2 => n46, Z => n48);
   U1366 : NAN2M1D2 port map( A1 => n1156, A2 => n834, Z => n6);
   U1367 : INVDL port map( A => a(1), Z => n842);
   U1368 : INVDL port map( A => n169, Z => n171);
   U1369 : EXNOR2DL port map( A1 => b(1), A2 => a(5), Z => n758);
   U1370 : NAN2DL port map( A1 => n412, A2 => n425, Z => n203);
   U1371 : EXOR2D1 port map( A1 => net12315, A2 => net9959, Z => product(15));
   U1372 : EXNOR2D2 port map( A1 => n195, A2 => net9957, Z => product(17));
   U1373 : EXNOR2D2 port map( A1 => n204, A2 => n1157, Z => product(16));
   U1374 : AND2DL port map( A1 => n203, A2 => n298, Z => n1157);
   U1375 : OAI21DL port map( A1 => n1064, A2 => n1148, B => n1147, Z => n87);
   U1376 : OAI21DL port map( A1 => n1064, A2 => n97, B => n100, Z => n96);
   U1377 : OAI21DL port map( A1 => n1064, A2 => n108, B => n109, Z => n107);
   U1378 : AOI21DL port map( A1 => net12184, A2 => n86, B => n87, Z => n85);
   U1379 : AOI21DL port map( A1 => n106, A2 => net12273, B => n107, Z => n105);
   U1380 : AOI21DL port map( A1 => n135, A2 => net12273, B => n136, Z => n134);
   U1381 : AOI21DL port map( A1 => n128, A2 => net12273, B => n129, Z => n127);
   U1382 : EXNOR2D4 port map( A1 => a(1), A2 => a(2), Z => n9);
   U1383 : EXNOR2D4 port map( A1 => a(7), A2 => a(8), Z => n28);
   U1384 : EXNOR2D4 port map( A1 => a(11), A2 => a(12), Z => n40);

end hier_sec_par_16_5;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_siso_gen.all;

architecture hier_sec_par_16_5 of siso_gen_DW_mult_tc_9 is

   component BUFD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22M10D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OA22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AO21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INVDL
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFD4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AO21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22DL
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFD20
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component ADHALFD1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component NOR2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n15, n16, n17, n18, 
      n19, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33, n34, n35, n36
      , n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n51, n54, n55, n56, 
      n57, n58, n59, n60, n61, n62, n64, n65, n66, n67, n68, n69, n84, n85, n86
      , n87, n92, n93, n94, n95, n96, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n112, n113, n114, n115, n116, n121, n123, 
      n124, n125, n126, n127, n128, n129, n132, n133, n134, n135, n136, n139, 
      n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n170, n171, n172, n173, n174, n175, n176, n177, n178, 
      n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, 
      n191, n192, n193, n194, n195, n197, n198, n199, n200, n201, n202, n203, 
      n204, n205, n206, n207, n208, n209, n210, n213, n214, n215, n216, n217, 
      n229, n230, n231, n232, n243, n248, n249, n250, n261, n266, n267, n268, 
      n269, n274, n275, n276, n277, n294, n315, n316, n317, n318, n319, n320, 
      n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, 
      n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, 
      n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, 
      n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, 
      n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, 
      n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, 
      n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, 
      n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, 
      n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, 
      n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, 
      n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, 
      n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, 
      n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, 
      n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, 
      n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, 
      n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, 
      n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, 
      n525, n526, n527, n528, n529, n530, n532, n533, n534, n535, n536, n537, 
      n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, 
      n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, 
      n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, 
      n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, 
      n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, 
      n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, 
      n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, 
      n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, 
      n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, 
      n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, 
      n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, 
      n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, 
      n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, 
      n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, 
      n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, 
      n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, 
      n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, 
      n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, 
      n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, 
      n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, 
      n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, 
      n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, 
      n802, n803, n805, n806, n807, n808, n809, n811, n812, n813, n814, n815, 
      n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, 
      n828, n829, n830, n831, n832, n833, n834, n837, n838, n839, n840, n842, 
      n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, 
      n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, 
      n934, n935, n936, n937, n938, n939, n940 : std_logic;

begin
   
   U54 : EXOR2D1 port map( A1 => n85, A2 => n54, Z => product(29));
   U59 : EXOR2D1 port map( A1 => n94, A2 => n55, Z => product(28));
   U60 : AOI21D1 port map( A1 => n51, A2 => n86, B => n87, Z => n85);
   U62 : OAI21D1 port map( A1 => n913, A2 => n920, B => n919, Z => n87);
   U71 : EXOR2D1 port map( A1 => n105, A2 => n56, Z => product(27));
   U74 : OAI21D1 port map( A1 => n913, A2 => n99, B => n100, Z => n96);
   U78 : AOI21D1 port map( A1 => n124, A2 => n101, B => n102, Z => n100);
   U80 : OAI21D1 port map( A1 => n113, A2 => n103, B => n104, Z => n102);
   U85 : EXOR2D1 port map( A1 => n114, A2 => n57, Z => product(26));
   U88 : OAI21D1 port map( A1 => n913, A2 => n108, B => n109, Z => n107);
   U97 : EXOR2D1 port map( A1 => n127, A2 => n58, Z => product(25));
   U108 : OAI21D1 port map( A1 => n133, A2 => n125, B => n126, Z => n124);
   U113 : EXOR2D1 port map( A1 => n134, A2 => n59, Z => product(24));
   U116 : OAI21D1 port map( A1 => n913, A2 => n132, B => n133, Z => n129);
   U123 : EXOR2D1 port map( A1 => n147, A2 => n60, Z => product(23));
   U132 : AOI21D1 port map( A1 => n155, A2 => n143, B => n144, Z => n142);
   U137 : NOR2D2 port map( A1 => n338, A2 => n345, Z => n145);
   U139 : EXOR2D1 port map( A1 => n158, A2 => n61, Z => product(22));
   U142 : OAI21D1 port map( A1 => n171, A2 => n150, B => n151, Z => n149);
   U144 : AOI21D1 port map( A1 => n164, A2 => n152, B => n155, Z => n151);
   U153 : EXOR2D1 port map( A1 => n167, A2 => n62, Z => product(21));
   U156 : OAI21D1 port map( A1 => n171, A2 => n161, B => n162, Z => n160);
   U163 : NOR2D2 port map( A1 => n354, A2 => n363, Z => n165);
   U166 : AOI21D1 port map( A1 => n51, A2 => n168, B => n173, Z => n167);
   U172 : OAI21D1 port map( A1 => n174, A2 => n180, B => n175, Z => n173);
   U175 : NOR2D2 port map( A1 => n364, A2 => n373, Z => n174);
   U177 : EXNOR2D1 port map( A1 => n51, A2 => n64, Z => product(19));
   U178 : AOI21D1 port map( A1 => n51, A2 => n177, B => n178, Z => n176);
   U184 : NAN2D2 port map( A1 => n374, A2 => n385, Z => n180);
   U185 : EXOR2D1 port map( A1 => n188, A2 => n65, Z => product(18));
   U186 : OAI21D1 port map( A1 => n182, A2 => n210, B => n183, Z => n181);
   U188 : AOI21D1 port map( A1 => n201, A2 => n184, B => n185, Z => n183);
   U190 : OAI21D1 port map( A1 => n186, A2 => n194, B => n187, Z => n185);
   U193 : NOR2D2 port map( A1 => n386, A2 => n397, Z => n186);
   U195 : EXOR2D1 port map( A1 => n195, A2 => n66, Z => product(17));
   U198 : OAI21D1 port map( A1 => n199, A2 => n191, B => n194, Z => n190);
   U203 : NOR2D2 port map( A1 => n398, A2 => n411, Z => n193);
   U205 : EXOR2D1 port map( A1 => n204, A2 => n67, Z => product(16));
   U212 : OAI21D1 port map( A1 => n202, A2 => n208, B => n203, Z => n201);
   U215 : NOR2D2 port map( A1 => n412, A2 => n425, Z => n202);
   U217 : EXNOR2D1 port map( A1 => n209, A2 => n68, Z => product(15));
   U218 : AOI21D1 port map( A1 => n209, A2 => n205, B => n206, Z => n204);
   U223 : NOR2D2 port map( A1 => n426, A2 => n439, Z => n207);
   U224 : NAN2D2 port map( A1 => n426, A2 => n439, Z => n208);
   U225 : EXNOR2D1 port map( A1 => n215, A2 => n69, Z => product(14));
   U232 : NOR2D2 port map( A1 => n440, A2 => n451, Z => n213);
   U237 : AOI21D1 port map( A1 => n925, A2 => n910, B => n917, Z => n217);
   U256 : OAI21D1 port map( A1 => n243, A2 => n231, B => n232, Z => n230);
   U258 : AOI21D1 port map( A1 => n921, A2 => n923, B => n924, Z => n232);
   U275 : AOI21D1 port map( A1 => n248, A2 => n928, B => n931, Z => n243);
   U283 : OAI21D1 port map( A1 => n249, A2 => n261, B => n250, Z => n248);
   U285 : AOI21D1 port map( A1 => n926, A2 => n929, B => n927, Z => n250);
   U302 : AOI21D1 port map( A1 => n266, A2 => n933, B => n934, Z => n261);
   U310 : OAI21D1 port map( A1 => n267, A2 => n269, B => n268, Z => n266);
   U316 : AOI21D1 port map( A1 => n274, A2 => n935, B => n936, Z => n269);
   U324 : OAI21D1 port map( A1 => n275, A2 => n277, B => n276, Z => n274);
   U330 : AOI21D1 port map( A1 => n937, A2 => n939, B => n938, Z => n277);
   U344 : ADFULD1 port map( A => n532, B => n319, CI => n547, CO => n315, S => 
                           n316);
   U345 : ADFULD1 port map( A => n320, B => n533, CI => n323, CO => n317, S => 
                           n318);
   U347 : ADFULD1 port map( A => n327, B => n563, CI => n324, CO => n321, S => 
                           n322);
   U348 : ADFULD1 port map( A => n548, B => n329, CI => n534, CO => n323, S => 
                           n324);
   U349 : ADFULD1 port map( A => n328, B => n335, CI => n333, CO => n325, S => 
                           n326);
   U350 : ADFULD1 port map( A => n535, B => n549, CI => n330, CO => n327, S => 
                           n328);
   U352 : ADFULD1 port map( A => n339, B => n336, CI => n334, CO => n331, S => 
                           n332);
   U353 : ADFULD1 port map( A => n579, B => n564, CI => n341, CO => n333, S => 
                           n334);
   U354 : ADFULD1 port map( A => n550, B => n536, CI => n343, CO => n335, S => 
                           n336);
   U355 : ADFULD1 port map( A => n347, B => n342, CI => n340, CO => n337, S => 
                           n338);
   U356 : ADFULD1 port map( A => n351, B => n344, CI => n349, CO => n339, S => 
                           n340);
   U357 : ADFULD1 port map( A => n551, B => n537, CI => n565, CO => n341, S => 
                           n342);
   U359 : ADFULD1 port map( A => n348, B => n357, CI => n355, CO => n345, S => 
                           n346);
   U360 : ADFULD1 port map( A => n352, B => n359, CI => n350, CO => n347, S => 
                           n348);
   U361 : ADFULD1 port map( A => n566, B => n552, CI => n595, CO => n349, S => 
                           n350);
   U362 : ADFULD1 port map( A => n580, B => n538, CI => n361, CO => n351, S => 
                           n352);
   U363 : ADFULD1 port map( A => n365, B => n358, CI => n356, CO => n353, S => 
                           n354);
   U364 : ADFULD1 port map( A => n360, B => n369, CI => n367, CO => n355, S => 
                           n356);
   U365 : ADFULD1 port map( A => n362, B => n567, CI => n371, CO => n357, S => 
                           n358);
   U366 : ADFULD1 port map( A => n581, B => n553, CI => n539, CO => n359, S => 
                           n360);
   U368 : ADFULD1 port map( A => n375, B => n368, CI => n366, CO => n363, S => 
                           n364);
   U369 : ADFULD1 port map( A => n372, B => n370, CI => n377, CO => n365, S => 
                           n366);
   U370 : ADFULD1 port map( A => n381, B => n611, CI => n379, CO => n367, S => 
                           n368);
   U371 : ADFULD1 port map( A => n554, B => n582, CI => n596, CO => n369, S => 
                           n370);
   U372 : ADFULD1 port map( A => n383, B => n540, CI => n568, CO => n371, S => 
                           n372);
   U373 : ADFULD1 port map( A => n387, B => n378, CI => n376, CO => n373, S => 
                           n374);
   U374 : ADFULD1 port map( A => n391, B => n380, CI => n389, CO => n375, S => 
                           n376);
   U375 : ADFULD1 port map( A => n393, B => n395, CI => n382, CO => n377, S => 
                           n378);
   U376 : ADFULD1 port map( A => n541, B => n555, CI => n384, CO => n379, S => 
                           n380);
   U377 : ADFULD1 port map( A => n597, B => n569, CI => n583, CO => n381, S => 
                           n382);
   U379 : ADFULD1 port map( A => n399, B => n390, CI => n388, CO => n385, S => 
                           n386);
   U380 : ADFULD1 port map( A => n392, B => n403, CI => n401, CO => n387, S => 
                           n388);
   U381 : ADFULD1 port map( A => n394, B => n405, CI => n396, CO => n389, S => 
                           n390);
   U382 : ADFULD1 port map( A => n627, B => n584, CI => n407, CO => n391, S => 
                           n392);
   U383 : ADFULD1 port map( A => n570, B => n598, CI => n612, CO => n393, S => 
                           n394);
   U384 : ADFULD1 port map( A => n409, B => n542, CI => n556, CO => n395, S => 
                           n396);
   U385 : ADFULD1 port map( A => n413, B => n402, CI => n400, CO => n397, S => 
                           n398);
   U386 : ADFULD1 port map( A => n404, B => n417, CI => n415, CO => n399, S => 
                           n400);
   U387 : ADFULD1 port map( A => n406, B => n419, CI => n408, CO => n401, S => 
                           n402);
   U388 : ADFULD1 port map( A => n423, B => n410, CI => n421, CO => n403, S => 
                           n404);
   U389 : ADFULD1 port map( A => n557, B => n599, CI => n585, CO => n405, S => 
                           n406);
   U390 : ADFULD1 port map( A => n543, B => n571, CI => n613, CO => n407, S => 
                           n408);
   U392 : ADFULD1 port map( A => n427, B => n416, CI => n414, CO => n411, S => 
                           n412);
   U393 : ADFULD1 port map( A => n429, B => n431, CI => n418, CO => n413, S => 
                           n414);
   U394 : ADFULD1 port map( A => n422, B => n433, CI => n420, CO => n415, S => 
                           n416);
   U395 : ADFULD1 port map( A => n424, B => n437, CI => n435, CO => n417, S => 
                           n418);
   U396 : ADFULD1 port map( A => n614, B => n628, CI => n643, CO => n419, S => 
                           n420);
   U397 : ADFULD1 port map( A => n544, B => n586, CI => n572, CO => n421, S => 
                           n422);
   U400 : ADFULD1 port map( A => n441, B => n430, CI => n428, CO => n425, S => 
                           n426);
   U401 : ADFULD1 port map( A => n443, B => n436, CI => n432, CO => n427, S => 
                           n428);
   U402 : ADFULD1 port map( A => n445, B => n447, CI => n434, CO => n429, S => 
                           n430);
   U403 : ADFULD1 port map( A => n438, B => n615, CI => n449, CO => n431, S => 
                           n432);
   U404 : ADFULD1 port map( A => n629, B => n573, CI => n601, CO => n433, S => 
                           n434);
   U405 : ADFULD1 port map( A => n545, B => n587, CI => n559, CO => n435, S => 
                           n436);
   U406 : ADHALFD1 port map( A => n523, B => n644, CO => n437, S => n438);
   U407 : ADFULD1 port map( A => n453, B => n444, CI => n442, CO => n439, S => 
                           n440);
   U408 : ADFULD1 port map( A => n446, B => n448, CI => n455, CO => n441, S => 
                           n442);
   U409 : ADFULD1 port map( A => n457, B => n459, CI => n450, CO => n443, S => 
                           n444);
   U410 : ADFULD1 port map( A => n588, B => n602, CI => n461, CO => n445, S => 
                           n446);
   U411 : ADFULD1 port map( A => n560, B => n616, CI => n574, CO => n447, S => 
                           n448);
   U412 : ADFULD1 port map( A => n645, B => n546, CI => n630, CO => n449, S => 
                           n450);
   U413 : ADFULD1 port map( A => n465, B => n456, CI => n454, CO => n451, S => 
                           n452);
   U414 : ADFULD1 port map( A => n460, B => n458, CI => n467, CO => n453, S => 
                           n454);
   U415 : ADFULD1 port map( A => n471, B => n462, CI => n469, CO => n455, S => 
                           n456);
   U416 : ADFULD1 port map( A => n561, B => n603, CI => n575, CO => n457, S => 
                           n458);
   U417 : ADFULD1 port map( A => n631, B => n589, CI => n617, CO => n459, S => 
                           n460);
   U418 : ADHALFD1 port map( A => n524, B => n646, CO => n461, S => n462);
   U419 : ADFULD1 port map( A => n468, B => n475, CI => n466, CO => n463, S => 
                           n464);
   U420 : ADFULD1 port map( A => n470, B => n472, CI => n477, CO => n465, S => 
                           n466);
   U421 : ADFULD1 port map( A => n481, B => n604, CI => n479, CO => n467, S => 
                           n468);
   U422 : ADFULD1 port map( A => n576, B => n618, CI => n590, CO => n469, S => 
                           n470);
   U423 : ADFULD1 port map( A => n647, B => n562, CI => n632, CO => n471, S => 
                           n472);
   U424 : ADFULD1 port map( A => n485, B => n478, CI => n476, CO => n473, S => 
                           n474);
   U425 : ADFULD1 port map( A => n487, B => n489, CI => n480, CO => n475, S => 
                           n476);
   U426 : ADFULD1 port map( A => n591, B => n619, CI => n482, CO => n477, S => 
                           n478);
   U427 : ADFULD1 port map( A => n577, B => n605, CI => n633, CO => n479, S => 
                           n480);
   U429 : ADFULD1 port map( A => n493, B => n488, CI => n486, CO => n483, S => 
                           n484);
   U430 : ADFULD1 port map( A => n495, B => n497, CI => n490, CO => n485, S => 
                           n486);
   U431 : ADFULD1 port map( A => n592, B => n620, CI => n606, CO => n487, S => 
                           n488);
   U432 : ADFULD1 port map( A => n649, B => n578, CI => n634, CO => n489, S => 
                           n490);
   U433 : ADFULD1 port map( A => n496, B => n501, CI => n494, CO => n491, S => 
                           n492);
   U434 : ADFULD1 port map( A => n498, B => n635, CI => n503, CO => n493, S => 
                           n494);
   U435 : ADFULD1 port map( A => n593, B => n607, CI => n621, CO => n495, S => 
                           n496);
   U437 : ADFULD1 port map( A => n504, B => n507, CI => n502, CO => n499, S => 
                           n500);
   U438 : ADFULD1 port map( A => n608, B => n622, CI => n509, CO => n501, S => 
                           n502);
   U439 : ADFULD1 port map( A => n651, B => n594, CI => n636, CO => n503, S => 
                           n504);
   U440 : ADFULD1 port map( A => n513, B => n510, CI => n508, CO => n505, S => 
                           n506);
   U441 : ADFULD1 port map( A => n609, B => n637, CI => n623, CO => n507, S => 
                           n508);
   U443 : ADFULD1 port map( A => n517, B => n624, CI => n514, CO => n511, S => 
                           n512);
   U444 : ADFULD1 port map( A => n653, B => n610, CI => n638, CO => n513, S => 
                           n514);
   U445 : ADFULD1 port map( A => n625, B => n639, CI => n518, CO => n515, S => 
                           n516);
   U447 : ADFULD1 port map( A => n655, B => n626, CI => n640, CO => n519, S => 
                           n520);
   U451 : OAI22D1 port map( A1 => n46, A2 => n660, B1 => n48, B2 => n661, Z => 
                           n532);
   U452 : OAI22D1 port map( A1 => n46, A2 => n661, B1 => n48, B2 => n662, Z => 
                           n533);
   U453 : OAI22D1 port map( A1 => n46, A2 => n662, B1 => n48, B2 => n663, Z => 
                           n534);
   U454 : OAI22D1 port map( A1 => n46, A2 => n663, B1 => n48, B2 => n664, Z => 
                           n535);
   U455 : OAI22D1 port map( A1 => n46, A2 => n664, B1 => n48, B2 => n665, Z => 
                           n536);
   U456 : OAI22D1 port map( A1 => n46, A2 => n665, B1 => n48, B2 => n666, Z => 
                           n537);
   U457 : OAI22D1 port map( A1 => n45, A2 => n666, B1 => n47, B2 => n667, Z => 
                           n538);
   U458 : OAI22D1 port map( A1 => n45, A2 => n667, B1 => n47, B2 => n668, Z => 
                           n539);
   U459 : OAI22D1 port map( A1 => n45, A2 => n668, B1 => n47, B2 => n669, Z => 
                           n540);
   U460 : OAI22D1 port map( A1 => n45, A2 => n669, B1 => n47, B2 => n670, Z => 
                           n541);
   U461 : OAI22D1 port map( A1 => n45, A2 => n670, B1 => n47, B2 => n671, Z => 
                           n542);
   U462 : OAI22D1 port map( A1 => n45, A2 => n671, B1 => n47, B2 => n672, Z => 
                           n543);
   U463 : OAI22D1 port map( A1 => n45, A2 => n672, B1 => n47, B2 => n673, Z => 
                           n544);
   U464 : OAI22D1 port map( A1 => n45, A2 => n673, B1 => n47, B2 => n674, Z => 
                           n545);
   U465 : NOR2M1D1 port map( A1 => b(0), A2 => n45, Z => n546);
   U466 : EXNOR2D1 port map( A1 => n43, A2 => n795, Z => n659);
   U467 : EXNOR2D1 port map( A1 => n43, A2 => n796, Z => n660);
   U468 : EXNOR2D1 port map( A1 => n43, A2 => n797, Z => n661);
   U469 : EXNOR2D1 port map( A1 => n43, A2 => n798, Z => n662);
   U470 : EXNOR2D1 port map( A1 => n43, A2 => n799, Z => n663);
   U471 : EXNOR2D1 port map( A1 => n43, A2 => n800, Z => n664);
   U472 : EXNOR2D1 port map( A1 => n43, A2 => n801, Z => n665);
   U473 : EXNOR2D1 port map( A1 => n43, A2 => n802, Z => n666);
   U474 : EXNOR2D1 port map( A1 => n43, A2 => n803, Z => n667);
   U475 : EXNOR2D1 port map( A1 => n43, A2 => b(6), Z => n668);
   U476 : EXNOR2D1 port map( A1 => n43, A2 => n805, Z => n669);
   U477 : EXNOR2D1 port map( A1 => n43, A2 => n806, Z => n670);
   U478 : EXNOR2D1 port map( A1 => n43, A2 => n807, Z => n671);
   U479 : EXNOR2D1 port map( A1 => n43, A2 => n808, Z => n672);
   U480 : EXNOR2D1 port map( A1 => n43, A2 => n809, Z => n673);
   U481 : EXNOR2D1 port map( A1 => n43, A2 => b(0), Z => n674);
   U482 : NAN2M1D1 port map( A1 => b(0), A2 => n43, Z => n675);
   U485 : OAI22D1 port map( A1 => n40, A2 => n676, B1 => n42, B2 => n677, Z => 
                           n319);
   U486 : OAI22D1 port map( A1 => n40, A2 => n677, B1 => n42, B2 => n678, Z => 
                           n548);
   U487 : OAI22D1 port map( A1 => n40, A2 => n678, B1 => n42, B2 => n679, Z => 
                           n549);
   U488 : OAI22D1 port map( A1 => n40, A2 => n679, B1 => n42, B2 => n680, Z => 
                           n550);
   U489 : OAI22D1 port map( A1 => n40, A2 => n680, B1 => n42, B2 => n681, Z => 
                           n551);
   U490 : OAI22D1 port map( A1 => n40, A2 => n681, B1 => n42, B2 => n682, Z => 
                           n552);
   U491 : OAI22D1 port map( A1 => n40, A2 => n682, B1 => n42, B2 => n683, Z => 
                           n553);
   U492 : OAI22D1 port map( A1 => n39, A2 => n683, B1 => n41, B2 => n684, Z => 
                           n554);
   U493 : OAI22D1 port map( A1 => n39, A2 => n684, B1 => n41, B2 => n685, Z => 
                           n555);
   U494 : OAI22D1 port map( A1 => n39, A2 => n685, B1 => n41, B2 => n686, Z => 
                           n556);
   U495 : OAI22D1 port map( A1 => n39, A2 => n686, B1 => n41, B2 => n687, Z => 
                           n557);
   U496 : OAI22D1 port map( A1 => n39, A2 => n687, B1 => n41, B2 => n688, Z => 
                           n558);
   U497 : OAI22D1 port map( A1 => n39, A2 => n688, B1 => n41, B2 => n689, Z => 
                           n559);
   U498 : OAI22D1 port map( A1 => n39, A2 => n689, B1 => n41, B2 => n690, Z => 
                           n560);
   U499 : OAI22D1 port map( A1 => n39, A2 => n690, B1 => n41, B2 => n691, Z => 
                           n561);
   U500 : NOR2M1D1 port map( A1 => b(0), A2 => n39, Z => n562);
   U501 : EXNOR2D1 port map( A1 => n37, A2 => n795, Z => n676);
   U502 : EXNOR2D1 port map( A1 => n37, A2 => n796, Z => n677);
   U503 : EXNOR2D1 port map( A1 => n37, A2 => n797, Z => n678);
   U504 : EXNOR2D1 port map( A1 => n37, A2 => n798, Z => n679);
   U505 : EXNOR2D1 port map( A1 => n37, A2 => n799, Z => n680);
   U506 : EXNOR2D1 port map( A1 => n37, A2 => n800, Z => n681);
   U507 : EXNOR2D1 port map( A1 => n37, A2 => n801, Z => n682);
   U508 : EXNOR2D1 port map( A1 => n37, A2 => n802, Z => n683);
   U509 : EXNOR2D1 port map( A1 => n37, A2 => n803, Z => n684);
   U510 : EXNOR2D1 port map( A1 => n37, A2 => b(6), Z => n685);
   U511 : EXNOR2D1 port map( A1 => n37, A2 => n805, Z => n686);
   U512 : EXNOR2D1 port map( A1 => n37, A2 => n806, Z => n687);
   U513 : EXNOR2D1 port map( A1 => n37, A2 => n807, Z => n688);
   U514 : EXNOR2D1 port map( A1 => n37, A2 => n808, Z => n689);
   U515 : EXNOR2D1 port map( A1 => n37, A2 => n809, Z => n690);
   U516 : EXNOR2D1 port map( A1 => n37, A2 => b(0), Z => n691);
   U517 : NAN2M1D1 port map( A1 => b(0), A2 => n37, Z => n692);
   U518 : OAI22D1 port map( A1 => n34, A2 => n709, B1 => n36, B2 => n837, Z => 
                           n525);
   U520 : OAI22D1 port map( A1 => n34, A2 => n693, B1 => n36, B2 => n694, Z => 
                           n329);
   U521 : OAI22D1 port map( A1 => n34, A2 => n694, B1 => n36, B2 => n695, Z => 
                           n564);
   U522 : OAI22D1 port map( A1 => n34, A2 => n695, B1 => n36, B2 => n696, Z => 
                           n565);
   U523 : OAI22D1 port map( A1 => n34, A2 => n696, B1 => n36, B2 => n697, Z => 
                           n566);
   U524 : OAI22D1 port map( A1 => n34, A2 => n697, B1 => n36, B2 => n698, Z => 
                           n567);
   U525 : OAI22D1 port map( A1 => n34, A2 => n698, B1 => n36, B2 => n699, Z => 
                           n568);
   U526 : OAI22D1 port map( A1 => n34, A2 => n699, B1 => n36, B2 => n700, Z => 
                           n569);
   U527 : OAI22D1 port map( A1 => n33, A2 => n700, B1 => n35, B2 => n701, Z => 
                           n570);
   U528 : OAI22D1 port map( A1 => n33, A2 => n701, B1 => n35, B2 => n702, Z => 
                           n571);
   U529 : OAI22D1 port map( A1 => n33, A2 => n702, B1 => n35, B2 => n703, Z => 
                           n572);
   U530 : OAI22D1 port map( A1 => n33, A2 => n703, B1 => n35, B2 => n704, Z => 
                           n573);
   U531 : OAI22D1 port map( A1 => n33, A2 => n704, B1 => n35, B2 => n705, Z => 
                           n574);
   U532 : OAI22D1 port map( A1 => n33, A2 => n705, B1 => n35, B2 => n706, Z => 
                           n575);
   U533 : OAI22D1 port map( A1 => n33, A2 => n706, B1 => n35, B2 => n707, Z => 
                           n576);
   U534 : OAI22D1 port map( A1 => n33, A2 => n707, B1 => n35, B2 => n708, Z => 
                           n577);
   U535 : NOR2M1D1 port map( A1 => b(0), A2 => n33, Z => n578);
   U536 : EXNOR2D1 port map( A1 => n31, A2 => n795, Z => n693);
   U537 : EXNOR2D1 port map( A1 => n31, A2 => n796, Z => n694);
   U538 : EXNOR2D1 port map( A1 => n31, A2 => n797, Z => n695);
   U539 : EXNOR2D1 port map( A1 => n31, A2 => n798, Z => n696);
   U540 : EXNOR2D1 port map( A1 => n31, A2 => n799, Z => n697);
   U541 : EXNOR2D1 port map( A1 => n31, A2 => n800, Z => n698);
   U542 : EXNOR2D1 port map( A1 => n31, A2 => n801, Z => n699);
   U543 : EXNOR2D1 port map( A1 => n31, A2 => n802, Z => n700);
   U544 : EXNOR2D1 port map( A1 => n31, A2 => n803, Z => n701);
   U545 : EXNOR2D1 port map( A1 => n31, A2 => b(6), Z => n702);
   U546 : EXNOR2D1 port map( A1 => n31, A2 => n805, Z => n703);
   U547 : EXNOR2D1 port map( A1 => n31, A2 => n806, Z => n704);
   U548 : EXNOR2D1 port map( A1 => n31, A2 => n807, Z => n705);
   U549 : EXNOR2D1 port map( A1 => n31, A2 => n808, Z => n706);
   U550 : EXNOR2D1 port map( A1 => n31, A2 => n809, Z => n707);
   U551 : EXNOR2D1 port map( A1 => n31, A2 => b(0), Z => n708);
   U552 : NAN2M1D1 port map( A1 => b(0), A2 => n31, Z => n709);
   U553 : OAI22D1 port map( A1 => n28, A2 => n726, B1 => n30, B2 => n838, Z => 
                           n526);
   U555 : OAI22D1 port map( A1 => n28, A2 => n710, B1 => n30, B2 => n711, Z => 
                           n343);
   U556 : OAI22D1 port map( A1 => n28, A2 => n711, B1 => n30, B2 => n712, Z => 
                           n580);
   U557 : OAI22D1 port map( A1 => n28, A2 => n712, B1 => n30, B2 => n713, Z => 
                           n581);
   U558 : OAI22D1 port map( A1 => n28, A2 => n713, B1 => n30, B2 => n714, Z => 
                           n582);
   U559 : OAI22D1 port map( A1 => n28, A2 => n714, B1 => n30, B2 => n715, Z => 
                           n583);
   U560 : OAI22D1 port map( A1 => n28, A2 => n715, B1 => n30, B2 => n716, Z => 
                           n584);
   U561 : OAI22D1 port map( A1 => n28, A2 => n716, B1 => n30, B2 => n717, Z => 
                           n585);
   U562 : OAI22D1 port map( A1 => n27, A2 => n717, B1 => n29, B2 => n718, Z => 
                           n586);
   U563 : OAI22D1 port map( A1 => n27, A2 => n718, B1 => n29, B2 => n719, Z => 
                           n587);
   U564 : OAI22D1 port map( A1 => n27, A2 => n719, B1 => n29, B2 => n720, Z => 
                           n588);
   U565 : OAI22D1 port map( A1 => n27, A2 => n720, B1 => n29, B2 => n721, Z => 
                           n589);
   U566 : OAI22D1 port map( A1 => n27, A2 => n721, B1 => n29, B2 => n722, Z => 
                           n590);
   U567 : OAI22D1 port map( A1 => n27, A2 => n722, B1 => n29, B2 => n723, Z => 
                           n591);
   U568 : OAI22D1 port map( A1 => n27, A2 => n723, B1 => n29, B2 => n724, Z => 
                           n592);
   U569 : OAI22D1 port map( A1 => n27, A2 => n724, B1 => n29, B2 => n725, Z => 
                           n593);
   U570 : NOR2M1D1 port map( A1 => b(0), A2 => n27, Z => n594);
   U571 : EXNOR2D1 port map( A1 => n25, A2 => n795, Z => n710);
   U572 : EXNOR2D1 port map( A1 => n25, A2 => n796, Z => n711);
   U573 : EXNOR2D1 port map( A1 => n25, A2 => n797, Z => n712);
   U574 : EXNOR2D1 port map( A1 => n25, A2 => n798, Z => n713);
   U575 : EXNOR2D1 port map( A1 => n25, A2 => n799, Z => n714);
   U576 : EXNOR2D1 port map( A1 => n25, A2 => n800, Z => n715);
   U577 : EXNOR2D1 port map( A1 => n25, A2 => n801, Z => n716);
   U578 : EXNOR2D1 port map( A1 => n25, A2 => n802, Z => n717);
   U579 : EXNOR2D1 port map( A1 => n25, A2 => n803, Z => n718);
   U580 : EXNOR2D1 port map( A1 => n25, A2 => b(6), Z => n719);
   U581 : EXNOR2D1 port map( A1 => n25, A2 => n805, Z => n720);
   U582 : EXNOR2D1 port map( A1 => n25, A2 => n806, Z => n721);
   U583 : EXNOR2D1 port map( A1 => n25, A2 => n807, Z => n722);
   U584 : EXNOR2D1 port map( A1 => n25, A2 => n808, Z => n723);
   U585 : EXNOR2D1 port map( A1 => n25, A2 => n809, Z => n724);
   U586 : EXNOR2D1 port map( A1 => n25, A2 => b(0), Z => n725);
   U587 : NAN2M1D1 port map( A1 => b(0), A2 => n25, Z => n726);
   U588 : OAI22D1 port map( A1 => n22, A2 => n743, B1 => n24, B2 => n839, Z => 
                           n527);
   U590 : OAI22D1 port map( A1 => n22, A2 => n727, B1 => n24, B2 => n728, Z => 
                           n361);
   U591 : OAI22D1 port map( A1 => n22, A2 => n728, B1 => n24, B2 => n729, Z => 
                           n596);
   U592 : OAI22D1 port map( A1 => n22, A2 => n729, B1 => n24, B2 => n730, Z => 
                           n597);
   U593 : OAI22D1 port map( A1 => n22, A2 => n730, B1 => n24, B2 => n731, Z => 
                           n598);
   U594 : OAI22D1 port map( A1 => n22, A2 => n731, B1 => n24, B2 => n732, Z => 
                           n599);
   U595 : OAI22D1 port map( A1 => n22, A2 => n732, B1 => n24, B2 => n733, Z => 
                           n600);
   U596 : OAI22D1 port map( A1 => n22, A2 => n733, B1 => n24, B2 => n734, Z => 
                           n601);
   U597 : OAI22D1 port map( A1 => n21, A2 => n734, B1 => n23, B2 => n735, Z => 
                           n602);
   U598 : OAI22D1 port map( A1 => n21, A2 => n735, B1 => n23, B2 => n736, Z => 
                           n603);
   U599 : OAI22D1 port map( A1 => n21, A2 => n736, B1 => n23, B2 => n737, Z => 
                           n604);
   U600 : OAI22D1 port map( A1 => n21, A2 => n737, B1 => n23, B2 => n738, Z => 
                           n605);
   U601 : OAI22D1 port map( A1 => n21, A2 => n738, B1 => n23, B2 => n739, Z => 
                           n606);
   U602 : OAI22D1 port map( A1 => n21, A2 => n739, B1 => n23, B2 => n740, Z => 
                           n607);
   U603 : OAI22D1 port map( A1 => n21, A2 => n740, B1 => n23, B2 => n741, Z => 
                           n608);
   U604 : OAI22D1 port map( A1 => n21, A2 => n741, B1 => n23, B2 => n742, Z => 
                           n609);
   U605 : NOR2M1D1 port map( A1 => b(0), A2 => n21, Z => n610);
   U606 : EXNOR2D1 port map( A1 => n19, A2 => n795, Z => n727);
   U607 : EXNOR2D1 port map( A1 => n19, A2 => n796, Z => n728);
   U608 : EXNOR2D1 port map( A1 => n19, A2 => n797, Z => n729);
   U609 : EXNOR2D1 port map( A1 => n19, A2 => n798, Z => n730);
   U610 : EXNOR2D1 port map( A1 => n19, A2 => n799, Z => n731);
   U611 : EXNOR2D1 port map( A1 => n19, A2 => n800, Z => n732);
   U612 : EXNOR2D1 port map( A1 => n19, A2 => n801, Z => n733);
   U613 : EXNOR2D1 port map( A1 => n19, A2 => n802, Z => n734);
   U614 : EXNOR2D1 port map( A1 => n19, A2 => n803, Z => n735);
   U615 : EXNOR2D1 port map( A1 => n19, A2 => b(6), Z => n736);
   U616 : EXNOR2D1 port map( A1 => n19, A2 => n805, Z => n737);
   U617 : EXNOR2D1 port map( A1 => n19, A2 => n806, Z => n738);
   U618 : EXNOR2D1 port map( A1 => n19, A2 => n807, Z => n739);
   U619 : EXNOR2D1 port map( A1 => n19, A2 => n808, Z => n740);
   U620 : EXNOR2D1 port map( A1 => n19, A2 => n809, Z => n741);
   U621 : EXNOR2D1 port map( A1 => n19, A2 => b(0), Z => n742);
   U622 : NAN2M1D1 port map( A1 => b(0), A2 => n19, Z => n743);
   U623 : OAI22D1 port map( A1 => n16, A2 => n760, B1 => n18, B2 => n840, Z => 
                           n528);
   U625 : OAI22D1 port map( A1 => n16, A2 => n744, B1 => n18, B2 => n745, Z => 
                           n383);
   U626 : OAI22D1 port map( A1 => n16, A2 => n745, B1 => n18, B2 => n746, Z => 
                           n612);
   U627 : OAI22D1 port map( A1 => n16, A2 => n746, B1 => n18, B2 => n747, Z => 
                           n613);
   U628 : OAI22D1 port map( A1 => n16, A2 => n747, B1 => n18, B2 => n748, Z => 
                           n614);
   U629 : OAI22D1 port map( A1 => n16, A2 => n748, B1 => n18, B2 => n749, Z => 
                           n615);
   U630 : OAI22D1 port map( A1 => n16, A2 => n749, B1 => n18, B2 => n750, Z => 
                           n616);
   U631 : OAI22D1 port map( A1 => n16, A2 => n750, B1 => n18, B2 => n751, Z => 
                           n617);
   U632 : OAI22D1 port map( A1 => n15, A2 => n751, B1 => n17, B2 => n752, Z => 
                           n618);
   U633 : OAI22D1 port map( A1 => n15, A2 => n752, B1 => n17, B2 => n753, Z => 
                           n619);
   U634 : OAI22D1 port map( A1 => n15, A2 => n753, B1 => n17, B2 => n754, Z => 
                           n620);
   U635 : OAI22D1 port map( A1 => n15, A2 => n754, B1 => n17, B2 => n755, Z => 
                           n621);
   U636 : OAI22D1 port map( A1 => n15, A2 => n755, B1 => n17, B2 => n756, Z => 
                           n622);
   U637 : OAI22D1 port map( A1 => n15, A2 => n756, B1 => n17, B2 => n757, Z => 
                           n623);
   U638 : OAI22D1 port map( A1 => n15, A2 => n757, B1 => n17, B2 => n758, Z => 
                           n624);
   U639 : OAI22D1 port map( A1 => n15, A2 => n758, B1 => n17, B2 => n759, Z => 
                           n625);
   U640 : NOR2M1D1 port map( A1 => b(0), A2 => n15, Z => n626);
   U641 : EXNOR2D1 port map( A1 => n13, A2 => n795, Z => n744);
   U642 : EXNOR2D1 port map( A1 => n13, A2 => n796, Z => n745);
   U643 : EXNOR2D1 port map( A1 => n13, A2 => n797, Z => n746);
   U644 : EXNOR2D1 port map( A1 => n13, A2 => n798, Z => n747);
   U645 : EXNOR2D1 port map( A1 => n13, A2 => n799, Z => n748);
   U646 : EXNOR2D1 port map( A1 => n13, A2 => n800, Z => n749);
   U647 : EXNOR2D1 port map( A1 => n13, A2 => n801, Z => n750);
   U648 : EXNOR2D1 port map( A1 => n13, A2 => n802, Z => n751);
   U649 : EXNOR2D1 port map( A1 => n13, A2 => n803, Z => n752);
   U650 : EXNOR2D1 port map( A1 => n13, A2 => b(6), Z => n753);
   U651 : EXNOR2D1 port map( A1 => n13, A2 => n805, Z => n754);
   U652 : EXNOR2D1 port map( A1 => n13, A2 => n806, Z => n755);
   U653 : EXNOR2D1 port map( A1 => n13, A2 => n807, Z => n756);
   U654 : EXNOR2D1 port map( A1 => n13, A2 => n808, Z => n757);
   U655 : EXNOR2D1 port map( A1 => n13, A2 => n809, Z => n758);
   U656 : EXNOR2D1 port map( A1 => n13, A2 => b(0), Z => n759);
   U657 : NAN2M1D1 port map( A1 => b(0), A2 => n13, Z => n760);
   U660 : OAI22D1 port map( A1 => n10, A2 => n761, B1 => n12, B2 => n762, Z => 
                           n409);
   U661 : OAI22D1 port map( A1 => n10, A2 => n762, B1 => n12, B2 => n763, Z => 
                           n628);
   U662 : OAI22D1 port map( A1 => n10, A2 => n763, B1 => n12, B2 => n764, Z => 
                           n629);
   U663 : OAI22D1 port map( A1 => n10, A2 => n764, B1 => n12, B2 => n765, Z => 
                           n630);
   U664 : OAI22D1 port map( A1 => n10, A2 => n765, B1 => n12, B2 => n766, Z => 
                           n631);
   U665 : OAI22D1 port map( A1 => n10, A2 => n766, B1 => n12, B2 => n767, Z => 
                           n632);
   U666 : OAI22D1 port map( A1 => n10, A2 => n767, B1 => n12, B2 => n768, Z => 
                           n633);
   U667 : OAI22D1 port map( A1 => n9, A2 => n768, B1 => n11, B2 => n769, Z => 
                           n634);
   U668 : OAI22D1 port map( A1 => n9, A2 => n769, B1 => n11, B2 => n770, Z => 
                           n635);
   U669 : OAI22D1 port map( A1 => n9, A2 => n770, B1 => n11, B2 => n771, Z => 
                           n636);
   U670 : OAI22D1 port map( A1 => n9, A2 => n771, B1 => n11, B2 => n772, Z => 
                           n637);
   U671 : OAI22D1 port map( A1 => n9, A2 => n772, B1 => n11, B2 => n773, Z => 
                           n638);
   U672 : OAI22D1 port map( A1 => n9, A2 => n773, B1 => n11, B2 => n774, Z => 
                           n639);
   U673 : OAI22D1 port map( A1 => n9, A2 => n774, B1 => n11, B2 => n775, Z => 
                           n640);
   U674 : OAI22D1 port map( A1 => n9, A2 => n775, B1 => n11, B2 => n776, Z => 
                           n641);
   U675 : NOR2M1D1 port map( A1 => b(0), A2 => n9, Z => n642);
   U676 : EXNOR2D1 port map( A1 => n7, A2 => n795, Z => n761);
   U677 : EXNOR2D1 port map( A1 => n7, A2 => n796, Z => n762);
   U678 : EXNOR2D1 port map( A1 => n7, A2 => n797, Z => n763);
   U679 : EXNOR2D1 port map( A1 => n7, A2 => n798, Z => n764);
   U680 : EXNOR2D1 port map( A1 => n7, A2 => n799, Z => n765);
   U681 : EXNOR2D1 port map( A1 => n7, A2 => n800, Z => n766);
   U682 : EXNOR2D1 port map( A1 => n7, A2 => n801, Z => n767);
   U683 : EXNOR2D1 port map( A1 => n7, A2 => n802, Z => n768);
   U684 : EXNOR2D1 port map( A1 => n7, A2 => n803, Z => n769);
   U685 : EXNOR2D1 port map( A1 => n7, A2 => b(6), Z => n770);
   U686 : EXNOR2D1 port map( A1 => n7, A2 => n805, Z => n771);
   U687 : EXNOR2D1 port map( A1 => n7, A2 => n806, Z => n772);
   U688 : EXNOR2D1 port map( A1 => n7, A2 => n807, Z => n773);
   U689 : EXNOR2D1 port map( A1 => n7, A2 => n808, Z => n774);
   U690 : EXNOR2D1 port map( A1 => n7, A2 => n809, Z => n775);
   U691 : EXNOR2D1 port map( A1 => n7, A2 => b(0), Z => n776);
   U692 : NAN2M1D1 port map( A1 => b(0), A2 => n7, Z => n777);
   U693 : OAI22D1 port map( A1 => n794, A2 => n4, B1 => n6, B2 => n842, Z => 
                           n530);
   U696 : OAI22D1 port map( A1 => n779, A2 => n4, B1 => n6, B2 => n780, Z => 
                           n645);
   U697 : OAI22D1 port map( A1 => n780, A2 => n4, B1 => n6, B2 => n781, Z => 
                           n646);
   U698 : OAI22D1 port map( A1 => n781, A2 => n4, B1 => n6, B2 => n782, Z => 
                           n647);
   U699 : OAI22D1 port map( A1 => n782, A2 => n4, B1 => n6, B2 => n783, Z => 
                           n648);
   U700 : OAI22D1 port map( A1 => n783, A2 => n4, B1 => n6, B2 => n784, Z => 
                           n649);
   U701 : OAI22D1 port map( A1 => n784, A2 => n4, B1 => n6, B2 => n785, Z => 
                           n650);
   U702 : OAI22D1 port map( A1 => n785, A2 => n3, B1 => n5, B2 => n786, Z => 
                           n651);
   U703 : OAI22D1 port map( A1 => n786, A2 => n3, B1 => n5, B2 => n787, Z => 
                           n652);
   U704 : OAI22D1 port map( A1 => n787, A2 => n3, B1 => n5, B2 => n788, Z => 
                           n653);
   U705 : OAI22D1 port map( A1 => n788, A2 => n3, B1 => n5, B2 => n789, Z => 
                           n654);
   U706 : OAI22D1 port map( A1 => n789, A2 => n3, B1 => n5, B2 => n790, Z => 
                           n655);
   U707 : OAI22D1 port map( A1 => n790, A2 => n3, B1 => n5, B2 => n791, Z => 
                           n656);
   U708 : OAI22D1 port map( A1 => n791, A2 => n3, B1 => n5, B2 => n792, Z => 
                           n657);
   U709 : OAI22D1 port map( A1 => n792, A2 => n3, B1 => n5, B2 => n793, Z => 
                           n658);
   U711 : EXNOR2D1 port map( A1 => n1, A2 => n795, Z => n778);
   U712 : EXNOR2D1 port map( A1 => n1, A2 => n796, Z => n779);
   U713 : EXNOR2D1 port map( A1 => n1, A2 => n797, Z => n780);
   U714 : EXNOR2D1 port map( A1 => n1, A2 => n798, Z => n781);
   U715 : EXNOR2D1 port map( A1 => n1, A2 => n799, Z => n782);
   U716 : EXNOR2D1 port map( A1 => n1, A2 => n800, Z => n783);
   U717 : EXNOR2D1 port map( A1 => n1, A2 => n801, Z => n784);
   U718 : EXNOR2D1 port map( A1 => n1, A2 => n802, Z => n785);
   U719 : EXNOR2D1 port map( A1 => n1, A2 => n803, Z => n786);
   U720 : EXNOR2D1 port map( A1 => n1, A2 => b(6), Z => n787);
   U721 : EXNOR2D1 port map( A1 => n1, A2 => n805, Z => n788);
   U722 : EXNOR2D1 port map( A1 => n1, A2 => n806, Z => n789);
   U723 : EXNOR2D1 port map( A1 => n1, A2 => n807, Z => n790);
   U724 : EXNOR2D1 port map( A1 => n1, A2 => n808, Z => n791);
   U725 : EXNOR2D1 port map( A1 => n1, A2 => n809, Z => n792);
   U726 : EXNOR2D1 port map( A1 => n1, A2 => b(0), Z => n793);
   U727 : NAN2M1D1 port map( A1 => b(0), A2 => n1, Z => n794);
   U752 : EXOR2D1 port map( A1 => a(14), A2 => a(15), Z => n811);
   U753 : EXNOR2D1 port map( A1 => a(14), A2 => a(13), Z => n827);
   U755 : EXOR2D1 port map( A1 => a(12), A2 => a(13), Z => n812);
   U756 : EXNOR2D1 port map( A1 => a(12), A2 => a(11), Z => n828);
   U758 : EXOR2D1 port map( A1 => a(10), A2 => a(11), Z => n813);
   U759 : EXNOR2D1 port map( A1 => a(10), A2 => a(9), Z => n829);
   U761 : EXOR2D1 port map( A1 => a(8), A2 => a(9), Z => n814);
   U762 : EXNOR2D1 port map( A1 => a(8), A2 => a(7), Z => n830);
   U764 : EXOR2D1 port map( A1 => a(6), A2 => a(7), Z => n815);
   U765 : EXNOR2D1 port map( A1 => a(6), A2 => a(5), Z => n831);
   U767 : EXOR2D1 port map( A1 => a(4), A2 => a(5), Z => n816);
   U768 : EXNOR2D1 port map( A1 => a(4), A2 => a(3), Z => n832);
   U770 : EXOR2D1 port map( A1 => a(2), A2 => a(3), Z => n817);
   U771 : EXNOR2D1 port map( A1 => a(2), A2 => a(1), Z => n833);
   U773 : EXOR2D1 port map( A1 => a(0), A2 => a(1), Z => n818);
   U777 : BUFD20 port map( A => b(10), Z => n800);
   U778 : NOR2D1 port map( A1 => n193, A2 => n186, Z => n184);
   U779 : INVDL port map( A => n174, Z => n294);
   U780 : AND2D1 port map( A1 => n464, A2 => n473, Z => n910);
   U781 : INVDL port map( A => n156, Z => n154);
   U782 : NOR2D1 port map( A1 => n346, A2 => n353, Z => n156);
   U783 : NOR2D1 port map( A1 => n202, A2 => n207, Z => n200);
   U784 : INVD1 port map( A => n173, Z => n171);
   U785 : NOR2D1 port map( A1 => n332, A2 => n337, Z => n132);
   U786 : BUFD20 port map( A => b(5), Z => n805);
   U787 : BUFD20 port map( A => b(9), Z => n801);
   U788 : EXOR2D1 port map( A1 => n176, A2 => n912, Z => product(20));
   U789 : INVD1 port map( A => n172, Z => n170);
   U790 : AOI21D1 port map( A1 => n51, A2 => n159, B => n160, Z => n158);
   U791 : NAN2D1 port map( A1 => n172, A2 => n139, Z => n911);
   U792 : NAN2M1DL port map( A1 => n145, A2 => n146, Z => n60);
   U793 : AOI21DL port map( A1 => n51, A2 => n148, B => n149, Z => n147);
   U794 : AOI21DL port map( A1 => n51, A2 => n128, B => n129, Z => n127);
   U795 : AOI21DL port map( A1 => n51, A2 => n135, B => n136, Z => n134);
   U796 : AOI21DL port map( A1 => n209, A2 => n200, B => n197, Z => n195);
   U797 : AOI21DL port map( A1 => n189, A2 => n209, B => n190, Z => n188);
   U798 : INVD2 port map( A => n145, Z => n143);
   U799 : NAN2DL port map( A1 => n412, A2 => n425, Z => n203);
   U800 : AOI21DL port map( A1 => n51, A2 => n115, B => n116, Z => n114);
   U801 : AOI21DL port map( A1 => n51, A2 => n106, B => n107, Z => n105);
   U802 : OAI21DL port map( A1 => n229, A2 => n216, B => n217, Z => n215);
   U803 : AOI21DL port map( A1 => n51, A2 => n95, B => n96, Z => n94);
   U804 : NAN2DL port map( A1 => n440, A2 => n451, Z => n214);
   U805 : INVDL port map( A => n409, Z => n410);
   U806 : AND2DL port map( A1 => n512, A2 => n515, Z => n934);
   U807 : NAN2M1DL port map( A1 => n179, A2 => n180, Z => n64);
   U808 : INVDL port map( A => n199, Z => n197);
   U809 : NOR2DL port map( A1 => n198, A2 => n191, Z => n189);
   U810 : INVDL port map( A => n179, Z => n177);
   U811 : NAN2M1DL port map( A1 => n202, A2 => n203, Z => n67);
   U812 : NAN2DL port map( A1 => n294, A2 => n175, Z => n912);
   U813 : NAN2M1DL port map( A1 => n165, A2 => n166, Z => n62);
   U814 : NAN2M1DL port map( A1 => n156, A2 => n157, Z => n61);
   U815 : NAN2M1D1 port map( A1 => n132, A2 => n133, Z => n59);
   U816 : NAN2M1D1 port map( A1 => n125, A2 => n126, Z => n58);
   U817 : NAN2M1DL port map( A1 => n193, A2 => n194, Z => n66);
   U818 : NAN2M1DL port map( A1 => n186, A2 => n187, Z => n65);
   U819 : AOI21D1 port map( A1 => n173, A2 => n139, B => n914, Z => n913);
   U820 : OAI21DL port map( A1 => n141, A2 => n166, B => n142, Z => n914);
   U821 : INVDL port map( A => n200, Z => n198);
   U822 : INVDL port map( A => n166, Z => n164);
   U823 : AOI21D1 port map( A1 => n915, A2 => n230, B => n916, Z => n210);
   U824 : NOR2DL port map( A1 => n216, A2 => n213, Z => n915);
   U825 : OAI21D1 port map( A1 => n217, A2 => n213, B => n214, Z => n916);
   U826 : NAN2D1 port map( A1 => n398, A2 => n411, Z => n194);
   U827 : NAN2M1DL port map( A1 => n207, A2 => n208, Z => n68);
   U828 : NAN2M1D1 port map( A1 => n112, A2 => n113, Z => n57);
   U829 : NAN2M1D1 port map( A1 => n103, A2 => n104, Z => n56);
   U830 : NAN2M1DL port map( A1 => n213, A2 => n214, Z => n69);
   U831 : NAN2M1D1 port map( A1 => n92, A2 => n93, Z => n55);
   U832 : NAN2DL port map( A1 => n338, A2 => n345, Z => n146);
   U833 : AND2DL port map( A1 => n452, A2 => n463, Z => n917);
   U834 : OR2D1 port map( A1 => n464, A2 => n473, Z => n918);
   U835 : NAN2DL port map( A1 => n921, A2 => n922, Z => n231);
   U836 : AND2D1 port map( A1 => n484, A2 => n491, Z => n923);
   U837 : OR2DL port map( A1 => n600, A2 => n558, Z => n423);
   U838 : OAI22DL port map( A1 => n778, A2 => n4, B1 => n6, B2 => n779, Z => 
                           n644);
   U839 : NOR2D1 port map( A1 => n516, A2 => n519, Z => n267);
   U840 : NAN2DL port map( A1 => n522, A2 => n529, Z => n276);
   U841 : NOR2D1 port map( A1 => n911, A2 => n121, Z => n115);
   U842 : INVD1 port map( A => n911, Z => n135);
   U843 : NOR2D1 port map( A1 => n170, A2 => n150, Z => n148);
   U844 : NOR2D1 port map( A1 => n170, A2 => n161, Z => n159);
   U845 : INVD1 port map( A => n170, Z => n168);
   U846 : NOR2D1 port map( A1 => n911, A2 => n99, Z => n95);
   U847 : AO21M20D1 port map( A1 => n913, A2 => n121, B => n124, Z => n116);
   U848 : INVD1 port map( A => n913, Z => n136);
   U849 : NAN2D1 port map( A1 => n154, A2 => n143, Z => n141);
   U850 : NOR2D1 port map( A1 => n911, A2 => n132, Z => n128);
   U851 : NOR2DL port map( A1 => n911, A2 => n108, Z => n106);
   U852 : INVD1 port map( A => n164, Z => n162);
   U853 : NAN2D1 port map( A1 => n163, A2 => n152, Z => n150);
   U854 : INVD1 port map( A => n156, Z => n152);
   U855 : INVD1 port map( A => n163, Z => n161);
   U856 : INVD1 port map( A => n123, Z => n121);
   U857 : INVDL port map( A => n180, Z => n178);
   U858 : BUFD4 port map( A => n181, Z => n51);
   U859 : NAN2DL port map( A1 => n200, A2 => n184, Z => n182);
   U860 : INVD1 port map( A => n210, Z => n209);
   U861 : NOR2D1 port map( A1 => n141, A2 => n165, Z => n139);
   U862 : NOR2D1 port map( A1 => n374, A2 => n385, Z => n179);
   U863 : NOR2D1 port map( A1 => n179, A2 => n174, Z => n172);
   U864 : INVD1 port map( A => n157, Z => n155);
   U865 : INVDL port map( A => n201, Z => n199);
   U866 : INVD1 port map( A => n146, Z => n144);
   U867 : NOR2DL port map( A1 => n911, A2 => n920, Z => n86);
   U868 : INVD1 port map( A => n192, Z => n191);
   U869 : INVDL port map( A => n193, Z => n192);
   U870 : INVDL port map( A => n165, Z => n163);
   U871 : NOR2D1 port map( A1 => n132, A2 => n125, Z => n123);
   U872 : NAN2D1 port map( A1 => n123, A2 => n110, Z => n108);
   U873 : NAN2D1 port map( A1 => n123, A2 => n101, Z => n99);
   U874 : OA21M20D1 port map( A1 => n124, A2 => n110, B => n113, Z => n109);
   U875 : NAN2DL port map( A1 => n364, A2 => n373, Z => n175);
   U876 : OA21D1 port map( A1 => n100, A2 => n92, B => n93, Z => n919);
   U877 : NAN2D1 port map( A1 => n354, A2 => n363, Z => n166);
   U878 : NAN2D1 port map( A1 => n346, A2 => n353, Z => n157);
   U879 : INVDL port map( A => n230, Z => n229);
   U880 : NAN2DL port map( A1 => n386, A2 => n397, Z => n187);
   U881 : INVDL port map( A => n207, Z => n205);
   U882 : INVDL port map( A => n208, Z => n206);
   U883 : NAN2D1 port map( A1 => n332, A2 => n337, Z => n133);
   U884 : NOR2D1 port map( A1 => n326, A2 => n331, Z => n125);
   U885 : OR2D1 port map( A1 => n99, A2 => n92, Z => n920);
   U886 : NAN2DL port map( A1 => n326, A2 => n331, Z => n126);
   U887 : NOR2D1 port map( A1 => n112, A2 => n103, Z => n101);
   U888 : INVD1 port map( A => n112, Z => n110);
   U889 : OR2D1 port map( A1 => n474, A2 => n483, Z => n921);
   U890 : OR2D1 port map( A1 => n484, A2 => n491, Z => n922);
   U891 : AND2DL port map( A1 => n474, A2 => n483, Z => n924);
   U892 : OR2D1 port map( A1 => n452, A2 => n463, Z => n925);
   U893 : NAN2D1 port map( A1 => n925, A2 => n918, Z => n216);
   U894 : INVDL port map( A => n343, Z => n344);
   U895 : NOR2D1 port map( A1 => n325, A2 => n322, Z => n112);
   U896 : NAN2D1 port map( A1 => n325, A2 => n322, Z => n113);
   U897 : NOR2D1 port map( A1 => n318, A2 => n321, Z => n103);
   U898 : NAN2D1 port map( A1 => n318, A2 => n321, Z => n104);
   U899 : NOR2D1 port map( A1 => n317, A2 => n316, Z => n92);
   U900 : NAN2D1 port map( A1 => n317, A2 => n316, Z => n93);
   U901 : NAN2D1 port map( A1 => n926, A2 => n930, Z => n249);
   U902 : OR2D1 port map( A1 => n500, A2 => n505, Z => n926);
   U903 : AND2DL port map( A1 => n500, A2 => n505, Z => n927);
   U904 : OR2D1 port map( A1 => n492, A2 => n499, Z => n928);
   U905 : AND2D1 port map( A1 => n506, A2 => n511, Z => n929);
   U906 : OR2D1 port map( A1 => n506, A2 => n511, Z => n930);
   U907 : AND2DL port map( A1 => n492, A2 => n499, Z => n931);
   U908 : INVDL port map( A => n383, Z => n384);
   U909 : AO21D1 port map( A1 => n12, A2 => n10, B => n761, Z => n627);
   U910 : EXNOR2D1 port map( A1 => n600, A2 => n558, Z => n424);
   U911 : AO21D1 port map( A1 => n6, A2 => n4, B => n778, Z => n643);
   U912 : AO21D1 port map( A1 => n18, A2 => n16, B => n744, Z => n611);
   U913 : NAN2D1 port map( A1 => n932, A2 => n84, Z => n54);
   U914 : NAN2D1 port map( A1 => n315, A2 => n940, Z => n84);
   U915 : AO21D1 port map( A1 => n24, A2 => n22, B => n727, Z => n595);
   U916 : INVDL port map( A => n361, Z => n362);
   U917 : INVDL port map( A => n329, Z => n330);
   U918 : AO21D1 port map( A1 => n30, A2 => n28, B => n710, Z => n579);
   U919 : AO21D1 port map( A1 => n36, A2 => n34, B => n693, Z => n563);
   U920 : INVD1 port map( A => n319, Z => n320);
   U921 : AO21D1 port map( A1 => n42, A2 => n40, B => n676, Z => n547);
   U922 : OR2D1 port map( A1 => n315, A2 => n940, Z => n932);
   U923 : ADHALFDL port map( A => n527, B => n652, CO => n509, S => n510);
   U924 : INVD1 port map( A => n19, Z => n839);
   U925 : OR2D1 port map( A1 => n512, A2 => n515, Z => n933);
   U926 : ADHALFDL port map( A => n526, B => n650, CO => n497, S => n498);
   U927 : INVD1 port map( A => n25, Z => n838);
   U928 : ADHALFDL port map( A => n525, B => n648, CO => n481, S => n482);
   U929 : INVD1 port map( A => n31, Z => n837);
   U930 : NAN2DL port map( A1 => n516, A2 => n519, Z => n268);
   U931 : OR2D1 port map( A1 => n520, A2 => n521, Z => n935);
   U932 : OAI22M10D1 port map( A1 => n43, A2 => n48, B1 => n46, B2 => n675, Z 
                           => n523);
   U933 : AND2DL port map( A1 => n520, A2 => n521, Z => n936);
   U934 : ADHALFDL port map( A => n528, B => n654, CO => n517, S => n518);
   U935 : INVD1 port map( A => n13, Z => n840);
   U936 : OAI22M10D1 port map( A1 => n37, A2 => n42, B1 => n40, B2 => n692, Z 
                           => n524);
   U937 : NOR2D1 port map( A1 => n522, A2 => n529, Z => n275);
   U938 : OR2D1 port map( A1 => n657, A2 => n642, Z => n937);
   U939 : AND2DL port map( A1 => n657, A2 => n642, Z => n938);
   U940 : AND2D1 port map( A1 => n658, A2 => n530, Z => n939);
   U941 : BUFD1 port map( A => n825, Z => n12);
   U942 : BUFD1 port map( A => n823, Z => n23);
   U943 : BUFD1 port map( A => n825, Z => n11);
   U944 : BUFD1 port map( A => n821, Z => n35);
   U945 : BUFD1 port map( A => n824, Z => n17);
   U946 : BUFD1 port map( A => n823, Z => n24);
   U947 : BUFD1 port map( A => n822, Z => n29);
   U948 : BUFD1 port map( A => n822, Z => n30);
   U949 : BUFD1 port map( A => n821, Z => n36);
   U950 : BUFD1 port map( A => n820, Z => n41);
   U951 : BUFD1 port map( A => n819, Z => n48);
   U952 : BUFD1 port map( A => n819, Z => n47);
   U953 : BUFD1 port map( A => n820, Z => n42);
   U954 : BUFD1 port map( A => n824, Z => n18);
   U955 : BUFD1 port map( A => n833, Z => n10);
   U956 : BUFD1 port map( A => n831, Z => n21);
   U957 : BUFD1 port map( A => n833, Z => n9);
   U958 : BUFD1 port map( A => n829, Z => n33);
   U959 : BUFD1 port map( A => n832, Z => n15);
   U960 : BUFD1 port map( A => n830, Z => n27);
   U961 : BUFD1 port map( A => n831, Z => n22);
   U962 : BUFD1 port map( A => n830, Z => n28);
   U963 : BUFD1 port map( A => n829, Z => n34);
   U964 : BUFD1 port map( A => n826, Z => n6);
   U965 : BUFD1 port map( A => n826, Z => n5);
   U966 : BUFD1 port map( A => n828, Z => n39);
   U967 : BUFD1 port map( A => n827, Z => n45);
   U968 : BUFD1 port map( A => n828, Z => n40);
   U969 : BUFD1 port map( A => n827, Z => n46);
   U970 : OA22D1 port map( A1 => n46, A2 => n659, B1 => n48, B2 => n660, Z => 
                           n940);
   U971 : BUFD1 port map( A => n832, Z => n16);
   U972 : BUFD1 port map( A => n834, Z => n4);
   U973 : BUFD1 port map( A => n834, Z => n3);
   U974 : INVD1 port map( A => n1, Z => n842);
   U975 : BUFD1 port map( A => b(1), Z => n809);
   U976 : BUFD1 port map( A => b(4), Z => n806);
   U977 : BUFD1 port map( A => b(7), Z => n803);
   U978 : BUFD1 port map( A => b(8), Z => n802);
   U979 : BUFD1 port map( A => b(2), Z => n808);
   U980 : BUFD1 port map( A => b(3), Z => n807);
   U981 : BUFD1 port map( A => b(11), Z => n799);
   U982 : BUFD1 port map( A => b(15), Z => n795);
   U983 : BUFD1 port map( A => b(14), Z => n796);
   U984 : BUFD1 port map( A => b(12), Z => n798);
   U985 : BUFD1 port map( A => b(13), Z => n797);
   U986 : ADHALFDL port map( A => n641, B => n656, CO => n521, S => n522);
   U987 : OAI22M10D1 port map( A1 => n7, A2 => n12, B1 => n10, B2 => n777, Z =>
                           n529);
   U988 : NAN2D1 port map( A1 => n817, A2 => n833, Z => n825);
   U989 : NAN2D1 port map( A1 => n815, A2 => n831, Z => n823);
   U990 : NAN2D1 port map( A1 => n813, A2 => n829, Z => n821);
   U991 : NAN2D1 port map( A1 => n816, A2 => n832, Z => n824);
   U992 : NAN2D1 port map( A1 => n814, A2 => n830, Z => n822);
   U993 : NAN2D1 port map( A1 => n812, A2 => n828, Z => n820);
   U994 : NAN2D1 port map( A1 => n811, A2 => n827, Z => n819);
   U995 : NAN2D1 port map( A1 => n818, A2 => n834, Z => n826);
   U996 : INVD1 port map( A => a(0), Z => n834);
   U997 : BUFD1 port map( A => a(1), Z => n1);
   U998 : BUFD1 port map( A => a(7), Z => n19);
   U999 : BUFD1 port map( A => a(11), Z => n31);
   U1000 : BUFD1 port map( A => a(5), Z => n13);
   U1001 : BUFD1 port map( A => a(9), Z => n25);
   U1002 : BUFD1 port map( A => a(3), Z => n7);
   U1003 : BUFD1 port map( A => a(13), Z => n37);
   U1004 : BUFD1 port map( A => a(15), Z => n43);

end hier_sec_par_16_5;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_siso_gen.all;

architecture hier_sec_par_16_5 of siso_gen_DW01_add_7 is

   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVDL
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFD4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21M20DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n21, n22, n23, n24, n25, n26, n27, n29, n30, n31, n32, n33, 
      n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48
      , n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, 
      n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77
      , n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n92, n93, 
      n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n117, n122, n124, n126, n128, 
      n130, n189, n190, n191, n193 : std_logic;

begin
   
   U2 : EXOR2D1 port map( A1 => n22, A2 => n4, Z => SUM(15));
   U7 : EXOR2D1 port map( A1 => n31, A2 => n5, Z => SUM(14));
   U8 : AOI21D1 port map( A1 => n1, A2 => n23, B => n24, Z => n22);
   U10 : OAI21D1 port map( A1 => n2, A2 => n25, B => n26, Z => n24);
   U19 : EXOR2D1 port map( A1 => n40, A2 => n6, Z => SUM(13));
   U22 : OAI21D1 port map( A1 => n2, A2 => n34, B => n35, Z => n33);
   U26 : OAI21D1 port map( A1 => n38, A2 => n46, B => n39, Z => n37);
   U31 : EXOR2D1 port map( A1 => n47, A2 => n7, Z => SUM(12));
   U32 : AOI21D1 port map( A1 => n1, A2 => n41, B => n42, Z => n40);
   U34 : OAI21D1 port map( A1 => n2, A2 => n43, B => n46, Z => n42);
   U39 : NOR2D2 port map( A1 => A(12), A2 => B(12), Z => n45);
   U41 : EXOR2D1 port map( A1 => n54, A2 => n8, Z => SUM(11));
   U46 : AOI21D1 port map( A1 => n50, A2 => n67, B => n51, Z => n2);
   U48 : OAI21D1 port map( A1 => n52, A2 => n60, B => n53, Z => n51);
   U53 : EXOR2D1 port map( A1 => n61, A2 => n9, Z => SUM(10));
   U54 : AOI21D1 port map( A1 => n1, A2 => n55, B => n56, Z => n54);
   U56 : OAI21D1 port map( A1 => n65, A2 => n57, B => n60, Z => n56);
   U61 : NOR2D2 port map( A1 => A(10), A2 => B(10), Z => n59);
   U63 : EXOR2D1 port map( A1 => n70, A2 => n10, Z => SUM(9));
   U64 : AOI21D1 port map( A1 => n1, A2 => n62, B => n63, Z => n61);
   U70 : OAI21D1 port map( A1 => n68, A2 => n74, B => n69, Z => n67);
   U73 : NOR2D2 port map( A1 => A(9), A2 => B(9), Z => n68);
   U75 : EXNOR2D1 port map( A1 => n1, A2 => n11, Z => SUM(8));
   U76 : AOI21D1 port map( A1 => n1, A2 => n71, B => n72, Z => n70);
   U83 : EXOR2D1 port map( A1 => n82, A2 => n12, Z => SUM(7));
   U84 : OAI21D1 port map( A1 => n104, A2 => n76, B => n77, Z => n75);
   U86 : AOI21D1 port map( A1 => n78, A2 => n95, B => n79, Z => n77);
   U88 : OAI21D1 port map( A1 => n80, A2 => n88, B => n81, Z => n79);
   U91 : NOR2D2 port map( A1 => A(7), A2 => B(7), Z => n80);
   U93 : EXOR2D1 port map( A1 => n89, A2 => n13, Z => SUM(6));
   U94 : AOI21D1 port map( A1 => n103, A2 => n83, B => n84, Z => n82);
   U96 : OAI21D1 port map( A1 => n93, A2 => n85, B => n88, Z => n84);
   U101 : NOR2D2 port map( A1 => A(6), A2 => B(6), Z => n87);
   U103 : EXOR2D1 port map( A1 => n98, A2 => n14, Z => SUM(5));
   U104 : AOI21D1 port map( A1 => n103, A2 => n94, B => n95, Z => n89);
   U110 : OAI21D1 port map( A1 => n96, A2 => n102, B => n97, Z => n95);
   U113 : NOR2D2 port map( A1 => A(5), A2 => B(5), Z => n96);
   U115 : EXNOR2D1 port map( A1 => n103, A2 => n15, Z => SUM(4));
   U116 : AOI21D1 port map( A1 => n103, A2 => n99, B => n100, Z => n98);
   U121 : NOR2D2 port map( A1 => A(4), A2 => B(4), Z => n101);
   U123 : EXNOR2D1 port map( A1 => n109, A2 => n16, Z => SUM(3));
   U130 : NOR2D2 port map( A1 => A(3), A2 => B(3), Z => n107);
   U132 : EXOR2D1 port map( A1 => n112, A2 => n17, Z => SUM(2));
   U138 : EXOR2D1 port map( A1 => n18, A2 => n117, Z => SUM(1));
   U140 : OAI21D1 port map( A1 => n114, A2 => n117, B => n115, Z => n113);
   U153 : OR2DL port map( A1 => A(0), A2 => B(0), Z => n189);
   U154 : NAN2D1 port map( A1 => A(6), A2 => B(6), Z => n88);
   U155 : NAN2D1 port map( A1 => A(8), A2 => B(8), Z => n74);
   U156 : NOR2D1 port map( A1 => A(2), A2 => B(2), Z => n110);
   U157 : NAN2D1 port map( A1 => A(4), A2 => B(4), Z => n102);
   U158 : NAN2DL port map( A1 => n86, A2 => n88, Z => n13);
   U159 : NAN2DL port map( A1 => n124, A2 => n69, Z => n10);
   U160 : NAN2DL port map( A1 => n126, A2 => n81, Z => n12);
   U161 : NAN2DL port map( A1 => n130, A2 => n108, Z => n16);
   U162 : NAN2DL port map( A1 => n128, A2 => n97, Z => n14);
   U163 : INVD1 port map( A => n94, Z => n92);
   U164 : NOR2D1 port map( A1 => n101, A2 => n96, Z => n94);
   U165 : NAN2M1DL port map( A1 => n38, A2 => n39, Z => n6);
   U166 : AOI21DL port map( A1 => n1, A2 => n48, B => n49, Z => n47);
   U167 : NAN2M1DL port map( A1 => n29, A2 => n30, Z => n5);
   U168 : AOI21DL port map( A1 => n1, A2 => n32, B => n33, Z => n31);
   U169 : INVDL port map( A => n3, Z => n48);
   U170 : INVDL port map( A => n65, Z => n63);
   U171 : INVDL port map( A => n64, Z => n62);
   U172 : NOR2DL port map( A1 => n3, A2 => n34, Z => n32);
   U173 : NOR2DL port map( A1 => n3, A2 => n25, Z => n23);
   U174 : NOR2DL port map( A1 => n64, A2 => n57, Z => n55);
   U175 : INVDL port map( A => n52, Z => n122);
   U176 : NAN2M1DL port map( A1 => n59, A2 => n60, Z => n9);
   U177 : NAN2M1DL port map( A1 => n45, A2 => n46, Z => n7);
   U178 : NAN2M1DL port map( A1 => n73, A2 => n74, Z => n11);
   U179 : AOI21D1 port map( A1 => n190, A2 => n113, B => n191, Z => n104);
   U180 : NOR2DL port map( A1 => n110, A2 => n107, Z => n190);
   U181 : OAI21DL port map( A1 => n107, A2 => n111, B => n108, Z => n191);
   U182 : INVD1 port map( A => n86, Z => n85);
   U183 : NAN2M1DL port map( A1 => n101, A2 => n102, Z => n15);
   U184 : INVDL port map( A => n73, Z => n71);
   U185 : NAN2M1DL port map( A1 => n110, A2 => n111, Z => n17);
   U186 : OA21M20DL port map( A1 => n37, A2 => n27, B => n30, Z => n26);
   U187 : NAN2M1DL port map( A1 => n114, A2 => n115, Z => n18);
   U188 : NOR2DL port map( A1 => n45, A2 => n38, Z => n36);
   U189 : OAI21DL port map( A1 => n112, A2 => n110, B => n111, Z => n109);
   U190 : INVDL port map( A => n29, Z => n27);
   U191 : NAN2D1 port map( A1 => A(7), A2 => B(7), Z => n81);
   U192 : NAN2D1 port map( A1 => A(5), A2 => B(5), Z => n97);
   U193 : NAN2D1 port map( A1 => A(9), A2 => B(9), Z => n69);
   U194 : NAN2D1 port map( A1 => A(10), A2 => B(10), Z => n60);
   U195 : NAN2D1 port map( A1 => A(3), A2 => B(3), Z => n108);
   U196 : NAN2DL port map( A1 => A(14), A2 => B(14), Z => n30);
   U197 : AND2DL port map( A1 => n189, A2 => n117, Z => SUM(0));
   U198 : INVDL port map( A => n2, Z => n49);
   U199 : INVD1 port map( A => n37, Z => n35);
   U200 : BUFD4 port map( A => n75, Z => n1);
   U201 : NAN2D1 port map( A1 => n94, A2 => n78, Z => n76);
   U202 : NAN2D1 port map( A1 => n66, A2 => n50, Z => n3);
   U203 : NOR2D1 port map( A1 => n3, A2 => n43, Z => n41);
   U204 : INVDL port map( A => n67, Z => n65);
   U205 : INVD1 port map( A => n66, Z => n64);
   U206 : INVDL port map( A => n95, Z => n93);
   U207 : NOR2D1 port map( A1 => n92, A2 => n85, Z => n83);
   U208 : INVD1 port map( A => n104, Z => n103);
   U209 : INVD1 port map( A => n36, Z => n34);
   U210 : NAN2D1 port map( A1 => n36, A2 => n27, Z => n25);
   U211 : INVD1 port map( A => n113, Z => n112);
   U212 : NOR2D1 port map( A1 => n87, A2 => n80, Z => n78);
   U213 : INVDL port map( A => n68, Z => n124);
   U214 : NOR2D1 port map( A1 => n73, A2 => n68, Z => n66);
   U215 : INVDL port map( A => n80, Z => n126);
   U216 : INVDL port map( A => n87, Z => n86);
   U217 : INVDL port map( A => n96, Z => n128);
   U218 : INVD1 port map( A => n58, Z => n57);
   U219 : INVDL port map( A => n59, Z => n58);
   U220 : INVD1 port map( A => n44, Z => n43);
   U221 : INVDL port map( A => n45, Z => n44);
   U222 : INVDL port map( A => n74, Z => n72);
   U223 : INVDL port map( A => n107, Z => n130);
   U224 : INVDL port map( A => n101, Z => n99);
   U225 : INVDL port map( A => n102, Z => n100);
   U226 : NOR2D1 port map( A1 => A(1), A2 => B(1), Z => n114);
   U227 : NOR2D1 port map( A1 => A(8), A2 => B(8), Z => n73);
   U228 : NAN2D1 port map( A1 => n193, A2 => n21, Z => n4);
   U229 : NAN2DL port map( A1 => A(15), A2 => B(15), Z => n21);
   U230 : NOR2D1 port map( A1 => A(11), A2 => B(11), Z => n52);
   U231 : NAN2DL port map( A1 => A(1), A2 => B(1), Z => n115);
   U232 : NAN2D1 port map( A1 => A(2), A2 => B(2), Z => n111);
   U233 : NAN2D1 port map( A1 => A(0), A2 => B(0), Z => n117);
   U234 : NOR2D1 port map( A1 => A(13), A2 => B(13), Z => n38);
   U235 : NAN2DL port map( A1 => A(12), A2 => B(12), Z => n46);
   U236 : NAN2DL port map( A1 => A(13), A2 => B(13), Z => n39);
   U237 : NOR2D1 port map( A1 => A(14), A2 => B(14), Z => n29);
   U238 : OR2D1 port map( A1 => A(15), A2 => B(15), Z => n193);
   U239 : NAN2DL port map( A1 => A(11), A2 => B(11), Z => n53);
   U240 : NAN2D1 port map( A1 => n122, A2 => n53, Z => n8);
   U241 : NOR2D1 port map( A1 => n59, A2 => n52, Z => n50);

end hier_sec_par_16_5;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_siso_gen.all;

architecture hier_sec_par_16_5 of siso_gen_DW_mult_tc_8 is

   component BUFD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22M10D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OA22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AO21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INVDL
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFD4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22DL
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21M20DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1DL
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AO21M20DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21DL
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFD20
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component ADHALFD1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component NOR2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n15, n16, n17, n18, 
      n19, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33, n34, n35, n36
      , n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n51, n52, n54, n55, 
      n56, n57, n58, n59, n60, n62, n63, n64, n65, n66, n67, n68, n69, n84, n85
      , n86, n87, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n112, n113, n114, n115, 
      n116, n117, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149, n150, n151, n152, n155, n156, n157, n158, n159, 
      n160, n161, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, 
      n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, 
      n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      n210, n213, n214, n215, n216, n217, n229, n230, n231, n232, n243, n248, 
      n249, n250, n261, n266, n267, n268, n269, n274, n275, n276, n277, n292, 
      n293, n294, n296, n297, n298, n315, n316, n317, n318, n319, n320, n321, 
      n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, 
      n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, 
      n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, 
      n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, 
      n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, 
      n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, 
      n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, 
      n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, 
      n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, 
      n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, 
      n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, 
      n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, 
      n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, 
      n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, 
      n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, 
      n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, 
      n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, 
      n526, n527, n528, n529, n530, n532, n533, n534, n535, n536, n537, n538, 
      n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, 
      n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, 
      n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, 
      n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, 
      n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, 
      n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, 
      n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, 
      n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, 
      n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, 
      n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, 
      n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, 
      n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, 
      n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, 
      n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, 
      n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, 
      n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, 
      n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, 
      n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, 
      n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, 
      n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, 
      n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, 
      n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, 
      n803, n805, n806, n807, n808, n809, n811, n812, n813, n814, n815, n816, 
      n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, 
      n829, n830, n831, n832, n833, n834, n837, n838, n839, n840, n842, n910, 
      n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, 
      n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, 
      n935, n936, n937, n938 : std_logic;

begin
   
   U54 : EXOR2D1 port map( A1 => n85, A2 => n54, Z => product(29));
   U59 : EXOR2D1 port map( A1 => n94, A2 => n55, Z => product(28));
   U60 : AOI21D1 port map( A1 => n51, A2 => n86, B => n87, Z => n85);
   U62 : OAI21D1 port map( A1 => n52, A2 => n918, B => n917, Z => n87);
   U71 : EXOR2D1 port map( A1 => n105, A2 => n56, Z => product(27));
   U74 : OAI21D1 port map( A1 => n52, A2 => n97, B => n100, Z => n96);
   U78 : AOI21D1 port map( A1 => n124, A2 => n101, B => n102, Z => n100);
   U80 : OAI21D1 port map( A1 => n113, A2 => n103, B => n104, Z => n102);
   U85 : EXOR2D1 port map( A1 => n114, A2 => n57, Z => product(26));
   U88 : OAI21D1 port map( A1 => n52, A2 => n108, B => n109, Z => n107);
   U97 : EXOR2D1 port map( A1 => n127, A2 => n58, Z => product(25));
   U108 : OAI21D1 port map( A1 => n133, A2 => n125, B => n126, Z => n124);
   U113 : EXOR2D1 port map( A1 => n134, A2 => n59, Z => product(24));
   U116 : OAI21D1 port map( A1 => n52, A2 => n130, B => n133, Z => n129);
   U121 : NOR2D2 port map( A1 => n332, A2 => n337, Z => n132);
   U123 : EXOR2D1 port map( A1 => n147, A2 => n60, Z => product(23));
   U128 : AOI21D1 port map( A1 => n173, A2 => n139, B => n140, Z => n138);
   U130 : OAI21D1 port map( A1 => n141, A2 => n166, B => n142, Z => n140);
   U132 : AOI21D1 port map( A1 => n155, A2 => n143, B => n144, Z => n142);
   U142 : OAI21D1 port map( A1 => n171, A2 => n150, B => n151, Z => n149);
   U144 : AOI21D1 port map( A1 => n164, A2 => n152, B => n155, Z => n151);
   U153 : EXOR2D1 port map( A1 => n167, A2 => n62, Z => product(21));
   U154 : AOI21D1 port map( A1 => n51, A2 => n159, B => n160, Z => n158);
   U163 : NOR2D2 port map( A1 => n354, A2 => n363, Z => n165);
   U165 : EXOR2D1 port map( A1 => n176, A2 => n63, Z => product(20));
   U172 : OAI21D1 port map( A1 => n174, A2 => n180, B => n175, Z => n173);
   U175 : NOR2D2 port map( A1 => n364, A2 => n373, Z => n174);
   U177 : EXNOR2D1 port map( A1 => n51, A2 => n64, Z => product(19));
   U178 : AOI21D1 port map( A1 => n51, A2 => n177, B => n178, Z => n176);
   U184 : NAN2D2 port map( A1 => n374, A2 => n385, Z => n180);
   U185 : EXOR2D1 port map( A1 => n188, A2 => n65, Z => product(18));
   U186 : OAI21D1 port map( A1 => n182, A2 => n210, B => n183, Z => n181);
   U188 : AOI21D1 port map( A1 => n201, A2 => n184, B => n185, Z => n183);
   U190 : OAI21D1 port map( A1 => n186, A2 => n194, B => n187, Z => n185);
   U193 : NOR2D2 port map( A1 => n386, A2 => n397, Z => n186);
   U195 : EXOR2D1 port map( A1 => n195, A2 => n66, Z => product(17));
   U196 : AOI21D1 port map( A1 => n189, A2 => n209, B => n190, Z => n188);
   U198 : OAI21D1 port map( A1 => n199, A2 => n191, B => n194, Z => n190);
   U203 : NOR2D2 port map( A1 => n398, A2 => n411, Z => n193);
   U205 : EXOR2D1 port map( A1 => n204, A2 => n67, Z => product(16));
   U206 : AOI21D1 port map( A1 => n209, A2 => n200, B => n197, Z => n195);
   U212 : OAI21D1 port map( A1 => n202, A2 => n208, B => n203, Z => n201);
   U215 : NOR2D2 port map( A1 => n412, A2 => n425, Z => n202);
   U217 : EXNOR2D1 port map( A1 => n209, A2 => n68, Z => product(15));
   U218 : AOI21D1 port map( A1 => n209, A2 => n205, B => n206, Z => n204);
   U223 : NOR2D2 port map( A1 => n426, A2 => n439, Z => n207);
   U225 : EXNOR2D1 port map( A1 => n215, A2 => n69, Z => product(14));
   U232 : NOR2D2 port map( A1 => n440, A2 => n451, Z => n213);
   U237 : AOI21D1 port map( A1 => n923, A2 => n910, B => n914, Z => n217);
   U256 : OAI21D1 port map( A1 => n243, A2 => n231, B => n232, Z => n230);
   U258 : AOI21D1 port map( A1 => n919, A2 => n921, B => n922, Z => n232);
   U275 : AOI21D1 port map( A1 => n248, A2 => n926, B => n929, Z => n243);
   U283 : OAI21D1 port map( A1 => n249, A2 => n261, B => n250, Z => n248);
   U302 : AOI21D1 port map( A1 => n266, A2 => n931, B => n932, Z => n261);
   U310 : OAI21D1 port map( A1 => n267, A2 => n269, B => n268, Z => n266);
   U316 : AOI21D1 port map( A1 => n274, A2 => n933, B => n934, Z => n269);
   U324 : OAI21D1 port map( A1 => n275, A2 => n277, B => n276, Z => n274);
   U330 : AOI21D1 port map( A1 => n935, A2 => n937, B => n936, Z => n277);
   U344 : ADFULD1 port map( A => n532, B => n319, CI => n547, CO => n315, S => 
                           n316);
   U345 : ADFULD1 port map( A => n320, B => n533, CI => n323, CO => n317, S => 
                           n318);
   U347 : ADFULD1 port map( A => n327, B => n563, CI => n324, CO => n321, S => 
                           n322);
   U348 : ADFULD1 port map( A => n548, B => n329, CI => n534, CO => n323, S => 
                           n324);
   U349 : ADFULD1 port map( A => n328, B => n335, CI => n333, CO => n325, S => 
                           n326);
   U350 : ADFULD1 port map( A => n535, B => n549, CI => n330, CO => n327, S => 
                           n328);
   U352 : ADFULD1 port map( A => n339, B => n336, CI => n334, CO => n331, S => 
                           n332);
   U353 : ADFULD1 port map( A => n579, B => n564, CI => n341, CO => n333, S => 
                           n334);
   U354 : ADFULD1 port map( A => n550, B => n536, CI => n343, CO => n335, S => 
                           n336);
   U355 : ADFULD1 port map( A => n347, B => n342, CI => n340, CO => n337, S => 
                           n338);
   U356 : ADFULD1 port map( A => n351, B => n344, CI => n349, CO => n339, S => 
                           n340);
   U357 : ADFULD1 port map( A => n551, B => n537, CI => n565, CO => n341, S => 
                           n342);
   U359 : ADFULD1 port map( A => n348, B => n357, CI => n355, CO => n345, S => 
                           n346);
   U360 : ADFULD1 port map( A => n352, B => n359, CI => n350, CO => n347, S => 
                           n348);
   U361 : ADFULD1 port map( A => n566, B => n552, CI => n595, CO => n349, S => 
                           n350);
   U362 : ADFULD1 port map( A => n580, B => n538, CI => n361, CO => n351, S => 
                           n352);
   U363 : ADFULD1 port map( A => n365, B => n358, CI => n356, CO => n353, S => 
                           n354);
   U364 : ADFULD1 port map( A => n360, B => n369, CI => n367, CO => n355, S => 
                           n356);
   U365 : ADFULD1 port map( A => n362, B => n567, CI => n371, CO => n357, S => 
                           n358);
   U366 : ADFULD1 port map( A => n581, B => n553, CI => n539, CO => n359, S => 
                           n360);
   U368 : ADFULD1 port map( A => n375, B => n368, CI => n366, CO => n363, S => 
                           n364);
   U369 : ADFULD1 port map( A => n372, B => n370, CI => n377, CO => n365, S => 
                           n366);
   U370 : ADFULD1 port map( A => n381, B => n611, CI => n379, CO => n367, S => 
                           n368);
   U371 : ADFULD1 port map( A => n554, B => n582, CI => n596, CO => n369, S => 
                           n370);
   U372 : ADFULD1 port map( A => n383, B => n540, CI => n568, CO => n371, S => 
                           n372);
   U373 : ADFULD1 port map( A => n387, B => n378, CI => n376, CO => n373, S => 
                           n374);
   U374 : ADFULD1 port map( A => n391, B => n380, CI => n389, CO => n375, S => 
                           n376);
   U375 : ADFULD1 port map( A => n393, B => n395, CI => n382, CO => n377, S => 
                           n378);
   U376 : ADFULD1 port map( A => n541, B => n555, CI => n384, CO => n379, S => 
                           n380);
   U377 : ADFULD1 port map( A => n597, B => n569, CI => n583, CO => n381, S => 
                           n382);
   U379 : ADFULD1 port map( A => n399, B => n390, CI => n388, CO => n385, S => 
                           n386);
   U380 : ADFULD1 port map( A => n392, B => n403, CI => n401, CO => n387, S => 
                           n388);
   U381 : ADFULD1 port map( A => n394, B => n405, CI => n396, CO => n389, S => 
                           n390);
   U382 : ADFULD1 port map( A => n627, B => n584, CI => n407, CO => n391, S => 
                           n392);
   U383 : ADFULD1 port map( A => n570, B => n598, CI => n612, CO => n393, S => 
                           n394);
   U384 : ADFULD1 port map( A => n409, B => n542, CI => n556, CO => n395, S => 
                           n396);
   U385 : ADFULD1 port map( A => n413, B => n402, CI => n400, CO => n397, S => 
                           n398);
   U386 : ADFULD1 port map( A => n404, B => n417, CI => n415, CO => n399, S => 
                           n400);
   U387 : ADFULD1 port map( A => n406, B => n419, CI => n408, CO => n401, S => 
                           n402);
   U388 : ADFULD1 port map( A => n423, B => n410, CI => n421, CO => n403, S => 
                           n404);
   U389 : ADFULD1 port map( A => n557, B => n599, CI => n585, CO => n405, S => 
                           n406);
   U390 : ADFULD1 port map( A => n543, B => n571, CI => n613, CO => n407, S => 
                           n408);
   U392 : ADFULD1 port map( A => n427, B => n416, CI => n414, CO => n411, S => 
                           n412);
   U393 : ADFULD1 port map( A => n429, B => n431, CI => n418, CO => n413, S => 
                           n414);
   U394 : ADFULD1 port map( A => n422, B => n433, CI => n420, CO => n415, S => 
                           n416);
   U395 : ADFULD1 port map( A => n424, B => n437, CI => n435, CO => n417, S => 
                           n418);
   U396 : ADFULD1 port map( A => n614, B => n628, CI => n643, CO => n419, S => 
                           n420);
   U397 : ADFULD1 port map( A => n544, B => n586, CI => n572, CO => n421, S => 
                           n422);
   U400 : ADFULD1 port map( A => n441, B => n430, CI => n428, CO => n425, S => 
                           n426);
   U401 : ADFULD1 port map( A => n443, B => n436, CI => n432, CO => n427, S => 
                           n428);
   U402 : ADFULD1 port map( A => n445, B => n447, CI => n434, CO => n429, S => 
                           n430);
   U403 : ADFULD1 port map( A => n438, B => n615, CI => n449, CO => n431, S => 
                           n432);
   U404 : ADFULD1 port map( A => n629, B => n573, CI => n601, CO => n433, S => 
                           n434);
   U405 : ADFULD1 port map( A => n545, B => n587, CI => n559, CO => n435, S => 
                           n436);
   U406 : ADHALFD1 port map( A => n523, B => n644, CO => n437, S => n438);
   U407 : ADFULD1 port map( A => n453, B => n444, CI => n442, CO => n439, S => 
                           n440);
   U408 : ADFULD1 port map( A => n446, B => n448, CI => n455, CO => n441, S => 
                           n442);
   U409 : ADFULD1 port map( A => n457, B => n459, CI => n450, CO => n443, S => 
                           n444);
   U410 : ADFULD1 port map( A => n588, B => n602, CI => n461, CO => n445, S => 
                           n446);
   U411 : ADFULD1 port map( A => n560, B => n616, CI => n574, CO => n447, S => 
                           n448);
   U412 : ADFULD1 port map( A => n645, B => n546, CI => n630, CO => n449, S => 
                           n450);
   U413 : ADFULD1 port map( A => n465, B => n456, CI => n454, CO => n451, S => 
                           n452);
   U414 : ADFULD1 port map( A => n460, B => n458, CI => n467, CO => n453, S => 
                           n454);
   U415 : ADFULD1 port map( A => n471, B => n462, CI => n469, CO => n455, S => 
                           n456);
   U416 : ADFULD1 port map( A => n561, B => n603, CI => n575, CO => n457, S => 
                           n458);
   U417 : ADFULD1 port map( A => n631, B => n589, CI => n617, CO => n459, S => 
                           n460);
   U418 : ADHALFD1 port map( A => n524, B => n646, CO => n461, S => n462);
   U419 : ADFULD1 port map( A => n468, B => n475, CI => n466, CO => n463, S => 
                           n464);
   U420 : ADFULD1 port map( A => n470, B => n472, CI => n477, CO => n465, S => 
                           n466);
   U421 : ADFULD1 port map( A => n481, B => n604, CI => n479, CO => n467, S => 
                           n468);
   U422 : ADFULD1 port map( A => n576, B => n618, CI => n590, CO => n469, S => 
                           n470);
   U423 : ADFULD1 port map( A => n647, B => n562, CI => n632, CO => n471, S => 
                           n472);
   U424 : ADFULD1 port map( A => n485, B => n478, CI => n476, CO => n473, S => 
                           n474);
   U425 : ADFULD1 port map( A => n487, B => n489, CI => n480, CO => n475, S => 
                           n476);
   U426 : ADFULD1 port map( A => n591, B => n619, CI => n482, CO => n477, S => 
                           n478);
   U427 : ADFULD1 port map( A => n577, B => n605, CI => n633, CO => n479, S => 
                           n480);
   U429 : ADFULD1 port map( A => n493, B => n488, CI => n486, CO => n483, S => 
                           n484);
   U430 : ADFULD1 port map( A => n495, B => n497, CI => n490, CO => n485, S => 
                           n486);
   U431 : ADFULD1 port map( A => n592, B => n620, CI => n606, CO => n487, S => 
                           n488);
   U432 : ADFULD1 port map( A => n649, B => n578, CI => n634, CO => n489, S => 
                           n490);
   U433 : ADFULD1 port map( A => n496, B => n501, CI => n494, CO => n491, S => 
                           n492);
   U434 : ADFULD1 port map( A => n498, B => n635, CI => n503, CO => n493, S => 
                           n494);
   U435 : ADFULD1 port map( A => n593, B => n607, CI => n621, CO => n495, S => 
                           n496);
   U437 : ADFULD1 port map( A => n504, B => n507, CI => n502, CO => n499, S => 
                           n500);
   U438 : ADFULD1 port map( A => n608, B => n622, CI => n509, CO => n501, S => 
                           n502);
   U439 : ADFULD1 port map( A => n651, B => n594, CI => n636, CO => n503, S => 
                           n504);
   U440 : ADFULD1 port map( A => n513, B => n510, CI => n508, CO => n505, S => 
                           n506);
   U441 : ADFULD1 port map( A => n609, B => n637, CI => n623, CO => n507, S => 
                           n508);
   U443 : ADFULD1 port map( A => n517, B => n624, CI => n514, CO => n511, S => 
                           n512);
   U444 : ADFULD1 port map( A => n653, B => n610, CI => n638, CO => n513, S => 
                           n514);
   U445 : ADFULD1 port map( A => n625, B => n639, CI => n518, CO => n515, S => 
                           n516);
   U447 : ADFULD1 port map( A => n655, B => n626, CI => n640, CO => n519, S => 
                           n520);
   U451 : OAI22D1 port map( A1 => n46, A2 => n660, B1 => n48, B2 => n661, Z => 
                           n532);
   U452 : OAI22D1 port map( A1 => n46, A2 => n661, B1 => n48, B2 => n662, Z => 
                           n533);
   U453 : OAI22D1 port map( A1 => n46, A2 => n662, B1 => n48, B2 => n663, Z => 
                           n534);
   U454 : OAI22D1 port map( A1 => n46, A2 => n663, B1 => n48, B2 => n664, Z => 
                           n535);
   U455 : OAI22D1 port map( A1 => n46, A2 => n664, B1 => n48, B2 => n665, Z => 
                           n536);
   U456 : OAI22D1 port map( A1 => n46, A2 => n665, B1 => n48, B2 => n666, Z => 
                           n537);
   U457 : OAI22D1 port map( A1 => n45, A2 => n666, B1 => n47, B2 => n667, Z => 
                           n538);
   U458 : OAI22D1 port map( A1 => n45, A2 => n667, B1 => n47, B2 => n668, Z => 
                           n539);
   U459 : OAI22D1 port map( A1 => n45, A2 => n668, B1 => n47, B2 => n669, Z => 
                           n540);
   U460 : OAI22D1 port map( A1 => n45, A2 => n669, B1 => n47, B2 => n670, Z => 
                           n541);
   U461 : OAI22D1 port map( A1 => n45, A2 => n670, B1 => n47, B2 => n671, Z => 
                           n542);
   U462 : OAI22D1 port map( A1 => n45, A2 => n671, B1 => n47, B2 => n672, Z => 
                           n543);
   U463 : OAI22D1 port map( A1 => n45, A2 => n672, B1 => n47, B2 => n673, Z => 
                           n544);
   U464 : OAI22D1 port map( A1 => n45, A2 => n673, B1 => n47, B2 => n674, Z => 
                           n545);
   U465 : NOR2M1D1 port map( A1 => b(0), A2 => n45, Z => n546);
   U466 : EXNOR2D1 port map( A1 => n43, A2 => n795, Z => n659);
   U467 : EXNOR2D1 port map( A1 => n43, A2 => n796, Z => n660);
   U468 : EXNOR2D1 port map( A1 => n43, A2 => n797, Z => n661);
   U469 : EXNOR2D1 port map( A1 => n43, A2 => n798, Z => n662);
   U470 : EXNOR2D1 port map( A1 => n43, A2 => n799, Z => n663);
   U471 : EXNOR2D1 port map( A1 => n43, A2 => n800, Z => n664);
   U472 : EXNOR2D1 port map( A1 => n43, A2 => n801, Z => n665);
   U473 : EXNOR2D1 port map( A1 => n43, A2 => n802, Z => n666);
   U474 : EXNOR2D1 port map( A1 => n43, A2 => n803, Z => n667);
   U475 : EXNOR2D1 port map( A1 => n43, A2 => b(6), Z => n668);
   U476 : EXNOR2D1 port map( A1 => n43, A2 => n805, Z => n669);
   U477 : EXNOR2D1 port map( A1 => n43, A2 => n806, Z => n670);
   U478 : EXNOR2D1 port map( A1 => n43, A2 => n807, Z => n671);
   U479 : EXNOR2D1 port map( A1 => n43, A2 => n808, Z => n672);
   U480 : EXNOR2D1 port map( A1 => n43, A2 => n809, Z => n673);
   U481 : EXNOR2D1 port map( A1 => n43, A2 => b(0), Z => n674);
   U482 : NAN2M1D1 port map( A1 => b(0), A2 => n43, Z => n675);
   U485 : OAI22D1 port map( A1 => n40, A2 => n676, B1 => n42, B2 => n677, Z => 
                           n319);
   U486 : OAI22D1 port map( A1 => n40, A2 => n677, B1 => n42, B2 => n678, Z => 
                           n548);
   U487 : OAI22D1 port map( A1 => n40, A2 => n678, B1 => n42, B2 => n679, Z => 
                           n549);
   U488 : OAI22D1 port map( A1 => n40, A2 => n679, B1 => n42, B2 => n680, Z => 
                           n550);
   U489 : OAI22D1 port map( A1 => n40, A2 => n680, B1 => n42, B2 => n681, Z => 
                           n551);
   U490 : OAI22D1 port map( A1 => n40, A2 => n681, B1 => n42, B2 => n682, Z => 
                           n552);
   U491 : OAI22D1 port map( A1 => n40, A2 => n682, B1 => n42, B2 => n683, Z => 
                           n553);
   U492 : OAI22D1 port map( A1 => n39, A2 => n683, B1 => n41, B2 => n684, Z => 
                           n554);
   U493 : OAI22D1 port map( A1 => n39, A2 => n684, B1 => n41, B2 => n685, Z => 
                           n555);
   U494 : OAI22D1 port map( A1 => n39, A2 => n685, B1 => n41, B2 => n686, Z => 
                           n556);
   U495 : OAI22D1 port map( A1 => n39, A2 => n686, B1 => n41, B2 => n687, Z => 
                           n557);
   U496 : OAI22D1 port map( A1 => n39, A2 => n687, B1 => n41, B2 => n688, Z => 
                           n558);
   U497 : OAI22D1 port map( A1 => n39, A2 => n688, B1 => n41, B2 => n689, Z => 
                           n559);
   U498 : OAI22D1 port map( A1 => n39, A2 => n689, B1 => n41, B2 => n690, Z => 
                           n560);
   U499 : OAI22D1 port map( A1 => n39, A2 => n690, B1 => n41, B2 => n691, Z => 
                           n561);
   U500 : NOR2M1D1 port map( A1 => b(0), A2 => n39, Z => n562);
   U501 : EXNOR2D1 port map( A1 => n37, A2 => n795, Z => n676);
   U502 : EXNOR2D1 port map( A1 => n37, A2 => n796, Z => n677);
   U503 : EXNOR2D1 port map( A1 => n37, A2 => n797, Z => n678);
   U504 : EXNOR2D1 port map( A1 => n37, A2 => n798, Z => n679);
   U505 : EXNOR2D1 port map( A1 => n37, A2 => n799, Z => n680);
   U506 : EXNOR2D1 port map( A1 => n37, A2 => n800, Z => n681);
   U507 : EXNOR2D1 port map( A1 => n37, A2 => n801, Z => n682);
   U508 : EXNOR2D1 port map( A1 => n37, A2 => n802, Z => n683);
   U509 : EXNOR2D1 port map( A1 => n37, A2 => n803, Z => n684);
   U510 : EXNOR2D1 port map( A1 => n37, A2 => b(6), Z => n685);
   U511 : EXNOR2D1 port map( A1 => n37, A2 => n805, Z => n686);
   U512 : EXNOR2D1 port map( A1 => n37, A2 => n806, Z => n687);
   U513 : EXNOR2D1 port map( A1 => n37, A2 => n807, Z => n688);
   U514 : EXNOR2D1 port map( A1 => n37, A2 => n808, Z => n689);
   U515 : EXNOR2D1 port map( A1 => n37, A2 => n809, Z => n690);
   U516 : EXNOR2D1 port map( A1 => n37, A2 => b(0), Z => n691);
   U517 : NAN2M1D1 port map( A1 => b(0), A2 => n37, Z => n692);
   U518 : OAI22D1 port map( A1 => n34, A2 => n709, B1 => n36, B2 => n837, Z => 
                           n525);
   U520 : OAI22D1 port map( A1 => n34, A2 => n693, B1 => n36, B2 => n694, Z => 
                           n329);
   U521 : OAI22D1 port map( A1 => n34, A2 => n694, B1 => n36, B2 => n695, Z => 
                           n564);
   U522 : OAI22D1 port map( A1 => n34, A2 => n695, B1 => n36, B2 => n696, Z => 
                           n565);
   U523 : OAI22D1 port map( A1 => n34, A2 => n696, B1 => n36, B2 => n697, Z => 
                           n566);
   U524 : OAI22D1 port map( A1 => n34, A2 => n697, B1 => n36, B2 => n698, Z => 
                           n567);
   U525 : OAI22D1 port map( A1 => n34, A2 => n698, B1 => n36, B2 => n699, Z => 
                           n568);
   U526 : OAI22D1 port map( A1 => n34, A2 => n699, B1 => n36, B2 => n700, Z => 
                           n569);
   U527 : OAI22D1 port map( A1 => n33, A2 => n700, B1 => n35, B2 => n701, Z => 
                           n570);
   U528 : OAI22D1 port map( A1 => n33, A2 => n701, B1 => n35, B2 => n702, Z => 
                           n571);
   U529 : OAI22D1 port map( A1 => n33, A2 => n702, B1 => n35, B2 => n703, Z => 
                           n572);
   U530 : OAI22D1 port map( A1 => n33, A2 => n703, B1 => n35, B2 => n704, Z => 
                           n573);
   U531 : OAI22D1 port map( A1 => n33, A2 => n704, B1 => n35, B2 => n705, Z => 
                           n574);
   U532 : OAI22D1 port map( A1 => n33, A2 => n705, B1 => n35, B2 => n706, Z => 
                           n575);
   U533 : OAI22D1 port map( A1 => n33, A2 => n706, B1 => n35, B2 => n707, Z => 
                           n576);
   U534 : OAI22D1 port map( A1 => n33, A2 => n707, B1 => n35, B2 => n708, Z => 
                           n577);
   U535 : NOR2M1D1 port map( A1 => b(0), A2 => n33, Z => n578);
   U536 : EXNOR2D1 port map( A1 => n31, A2 => n795, Z => n693);
   U537 : EXNOR2D1 port map( A1 => n31, A2 => n796, Z => n694);
   U538 : EXNOR2D1 port map( A1 => n31, A2 => n797, Z => n695);
   U539 : EXNOR2D1 port map( A1 => n31, A2 => n798, Z => n696);
   U540 : EXNOR2D1 port map( A1 => n31, A2 => n799, Z => n697);
   U541 : EXNOR2D1 port map( A1 => n31, A2 => n800, Z => n698);
   U542 : EXNOR2D1 port map( A1 => n31, A2 => n801, Z => n699);
   U543 : EXNOR2D1 port map( A1 => n31, A2 => n802, Z => n700);
   U544 : EXNOR2D1 port map( A1 => n31, A2 => n803, Z => n701);
   U545 : EXNOR2D1 port map( A1 => n31, A2 => b(6), Z => n702);
   U546 : EXNOR2D1 port map( A1 => n31, A2 => n805, Z => n703);
   U547 : EXNOR2D1 port map( A1 => n31, A2 => n806, Z => n704);
   U548 : EXNOR2D1 port map( A1 => n31, A2 => n807, Z => n705);
   U549 : EXNOR2D1 port map( A1 => n31, A2 => n808, Z => n706);
   U550 : EXNOR2D1 port map( A1 => n31, A2 => n809, Z => n707);
   U551 : EXNOR2D1 port map( A1 => n31, A2 => b(0), Z => n708);
   U552 : NAN2M1D1 port map( A1 => b(0), A2 => n31, Z => n709);
   U553 : OAI22D1 port map( A1 => n28, A2 => n726, B1 => n30, B2 => n838, Z => 
                           n526);
   U555 : OAI22D1 port map( A1 => n28, A2 => n710, B1 => n30, B2 => n711, Z => 
                           n343);
   U556 : OAI22D1 port map( A1 => n28, A2 => n711, B1 => n30, B2 => n712, Z => 
                           n580);
   U557 : OAI22D1 port map( A1 => n28, A2 => n712, B1 => n30, B2 => n713, Z => 
                           n581);
   U558 : OAI22D1 port map( A1 => n28, A2 => n713, B1 => n30, B2 => n714, Z => 
                           n582);
   U559 : OAI22D1 port map( A1 => n28, A2 => n714, B1 => n30, B2 => n715, Z => 
                           n583);
   U560 : OAI22D1 port map( A1 => n28, A2 => n715, B1 => n30, B2 => n716, Z => 
                           n584);
   U561 : OAI22D1 port map( A1 => n28, A2 => n716, B1 => n30, B2 => n717, Z => 
                           n585);
   U562 : OAI22D1 port map( A1 => n27, A2 => n717, B1 => n29, B2 => n718, Z => 
                           n586);
   U563 : OAI22D1 port map( A1 => n27, A2 => n718, B1 => n29, B2 => n719, Z => 
                           n587);
   U564 : OAI22D1 port map( A1 => n27, A2 => n719, B1 => n29, B2 => n720, Z => 
                           n588);
   U565 : OAI22D1 port map( A1 => n27, A2 => n720, B1 => n29, B2 => n721, Z => 
                           n589);
   U566 : OAI22D1 port map( A1 => n27, A2 => n721, B1 => n29, B2 => n722, Z => 
                           n590);
   U567 : OAI22D1 port map( A1 => n27, A2 => n722, B1 => n29, B2 => n723, Z => 
                           n591);
   U568 : OAI22D1 port map( A1 => n27, A2 => n723, B1 => n29, B2 => n724, Z => 
                           n592);
   U569 : OAI22D1 port map( A1 => n27, A2 => n724, B1 => n29, B2 => n725, Z => 
                           n593);
   U570 : NOR2M1D1 port map( A1 => b(0), A2 => n27, Z => n594);
   U571 : EXNOR2D1 port map( A1 => n25, A2 => n795, Z => n710);
   U572 : EXNOR2D1 port map( A1 => n25, A2 => n796, Z => n711);
   U573 : EXNOR2D1 port map( A1 => n25, A2 => n797, Z => n712);
   U574 : EXNOR2D1 port map( A1 => n25, A2 => n798, Z => n713);
   U575 : EXNOR2D1 port map( A1 => n25, A2 => n799, Z => n714);
   U576 : EXNOR2D1 port map( A1 => n25, A2 => n800, Z => n715);
   U577 : EXNOR2D1 port map( A1 => n25, A2 => n801, Z => n716);
   U578 : EXNOR2D1 port map( A1 => n25, A2 => n802, Z => n717);
   U579 : EXNOR2D1 port map( A1 => n25, A2 => n803, Z => n718);
   U580 : EXNOR2D1 port map( A1 => n25, A2 => b(6), Z => n719);
   U581 : EXNOR2D1 port map( A1 => n25, A2 => n805, Z => n720);
   U582 : EXNOR2D1 port map( A1 => n25, A2 => n806, Z => n721);
   U583 : EXNOR2D1 port map( A1 => n25, A2 => n807, Z => n722);
   U584 : EXNOR2D1 port map( A1 => n25, A2 => n808, Z => n723);
   U585 : EXNOR2D1 port map( A1 => n25, A2 => n809, Z => n724);
   U586 : EXNOR2D1 port map( A1 => n25, A2 => b(0), Z => n725);
   U587 : NAN2M1D1 port map( A1 => b(0), A2 => n25, Z => n726);
   U588 : OAI22D1 port map( A1 => n22, A2 => n743, B1 => n24, B2 => n839, Z => 
                           n527);
   U590 : OAI22D1 port map( A1 => n22, A2 => n727, B1 => n24, B2 => n728, Z => 
                           n361);
   U591 : OAI22D1 port map( A1 => n22, A2 => n728, B1 => n24, B2 => n729, Z => 
                           n596);
   U592 : OAI22D1 port map( A1 => n22, A2 => n729, B1 => n24, B2 => n730, Z => 
                           n597);
   U593 : OAI22D1 port map( A1 => n22, A2 => n730, B1 => n24, B2 => n731, Z => 
                           n598);
   U594 : OAI22D1 port map( A1 => n22, A2 => n731, B1 => n24, B2 => n732, Z => 
                           n599);
   U595 : OAI22D1 port map( A1 => n22, A2 => n732, B1 => n24, B2 => n733, Z => 
                           n600);
   U596 : OAI22D1 port map( A1 => n22, A2 => n733, B1 => n24, B2 => n734, Z => 
                           n601);
   U597 : OAI22D1 port map( A1 => n21, A2 => n734, B1 => n23, B2 => n735, Z => 
                           n602);
   U598 : OAI22D1 port map( A1 => n21, A2 => n735, B1 => n23, B2 => n736, Z => 
                           n603);
   U599 : OAI22D1 port map( A1 => n21, A2 => n736, B1 => n23, B2 => n737, Z => 
                           n604);
   U600 : OAI22D1 port map( A1 => n21, A2 => n737, B1 => n23, B2 => n738, Z => 
                           n605);
   U601 : OAI22D1 port map( A1 => n21, A2 => n738, B1 => n23, B2 => n739, Z => 
                           n606);
   U602 : OAI22D1 port map( A1 => n21, A2 => n739, B1 => n23, B2 => n740, Z => 
                           n607);
   U603 : OAI22D1 port map( A1 => n21, A2 => n740, B1 => n23, B2 => n741, Z => 
                           n608);
   U604 : OAI22D1 port map( A1 => n21, A2 => n741, B1 => n23, B2 => n742, Z => 
                           n609);
   U605 : NOR2M1D1 port map( A1 => b(0), A2 => n21, Z => n610);
   U606 : EXNOR2D1 port map( A1 => n19, A2 => n795, Z => n727);
   U607 : EXNOR2D1 port map( A1 => n19, A2 => n796, Z => n728);
   U608 : EXNOR2D1 port map( A1 => n19, A2 => n797, Z => n729);
   U609 : EXNOR2D1 port map( A1 => n19, A2 => n798, Z => n730);
   U610 : EXNOR2D1 port map( A1 => n19, A2 => n799, Z => n731);
   U611 : EXNOR2D1 port map( A1 => n19, A2 => n800, Z => n732);
   U612 : EXNOR2D1 port map( A1 => n19, A2 => n801, Z => n733);
   U613 : EXNOR2D1 port map( A1 => n19, A2 => n802, Z => n734);
   U614 : EXNOR2D1 port map( A1 => n19, A2 => n803, Z => n735);
   U615 : EXNOR2D1 port map( A1 => n19, A2 => b(6), Z => n736);
   U616 : EXNOR2D1 port map( A1 => n19, A2 => n805, Z => n737);
   U617 : EXNOR2D1 port map( A1 => n19, A2 => n806, Z => n738);
   U618 : EXNOR2D1 port map( A1 => n19, A2 => n807, Z => n739);
   U619 : EXNOR2D1 port map( A1 => n19, A2 => n808, Z => n740);
   U620 : EXNOR2D1 port map( A1 => n19, A2 => n809, Z => n741);
   U621 : EXNOR2D1 port map( A1 => n19, A2 => b(0), Z => n742);
   U622 : NAN2M1D1 port map( A1 => b(0), A2 => n19, Z => n743);
   U623 : OAI22D1 port map( A1 => n16, A2 => n760, B1 => n18, B2 => n840, Z => 
                           n528);
   U625 : OAI22D1 port map( A1 => n16, A2 => n744, B1 => n18, B2 => n745, Z => 
                           n383);
   U626 : OAI22D1 port map( A1 => n16, A2 => n745, B1 => n18, B2 => n746, Z => 
                           n612);
   U627 : OAI22D1 port map( A1 => n16, A2 => n746, B1 => n18, B2 => n747, Z => 
                           n613);
   U628 : OAI22D1 port map( A1 => n16, A2 => n747, B1 => n18, B2 => n748, Z => 
                           n614);
   U629 : OAI22D1 port map( A1 => n16, A2 => n748, B1 => n18, B2 => n749, Z => 
                           n615);
   U630 : OAI22D1 port map( A1 => n16, A2 => n749, B1 => n18, B2 => n750, Z => 
                           n616);
   U631 : OAI22D1 port map( A1 => n16, A2 => n750, B1 => n18, B2 => n751, Z => 
                           n617);
   U632 : OAI22D1 port map( A1 => n15, A2 => n751, B1 => n17, B2 => n752, Z => 
                           n618);
   U633 : OAI22D1 port map( A1 => n15, A2 => n752, B1 => n17, B2 => n753, Z => 
                           n619);
   U634 : OAI22D1 port map( A1 => n15, A2 => n753, B1 => n17, B2 => n754, Z => 
                           n620);
   U635 : OAI22D1 port map( A1 => n15, A2 => n754, B1 => n17, B2 => n755, Z => 
                           n621);
   U636 : OAI22D1 port map( A1 => n15, A2 => n755, B1 => n17, B2 => n756, Z => 
                           n622);
   U637 : OAI22D1 port map( A1 => n15, A2 => n756, B1 => n17, B2 => n757, Z => 
                           n623);
   U638 : OAI22D1 port map( A1 => n15, A2 => n757, B1 => n17, B2 => n758, Z => 
                           n624);
   U639 : OAI22D1 port map( A1 => n15, A2 => n758, B1 => n17, B2 => n759, Z => 
                           n625);
   U640 : NOR2M1D1 port map( A1 => b(0), A2 => n15, Z => n626);
   U641 : EXNOR2D1 port map( A1 => n13, A2 => n795, Z => n744);
   U642 : EXNOR2D1 port map( A1 => n13, A2 => n796, Z => n745);
   U643 : EXNOR2D1 port map( A1 => n13, A2 => n797, Z => n746);
   U644 : EXNOR2D1 port map( A1 => n13, A2 => n798, Z => n747);
   U645 : EXNOR2D1 port map( A1 => n13, A2 => n799, Z => n748);
   U646 : EXNOR2D1 port map( A1 => n13, A2 => n800, Z => n749);
   U647 : EXNOR2D1 port map( A1 => n13, A2 => n801, Z => n750);
   U648 : EXNOR2D1 port map( A1 => n13, A2 => n802, Z => n751);
   U649 : EXNOR2D1 port map( A1 => n13, A2 => n803, Z => n752);
   U650 : EXNOR2D1 port map( A1 => n13, A2 => b(6), Z => n753);
   U651 : EXNOR2D1 port map( A1 => n13, A2 => n805, Z => n754);
   U652 : EXNOR2D1 port map( A1 => n13, A2 => n806, Z => n755);
   U653 : EXNOR2D1 port map( A1 => n13, A2 => n807, Z => n756);
   U654 : EXNOR2D1 port map( A1 => n13, A2 => n808, Z => n757);
   U655 : EXNOR2D1 port map( A1 => n13, A2 => n809, Z => n758);
   U656 : EXNOR2D1 port map( A1 => n13, A2 => b(0), Z => n759);
   U657 : NAN2M1D1 port map( A1 => b(0), A2 => n13, Z => n760);
   U660 : OAI22D1 port map( A1 => n10, A2 => n761, B1 => n12, B2 => n762, Z => 
                           n409);
   U661 : OAI22D1 port map( A1 => n10, A2 => n762, B1 => n12, B2 => n763, Z => 
                           n628);
   U662 : OAI22D1 port map( A1 => n10, A2 => n763, B1 => n12, B2 => n764, Z => 
                           n629);
   U663 : OAI22D1 port map( A1 => n10, A2 => n764, B1 => n12, B2 => n765, Z => 
                           n630);
   U664 : OAI22D1 port map( A1 => n10, A2 => n765, B1 => n12, B2 => n766, Z => 
                           n631);
   U665 : OAI22D1 port map( A1 => n10, A2 => n766, B1 => n12, B2 => n767, Z => 
                           n632);
   U666 : OAI22D1 port map( A1 => n10, A2 => n767, B1 => n12, B2 => n768, Z => 
                           n633);
   U667 : OAI22D1 port map( A1 => n9, A2 => n768, B1 => n11, B2 => n769, Z => 
                           n634);
   U668 : OAI22D1 port map( A1 => n9, A2 => n769, B1 => n11, B2 => n770, Z => 
                           n635);
   U669 : OAI22D1 port map( A1 => n9, A2 => n770, B1 => n11, B2 => n771, Z => 
                           n636);
   U670 : OAI22D1 port map( A1 => n9, A2 => n771, B1 => n11, B2 => n772, Z => 
                           n637);
   U671 : OAI22D1 port map( A1 => n9, A2 => n772, B1 => n11, B2 => n773, Z => 
                           n638);
   U672 : OAI22D1 port map( A1 => n9, A2 => n773, B1 => n11, B2 => n774, Z => 
                           n639);
   U673 : OAI22D1 port map( A1 => n9, A2 => n774, B1 => n11, B2 => n775, Z => 
                           n640);
   U674 : OAI22D1 port map( A1 => n9, A2 => n775, B1 => n11, B2 => n776, Z => 
                           n641);
   U675 : NOR2M1D1 port map( A1 => b(0), A2 => n9, Z => n642);
   U676 : EXNOR2D1 port map( A1 => n7, A2 => n795, Z => n761);
   U677 : EXNOR2D1 port map( A1 => n7, A2 => n796, Z => n762);
   U678 : EXNOR2D1 port map( A1 => n7, A2 => n797, Z => n763);
   U679 : EXNOR2D1 port map( A1 => n7, A2 => n798, Z => n764);
   U680 : EXNOR2D1 port map( A1 => n7, A2 => n799, Z => n765);
   U681 : EXNOR2D1 port map( A1 => n7, A2 => n800, Z => n766);
   U682 : EXNOR2D1 port map( A1 => n7, A2 => n801, Z => n767);
   U683 : EXNOR2D1 port map( A1 => n7, A2 => n802, Z => n768);
   U684 : EXNOR2D1 port map( A1 => n7, A2 => n803, Z => n769);
   U685 : EXNOR2D1 port map( A1 => n7, A2 => b(6), Z => n770);
   U686 : EXNOR2D1 port map( A1 => n7, A2 => n805, Z => n771);
   U687 : EXNOR2D1 port map( A1 => n7, A2 => n806, Z => n772);
   U688 : EXNOR2D1 port map( A1 => n7, A2 => n807, Z => n773);
   U689 : EXNOR2D1 port map( A1 => n7, A2 => n808, Z => n774);
   U690 : EXNOR2D1 port map( A1 => n7, A2 => n809, Z => n775);
   U691 : EXNOR2D1 port map( A1 => n7, A2 => b(0), Z => n776);
   U692 : NAN2M1D1 port map( A1 => b(0), A2 => n7, Z => n777);
   U693 : OAI22D1 port map( A1 => n794, A2 => n4, B1 => n6, B2 => n842, Z => 
                           n530);
   U696 : OAI22D1 port map( A1 => n779, A2 => n4, B1 => n6, B2 => n780, Z => 
                           n645);
   U697 : OAI22D1 port map( A1 => n780, A2 => n4, B1 => n6, B2 => n781, Z => 
                           n646);
   U698 : OAI22D1 port map( A1 => n781, A2 => n4, B1 => n6, B2 => n782, Z => 
                           n647);
   U699 : OAI22D1 port map( A1 => n782, A2 => n4, B1 => n6, B2 => n783, Z => 
                           n648);
   U700 : OAI22D1 port map( A1 => n783, A2 => n4, B1 => n6, B2 => n784, Z => 
                           n649);
   U701 : OAI22D1 port map( A1 => n784, A2 => n4, B1 => n6, B2 => n785, Z => 
                           n650);
   U702 : OAI22D1 port map( A1 => n785, A2 => n3, B1 => n5, B2 => n786, Z => 
                           n651);
   U703 : OAI22D1 port map( A1 => n786, A2 => n3, B1 => n5, B2 => n787, Z => 
                           n652);
   U704 : OAI22D1 port map( A1 => n787, A2 => n3, B1 => n5, B2 => n788, Z => 
                           n653);
   U705 : OAI22D1 port map( A1 => n788, A2 => n3, B1 => n5, B2 => n789, Z => 
                           n654);
   U706 : OAI22D1 port map( A1 => n789, A2 => n3, B1 => n5, B2 => n790, Z => 
                           n655);
   U707 : OAI22D1 port map( A1 => n790, A2 => n3, B1 => n5, B2 => n791, Z => 
                           n656);
   U708 : OAI22D1 port map( A1 => n791, A2 => n3, B1 => n5, B2 => n792, Z => 
                           n657);
   U709 : OAI22D1 port map( A1 => n792, A2 => n3, B1 => n5, B2 => n793, Z => 
                           n658);
   U711 : EXNOR2D1 port map( A1 => n1, A2 => n795, Z => n778);
   U712 : EXNOR2D1 port map( A1 => n1, A2 => n796, Z => n779);
   U713 : EXNOR2D1 port map( A1 => n1, A2 => n797, Z => n780);
   U714 : EXNOR2D1 port map( A1 => n1, A2 => n798, Z => n781);
   U715 : EXNOR2D1 port map( A1 => n1, A2 => n799, Z => n782);
   U716 : EXNOR2D1 port map( A1 => n1, A2 => n800, Z => n783);
   U717 : EXNOR2D1 port map( A1 => n1, A2 => n801, Z => n784);
   U718 : EXNOR2D1 port map( A1 => n1, A2 => n802, Z => n785);
   U719 : EXNOR2D1 port map( A1 => n1, A2 => n803, Z => n786);
   U720 : EXNOR2D1 port map( A1 => n1, A2 => b(6), Z => n787);
   U721 : EXNOR2D1 port map( A1 => n1, A2 => n805, Z => n788);
   U722 : EXNOR2D1 port map( A1 => n1, A2 => n806, Z => n789);
   U723 : EXNOR2D1 port map( A1 => n1, A2 => n807, Z => n790);
   U724 : EXNOR2D1 port map( A1 => n1, A2 => n808, Z => n791);
   U725 : EXNOR2D1 port map( A1 => n1, A2 => n809, Z => n792);
   U726 : EXNOR2D1 port map( A1 => n1, A2 => b(0), Z => n793);
   U727 : NAN2M1D1 port map( A1 => b(0), A2 => n1, Z => n794);
   U752 : EXOR2D1 port map( A1 => a(14), A2 => a(15), Z => n811);
   U753 : EXNOR2D1 port map( A1 => a(14), A2 => a(13), Z => n827);
   U755 : EXOR2D1 port map( A1 => a(12), A2 => a(13), Z => n812);
   U756 : EXNOR2D1 port map( A1 => a(12), A2 => a(11), Z => n828);
   U758 : EXOR2D1 port map( A1 => a(10), A2 => a(11), Z => n813);
   U759 : EXNOR2D1 port map( A1 => a(10), A2 => a(9), Z => n829);
   U761 : EXOR2D1 port map( A1 => a(8), A2 => a(9), Z => n814);
   U762 : EXNOR2D1 port map( A1 => a(8), A2 => a(7), Z => n830);
   U764 : EXOR2D1 port map( A1 => a(6), A2 => a(7), Z => n815);
   U765 : EXNOR2D1 port map( A1 => a(6), A2 => a(5), Z => n831);
   U767 : EXOR2D1 port map( A1 => a(4), A2 => a(5), Z => n816);
   U768 : EXNOR2D1 port map( A1 => a(4), A2 => a(3), Z => n832);
   U770 : EXOR2D1 port map( A1 => a(2), A2 => a(3), Z => n817);
   U771 : EXNOR2D1 port map( A1 => a(2), A2 => a(1), Z => n833);
   U773 : EXOR2D1 port map( A1 => a(0), A2 => a(1), Z => n818);
   U777 : NAN2DL port map( A1 => n294, A2 => n175, Z => n63);
   U778 : NAN2DL port map( A1 => n293, A2 => n166, Z => n62);
   U779 : NAN2DL port map( A1 => n298, A2 => n203, Z => n67);
   U780 : NAN2DL port map( A1 => n297, A2 => n194, Z => n66);
   U781 : NAN2D1 port map( A1 => n813, A2 => n829, Z => n821);
   U782 : NAN2D1 port map( A1 => n817, A2 => n833, Z => n825);
   U783 : INVDL port map( A => n409, Z => n410);
   U784 : NAN2D1 port map( A1 => n815, A2 => n831, Z => n823);
   U785 : NAN2D1 port map( A1 => n816, A2 => n832, Z => n824);
   U786 : NAN2D1 port map( A1 => n814, A2 => n830, Z => n822);
   U787 : NOR2D1 port map( A1 => n338, A2 => n345, Z => n145);
   U788 : NAN2D1 port map( A1 => n812, A2 => n828, Z => n820);
   U789 : NAN2D1 port map( A1 => n811, A2 => n827, Z => n819);
   U790 : NAN2D1 port map( A1 => n426, A2 => n439, Z => n208);
   U791 : NOR2D1 port map( A1 => n193, A2 => n186, Z => n184);
   U792 : NAN2DL port map( A1 => n296, A2 => n187, Z => n65);
   U793 : NOR2D1 port map( A1 => n346, A2 => n353, Z => n156);
   U794 : INVDL port map( A => n156, Z => n292);
   U795 : AND2D1 port map( A1 => n464, A2 => n473, Z => n910);
   U796 : INVD1 port map( A => n200, Z => n198);
   U797 : NOR2D1 port map( A1 => n202, A2 => n207, Z => n200);
   U798 : BUFD20 port map( A => b(10), Z => n800);
   U799 : BUFD20 port map( A => b(9), Z => n801);
   U800 : BUFD20 port map( A => b(5), Z => n805);
   U801 : AND2D1 port map( A1 => n657, A2 => n642, Z => n936);
   U802 : OR2DL port map( A1 => n657, A2 => n642, Z => n935);
   U803 : INVDL port map( A => n172, Z => n170);
   U804 : INVDL port map( A => n112, Z => n110);
   U805 : NAN2DL port map( A1 => n172, A2 => n139, Z => n911);
   U806 : AOI21D1 port map( A1 => n51, A2 => n168, B => n169, Z => n167);
   U807 : AOI21DL port map( A1 => n51, A2 => n128, B => n129, Z => n127);
   U808 : AOI21DL port map( A1 => n51, A2 => n148, B => n149, Z => n147);
   U809 : AOI21DL port map( A1 => n51, A2 => n135, B => n136, Z => n134);
   U810 : NAN2D1 port map( A1 => n123, A2 => n110, Z => n108);
   U811 : NAN2D1 port map( A1 => n398, A2 => n411, Z => n194);
   U812 : AOI21DL port map( A1 => n51, A2 => n115, B => n116, Z => n114);
   U813 : AOI21DL port map( A1 => n51, A2 => n106, B => n107, Z => n105);
   U814 : OAI21DL port map( A1 => n229, A2 => n216, B => n217, Z => n215);
   U815 : AOI21DL port map( A1 => n51, A2 => n95, B => n96, Z => n94);
   U816 : AOI21D1 port map( A1 => n924, A2 => n927, B => n925, Z => n250);
   U817 : NAN2DL port map( A1 => n924, A2 => n928, Z => n249);
   U818 : OR2D1 port map( A1 => n512, A2 => n515, Z => n931);
   U819 : AND2DL port map( A1 => n512, A2 => n515, Z => n932);
   U820 : INVDL port map( A => n171, Z => n169);
   U821 : NOR2DL port map( A1 => n170, A2 => n150, Z => n148);
   U822 : NOR2DL port map( A1 => n911, A2 => n117, Z => n115);
   U823 : NOR2DL port map( A1 => n911, A2 => n97, Z => n95);
   U824 : NAN2M1DL port map( A1 => n179, A2 => n180, Z => n64);
   U825 : INVDL port map( A => n199, Z => n197);
   U826 : INVDL port map( A => n179, Z => n177);
   U827 : AO21M20DL port map( A1 => n171, A2 => n161, B => n164, Z => n160);
   U828 : AO21M20DL port map( A1 => n52, A2 => n117, B => n124, Z => n116);
   U829 : INVDL port map( A => n163, Z => n161);
   U830 : INVDL port map( A => n165, Z => n293);
   U831 : NAN2M1DL port map( A1 => n145, A2 => n146, Z => n60);
   U832 : NAN2M1DL port map( A1 => n132, A2 => n133, Z => n59);
   U833 : NAN2M1DL port map( A1 => n125, A2 => n126, Z => n58);
   U834 : BUFD1 port map( A => n138, Z => n52);
   U835 : INVD1 port map( A => n192, Z => n191);
   U836 : INVDL port map( A => n146, Z => n144);
   U837 : INVDL port map( A => n166, Z => n164);
   U838 : NOR2DL port map( A1 => n132, A2 => n125, Z => n123);
   U839 : NAN2DL port map( A1 => n123, A2 => n101, Z => n99);
   U840 : NAN2D1 port map( A1 => n412, A2 => n425, Z => n203);
   U841 : AOI21D1 port map( A1 => n912, A2 => n230, B => n913, Z => n210);
   U842 : NOR2DL port map( A1 => n216, A2 => n213, Z => n912);
   U843 : OAI21D1 port map( A1 => n217, A2 => n213, B => n214, Z => n913);
   U844 : NAN2D1 port map( A1 => n386, A2 => n397, Z => n187);
   U845 : NAN2D1 port map( A1 => n364, A2 => n373, Z => n175);
   U846 : NAN2M1DL port map( A1 => n207, A2 => n208, Z => n68);
   U847 : NAN2DL port map( A1 => n346, A2 => n353, Z => n157);
   U848 : NAN2M1DL port map( A1 => n112, A2 => n113, Z => n57);
   U849 : NAN2M1D1 port map( A1 => n103, A2 => n104, Z => n56);
   U850 : NAN2M1DL port map( A1 => n213, A2 => n214, Z => n69);
   U851 : OA21M20DL port map( A1 => n124, A2 => n110, B => n113, Z => n109);
   U852 : NAN2M1D1 port map( A1 => n92, A2 => n93, Z => n55);
   U853 : OR2DL port map( A1 => n99, A2 => n92, Z => n918);
   U854 : AND2DL port map( A1 => n452, A2 => n463, Z => n914);
   U855 : OR2DL port map( A1 => n600, A2 => n558, Z => n423);
   U856 : OR2D1 port map( A1 => n464, A2 => n473, Z => n915);
   U857 : NAN2DL port map( A1 => n919, A2 => n920, Z => n231);
   U858 : AND2D1 port map( A1 => n484, A2 => n491, Z => n921);
   U859 : NAN2DL port map( A1 => n325, A2 => n322, Z => n113);
   U860 : OR2DL port map( A1 => n506, A2 => n511, Z => n928);
   U861 : OAI22DL port map( A1 => n778, A2 => n4, B1 => n6, B2 => n779, Z => 
                           n644);
   U862 : NOR2D1 port map( A1 => n516, A2 => n519, Z => n267);
   U863 : NAN2DL port map( A1 => n522, A2 => n529, Z => n276);
   U864 : INVD1 port map( A => n911, Z => n135);
   U865 : NOR2D1 port map( A1 => n170, A2 => n161, Z => n159);
   U866 : INVD1 port map( A => n170, Z => n168);
   U867 : INVD1 port map( A => n123, Z => n117);
   U868 : INVD1 port map( A => n52, Z => n136);
   U869 : NAN2D1 port map( A1 => n292, A2 => n143, Z => n141);
   U870 : INVDL port map( A => n173, Z => n171);
   U871 : NOR2DL port map( A1 => n911, A2 => n130, Z => n128);
   U872 : NOR2D1 port map( A1 => n198, A2 => n191, Z => n189);
   U873 : NAN2D1 port map( A1 => n163, A2 => n152, Z => n150);
   U874 : INVD1 port map( A => n156, Z => n152);
   U875 : NOR2DL port map( A1 => n911, A2 => n108, Z => n106);
   U876 : INVDL port map( A => n180, Z => n178);
   U877 : INVD1 port map( A => n98, Z => n97);
   U878 : INVD1 port map( A => n99, Z => n98);
   U879 : BUFD4 port map( A => n181, Z => n51);
   U880 : NAN2DL port map( A1 => n200, A2 => n184, Z => n182);
   U881 : EXNOR2D1 port map( A1 => n158, A2 => n916, Z => product(22));
   U882 : AND2D1 port map( A1 => n292, A2 => n157, Z => n916);
   U883 : INVDL port map( A => n174, Z => n294);
   U884 : INVD1 port map( A => n210, Z => n209);
   U885 : INVDL port map( A => n193, Z => n297);
   U886 : INVDL port map( A => n202, Z => n298);
   U887 : INVDL port map( A => n186, Z => n296);
   U888 : NOR2D1 port map( A1 => n141, A2 => n165, Z => n139);
   U889 : NOR2D1 port map( A1 => n374, A2 => n385, Z => n179);
   U890 : NOR2D1 port map( A1 => n179, A2 => n174, Z => n172);
   U891 : INVD1 port map( A => n145, Z => n143);
   U892 : INVDL port map( A => n201, Z => n199);
   U893 : INVD1 port map( A => n157, Z => n155);
   U894 : INVDL port map( A => n165, Z => n163);
   U895 : INVDL port map( A => n193, Z => n192);
   U896 : INVD1 port map( A => n131, Z => n130);
   U897 : INVDL port map( A => n132, Z => n131);
   U898 : NOR2DL port map( A1 => n911, A2 => n918, Z => n86);
   U899 : INVDL port map( A => n230, Z => n229);
   U900 : NAN2D1 port map( A1 => n354, A2 => n363, Z => n166);
   U901 : NAN2D1 port map( A1 => n338, A2 => n345, Z => n146);
   U902 : INVDL port map( A => n207, Z => n205);
   U903 : INVDL port map( A => n208, Z => n206);
   U904 : OA21DL port map( A1 => n100, A2 => n92, B => n93, Z => n917);
   U905 : NAN2DL port map( A1 => n332, A2 => n337, Z => n133);
   U906 : NOR2D1 port map( A1 => n326, A2 => n331, Z => n125);
   U907 : NAN2DL port map( A1 => n326, A2 => n331, Z => n126);
   U908 : NOR2D1 port map( A1 => n112, A2 => n103, Z => n101);
   U909 : OR2D1 port map( A1 => n474, A2 => n483, Z => n919);
   U910 : OR2D1 port map( A1 => n484, A2 => n491, Z => n920);
   U911 : AND2DL port map( A1 => n474, A2 => n483, Z => n922);
   U912 : OR2D1 port map( A1 => n452, A2 => n463, Z => n923);
   U913 : NAN2D1 port map( A1 => n923, A2 => n915, Z => n216);
   U914 : NAN2DL port map( A1 => n440, A2 => n451, Z => n214);
   U915 : INVDL port map( A => n343, Z => n344);
   U916 : NOR2D1 port map( A1 => n325, A2 => n322, Z => n112);
   U917 : NOR2D1 port map( A1 => n318, A2 => n321, Z => n103);
   U918 : NAN2DL port map( A1 => n318, A2 => n321, Z => n104);
   U919 : NOR2D1 port map( A1 => n317, A2 => n316, Z => n92);
   U920 : NAN2D1 port map( A1 => n317, A2 => n316, Z => n93);
   U921 : OR2D1 port map( A1 => n500, A2 => n505, Z => n924);
   U922 : AND2DL port map( A1 => n500, A2 => n505, Z => n925);
   U923 : OR2D1 port map( A1 => n492, A2 => n499, Z => n926);
   U924 : AND2D1 port map( A1 => n506, A2 => n511, Z => n927);
   U925 : AND2DL port map( A1 => n492, A2 => n499, Z => n929);
   U926 : EXNOR2D1 port map( A1 => n600, A2 => n558, Z => n424);
   U927 : INVDL port map( A => n383, Z => n384);
   U928 : AO21D1 port map( A1 => n12, A2 => n10, B => n761, Z => n627);
   U929 : AO21D1 port map( A1 => n6, A2 => n4, B => n778, Z => n643);
   U930 : AO21D1 port map( A1 => n18, A2 => n16, B => n744, Z => n611);
   U931 : AO21D1 port map( A1 => n24, A2 => n22, B => n727, Z => n595);
   U932 : INVDL port map( A => n361, Z => n362);
   U933 : NAN2D1 port map( A1 => n930, A2 => n84, Z => n54);
   U934 : NAN2D1 port map( A1 => n315, A2 => n938, Z => n84);
   U935 : AO21D1 port map( A1 => n30, A2 => n28, B => n710, Z => n579);
   U936 : INVDL port map( A => n329, Z => n330);
   U937 : AO21D1 port map( A1 => n36, A2 => n34, B => n693, Z => n563);
   U938 : INVD1 port map( A => n319, Z => n320);
   U939 : AO21D1 port map( A1 => n42, A2 => n40, B => n676, Z => n547);
   U940 : OR2D1 port map( A1 => n315, A2 => n938, Z => n930);
   U941 : ADHALFDL port map( A => n527, B => n652, CO => n509, S => n510);
   U942 : INVD1 port map( A => n19, Z => n839);
   U943 : ADHALFDL port map( A => n526, B => n650, CO => n497, S => n498);
   U944 : INVD1 port map( A => n25, Z => n838);
   U945 : ADHALFDL port map( A => n525, B => n648, CO => n481, S => n482);
   U946 : INVD1 port map( A => n31, Z => n837);
   U947 : NAN2DL port map( A1 => n516, A2 => n519, Z => n268);
   U948 : OR2D1 port map( A1 => n520, A2 => n521, Z => n933);
   U949 : OAI22M10D1 port map( A1 => n43, A2 => n48, B1 => n46, B2 => n675, Z 
                           => n523);
   U950 : AND2DL port map( A1 => n520, A2 => n521, Z => n934);
   U951 : ADHALFDL port map( A => n528, B => n654, CO => n517, S => n518);
   U952 : INVD1 port map( A => n13, Z => n840);
   U953 : OAI22M10D1 port map( A1 => n37, A2 => n42, B1 => n40, B2 => n692, Z 
                           => n524);
   U954 : NOR2D1 port map( A1 => n522, A2 => n529, Z => n275);
   U955 : AND2D1 port map( A1 => n658, A2 => n530, Z => n937);
   U956 : BUFD1 port map( A => n823, Z => n23);
   U957 : BUFD1 port map( A => n821, Z => n35);
   U958 : BUFD1 port map( A => n824, Z => n17);
   U959 : BUFD1 port map( A => n825, Z => n12);
   U960 : BUFD1 port map( A => n822, Z => n29);
   U961 : BUFD1 port map( A => n823, Z => n24);
   U962 : BUFD1 port map( A => n822, Z => n30);
   U963 : BUFD1 port map( A => n825, Z => n11);
   U964 : BUFD1 port map( A => n821, Z => n36);
   U965 : BUFD1 port map( A => n820, Z => n41);
   U966 : BUFD1 port map( A => n819, Z => n48);
   U967 : BUFD1 port map( A => n820, Z => n42);
   U968 : BUFD1 port map( A => n824, Z => n18);
   U969 : BUFD1 port map( A => n831, Z => n21);
   U970 : BUFD1 port map( A => n829, Z => n33);
   U971 : BUFD1 port map( A => n832, Z => n15);
   U972 : BUFD1 port map( A => n830, Z => n27);
   U973 : BUFD1 port map( A => n831, Z => n22);
   U974 : BUFD1 port map( A => n833, Z => n10);
   U975 : BUFD1 port map( A => n819, Z => n47);
   U976 : BUFD1 port map( A => n833, Z => n9);
   U977 : BUFD1 port map( A => n830, Z => n28);
   U978 : BUFD1 port map( A => n829, Z => n34);
   U979 : BUFD1 port map( A => n828, Z => n39);
   U980 : BUFD1 port map( A => n826, Z => n6);
   U981 : BUFD1 port map( A => n827, Z => n45);
   U982 : BUFD1 port map( A => n826, Z => n5);
   U983 : BUFD1 port map( A => n828, Z => n40);
   U984 : BUFD1 port map( A => n827, Z => n46);
   U985 : BUFD1 port map( A => n832, Z => n16);
   U986 : BUFD1 port map( A => n834, Z => n4);
   U987 : BUFD1 port map( A => n834, Z => n3);
   U988 : INVD1 port map( A => n1, Z => n842);
   U989 : OA22D1 port map( A1 => n46, A2 => n659, B1 => n48, B2 => n660, Z => 
                           n938);
   U990 : BUFD1 port map( A => b(1), Z => n809);
   U991 : BUFD1 port map( A => b(4), Z => n806);
   U992 : BUFD1 port map( A => b(8), Z => n802);
   U993 : BUFD1 port map( A => b(2), Z => n808);
   U994 : BUFD1 port map( A => b(7), Z => n803);
   U995 : BUFD1 port map( A => b(3), Z => n807);
   U996 : BUFD1 port map( A => b(11), Z => n799);
   U997 : BUFD1 port map( A => b(14), Z => n796);
   U998 : BUFD1 port map( A => b(13), Z => n797);
   U999 : BUFD1 port map( A => b(12), Z => n798);
   U1000 : BUFD1 port map( A => b(15), Z => n795);
   U1001 : ADHALFDL port map( A => n641, B => n656, CO => n521, S => n522);
   U1002 : OAI22M10D1 port map( A1 => n7, A2 => n12, B1 => n10, B2 => n777, Z 
                           => n529);
   U1003 : NAN2D1 port map( A1 => n818, A2 => n834, Z => n826);
   U1004 : INVD1 port map( A => a(0), Z => n834);
   U1005 : BUFD1 port map( A => a(7), Z => n19);
   U1006 : BUFD1 port map( A => a(11), Z => n31);
   U1007 : BUFD1 port map( A => a(5), Z => n13);
   U1008 : BUFD1 port map( A => a(9), Z => n25);
   U1009 : BUFD1 port map( A => a(1), Z => n1);
   U1010 : BUFD1 port map( A => a(3), Z => n7);
   U1011 : BUFD1 port map( A => a(13), Z => n37);
   U1012 : BUFD1 port map( A => a(15), Z => n43);

end hier_sec_par_16_5;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_siso_gen.all;

architecture hier_sec_par_16_5 of siso_gen is

   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFDL
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFD4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component TIELO
      port( Z : out std_logic);
   end component;
   
   component TIEHI
      port( Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFD8
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INVBD4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFERPQ1
      port( D, CEB, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component DFERPQ4
      port( D, CEB, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component DFERPQL
      port( D, CEB, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component DFERPQ2
      port( D, CEB, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFRPQ1
      port( D, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component siso_gen_DW_mult_tc_18
      port( a, b : in std_logic_vector (15 downto 0);  product : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component siso_gen_DW_mult_tc_17
      port( a, b : in std_logic_vector (15 downto 0);  product : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component siso_gen_DW01_add_12
      port( A, B : in std_logic_vector (15 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (15 downto 0);  CO : out std_logic);
   end component;
   
   component siso_gen_DW01_add_11
      port( A, B : in std_logic_vector (15 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (15 downto 0);  CO : out std_logic);
   end component;
   
   component siso_gen_DW01_add_13
      port( A, B : in std_logic_vector (15 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (15 downto 0);  CO : out std_logic);
   end component;
   
   component siso_gen_DW_mult_tc_10
      port( a, b : in std_logic_vector (15 downto 0);  product : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component siso_gen_DW01_add_7
      port( A, B : in std_logic_vector (15 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (15 downto 0);  CO : out std_logic);
   end component;
   
   component siso_gen_DW_mult_tc_8
      port( a, b : in std_logic_vector (15 downto 0);  product : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component siso_gen_DW_mult_tc_9
      port( a, b : in std_logic_vector (15 downto 0);  product : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal ready_port, coeff_memory_79_port, coeff_memory_78_port, 
      coeff_memory_77_port, coeff_memory_76_port, coeff_memory_75_port, 
      coeff_memory_74_port, coeff_memory_73_port, coeff_memory_72_port, 
      coeff_memory_71_port, coeff_memory_70_port, coeff_memory_69_port, 
      coeff_memory_68_port, coeff_memory_67_port, coeff_memory_66_port, 
      coeff_memory_65_port, coeff_memory_64_port, coeff_memory_63_port, 
      coeff_memory_62_port, coeff_memory_61_port, coeff_memory_60_port, 
      coeff_memory_59_port, coeff_memory_58_port, coeff_memory_57_port, 
      coeff_memory_56_port, coeff_memory_55_port, coeff_memory_54_port, 
      coeff_memory_53_port, coeff_memory_52_port, coeff_memory_51_port, 
      coeff_memory_50_port, coeff_memory_49_port, coeff_memory_48_port, 
      coeff_memory_47_port, coeff_memory_46_port, coeff_memory_45_port, 
      coeff_memory_44_port, coeff_memory_43_port, coeff_memory_42_port, 
      coeff_memory_41_port, coeff_memory_40_port, coeff_memory_39_port, 
      coeff_memory_38_port, coeff_memory_37_port, coeff_memory_36_port, 
      coeff_memory_35_port, coeff_memory_34_port, coeff_memory_33_port, 
      coeff_memory_32_port, coeff_memory_31_port, coeff_memory_30_port, 
      coeff_memory_29_port, coeff_memory_28_port, coeff_memory_27_port, 
      coeff_memory_26_port, coeff_memory_25_port, coeff_memory_24_port, 
      coeff_memory_23_port, coeff_memory_22_port, coeff_memory_21_port, 
      coeff_memory_20_port, coeff_memory_19_port, coeff_memory_18_port, 
      coeff_memory_17_port, coeff_memory_16_port, coeff_memory_15_port, 
      coeff_memory_14_port, coeff_memory_13_port, coeff_memory_12_port, 
      coeff_memory_11_port, coeff_memory_10_port, coeff_memory_9_port, 
      coeff_memory_8_port, coeff_memory_7_port, coeff_memory_6_port, 
      coeff_memory_5_port, coeff_memory_4_port, coeff_memory_3_port, 
      coeff_memory_2_port, coeff_memory_1_port, coeff_memory_0_port, 
      coeff_counter_2_port, coeff_counter_1_port, coeff_counter_0_port, 
      z1_15_port, z1_14_port, z1_13_port, z1_12_port, z1_11_port, z1_10_port, 
      z1_9_port, z1_8_port, z1_7_port, z1_6_port, z1_5_port, z1_4_port, 
      z1_3_port, z1_2_port, z1_1_port, z1_0_port, z2_15_port, z2_14_port, 
      z2_13_port, z2_12_port, z2_11_port, z2_10_port, z2_9_port, z2_8_port, 
      z2_7_port, z2_6_port, z2_5_port, z2_4_port, z2_3_port, z2_2_port, 
      z2_1_port, z2_0_port, z1_next_15_port, z1_next_14_port, z1_next_13_port, 
      z1_next_12_port, z1_next_11_port, z1_next_10_port, z1_next_9_port, 
      z1_next_8_port, z1_next_7_port, z1_next_6_port, z1_next_5_port, 
      z1_next_4_port, z1_next_3_port, z1_next_2_port, z1_next_1_port, 
      z1_next_0_port, z2_next_15_port, z2_next_14_port, z2_next_13_port, 
      z2_next_12_port, z2_next_11_port, z2_next_10_port, z2_next_9_port, 
      z2_next_8_port, z2_next_7_port, z2_next_6_port, z2_next_5_port, 
      z2_next_4_port, z2_next_3_port, z2_next_2_port, z2_next_1_port, 
      z2_next_0_port, y_15_port, y_14_port, y_13_port, y_12_port, y_11_port, 
      y_10_port, y_9_port, y_8_port, y_7_port, y_6_port, y_5_port, y_4_port, 
      y_3_port, y_2_port, y_1_port, y_0_port, n22, n23, n25, n26, n27, n28, n29
      , n30, n31, n32, z2_temp_9_port, z2_temp_8_port, z2_temp_7_port, 
      z2_temp_6_port, z2_temp_5_port, z2_temp_4_port, z2_temp_3_port, 
      z2_temp_2_port, z2_temp_1_port, z2_temp_15_port, z2_temp_14_port, 
      z2_temp_13_port, z2_temp_12_port, z2_temp_11_port, z2_temp_10_port, 
      z2_temp_0_port, m3_9_port, m3_8_port, m3_7_port, m3_6_port, m3_5_port, 
      m3_4_port, m3_3_port, m3_2_port, m3_1_port, m3_15_port, m3_14_port, 
      m3_13_port, m3_12_port, m3_11_port, m3_10_port, m3_0_port, m2_9_port, 
      m2_8_port, m2_7_port, m2_6_port, m2_5_port, m2_4_port, m2_3_port, 
      m2_2_port, m2_1_port, m2_15_port, m2_14_port, m2_13_port, m2_12_port, 
      m2_11_port, m2_10_port, m2_0_port, m5_9_port, m5_8_port, m5_7_port, 
      m5_6_port, m5_5_port, m5_4_port, m5_3_port, m5_2_port, m5_1_port, 
      m5_15_port, m5_14_port, m5_13_port, m5_12_port, m5_11_port, m5_10_port, 
      m5_0_port, m4_9_port, m4_8_port, m4_7_port, m4_6_port, m4_5_port, 
      m4_4_port, m4_3_port, m4_2_port, m4_1_port, m4_15_port, m4_14_port, 
      m4_13_port, m4_12_port, m4_11_port, m4_10_port, m4_0_port, m1_9_port, 
      m1_8_port, m1_7_port, m1_6_port, m1_5_port, m1_4_port, m1_3_port, 
      m1_2_port, m1_1_port, m1_15_port, m1_14_port, m1_13_port, m1_12_port, 
      m1_11_port, m1_10_port, m1_0_port, n33, n34, n35, n36, n37, n38, n39, n40
      , n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, 
      n55, n56, n57, n58, n59, n60, n61, n_1091, n_1092, n_1093, n_1094, n_1095
      , n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104,
      n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, 
      n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, 
      n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, 
      n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, 
      n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, 
      n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, 
      n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, 
      n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174 : std_logic;

begin
   ready <= ready_port;
   
   mult_28_C94 : siso_gen_DW_mult_tc_9 port map( a(15) => coeff_memory_47_port,
                           a(14) => coeff_memory_46_port, a(13) => 
                           coeff_memory_45_port, a(12) => coeff_memory_44_port,
                           a(11) => coeff_memory_43_port, a(10) => 
                           coeff_memory_42_port, a(9) => coeff_memory_41_port, 
                           a(8) => coeff_memory_40_port, a(7) => 
                           coeff_memory_39_port, a(6) => coeff_memory_38_port, 
                           a(5) => coeff_memory_37_port, a(4) => 
                           coeff_memory_36_port, a(3) => coeff_memory_35_port, 
                           a(2) => coeff_memory_34_port, a(1) => 
                           coeff_memory_33_port, a(0) => coeff_memory_32_port, 
                           b(15) => data_in(15), b(14) => data_in(14), b(13) =>
                           data_in(13), b(12) => data_in(12), b(11) => 
                           data_in(11), b(10) => data_in(10), b(9) => 
                           data_in(9), b(8) => data_in(8), b(7) => data_in(7), 
                           b(6) => data_in(6), b(5) => data_in(5), b(4) => 
                           data_in(4), b(3) => data_in(3), b(2) => data_in(2), 
                           b(1) => data_in(1), b(0) => data_in(0), product(31) 
                           => n_1091, product(30) => n_1092, product(29) => 
                           m4_15_port, product(28) => m4_14_port, product(27) 
                           => m4_13_port, product(26) => m4_12_port, 
                           product(25) => m4_11_port, product(24) => m4_10_port
                           , product(23) => m4_9_port, product(22) => m4_8_port
                           , product(21) => m4_7_port, product(20) => m4_6_port
                           , product(19) => m4_5_port, product(18) => m4_4_port
                           , product(17) => m4_3_port, product(16) => m4_2_port
                           , product(15) => m4_1_port, product(14) => m4_0_port
                           , product(13) => n_1093, product(12) => n_1094, 
                           product(11) => n_1095, product(10) => n_1096, 
                           product(9) => n_1097, product(8) => n_1098, 
                           product(7) => n_1099, product(6) => n_1100, 
                           product(5) => n_1101, product(4) => n_1102, 
                           product(3) => n_1103, product(2) => n_1104, 
                           product(1) => n_1105, product(0) => n_1106);
   mult_28_C93 : siso_gen_DW_mult_tc_8 port map( a(15) => coeff_memory_63_port,
                           a(14) => coeff_memory_62_port, a(13) => 
                           coeff_memory_61_port, a(12) => coeff_memory_60_port,
                           a(11) => coeff_memory_59_port, a(10) => 
                           coeff_memory_58_port, a(9) => coeff_memory_57_port, 
                           a(8) => coeff_memory_56_port, a(7) => 
                           coeff_memory_55_port, a(6) => coeff_memory_54_port, 
                           a(5) => coeff_memory_53_port, a(4) => 
                           coeff_memory_52_port, a(3) => coeff_memory_51_port, 
                           a(2) => coeff_memory_50_port, a(1) => 
                           coeff_memory_49_port, a(0) => coeff_memory_48_port, 
                           b(15) => data_in(15), b(14) => data_in(14), b(13) =>
                           data_in(13), b(12) => data_in(12), b(11) => 
                           data_in(11), b(10) => data_in(10), b(9) => 
                           data_in(9), b(8) => data_in(8), b(7) => data_in(7), 
                           b(6) => data_in(6), b(5) => data_in(5), b(4) => 
                           data_in(4), b(3) => data_in(3), b(2) => data_in(2), 
                           b(1) => data_in(1), b(0) => data_in(0), product(31) 
                           => n_1107, product(30) => n_1108, product(29) => 
                           m2_15_port, product(28) => m2_14_port, product(27) 
                           => m2_13_port, product(26) => m2_12_port, 
                           product(25) => m2_11_port, product(24) => m2_10_port
                           , product(23) => m2_9_port, product(22) => m2_8_port
                           , product(21) => m2_7_port, product(20) => m2_6_port
                           , product(19) => m2_5_port, product(18) => m2_4_port
                           , product(17) => m2_3_port, product(16) => m2_2_port
                           , product(15) => m2_1_port, product(14) => m2_0_port
                           , product(13) => n_1109, product(12) => n_1110, 
                           product(11) => n_1111, product(10) => n_1112, 
                           product(9) => n_1113, product(8) => n_1114, 
                           product(7) => n_1115, product(6) => n_1116, 
                           product(5) => n_1117, product(4) => n_1118, 
                           product(3) => n_1119, product(2) => n_1120, 
                           product(1) => n_1121, product(0) => n_1122);
   add_1_root_add_0_root_add_101 : siso_gen_DW01_add_7 port map( A(15) => 
                           z1_15_port, A(14) => z1_14_port, A(13) => z1_13_port
                           , A(12) => z1_12_port, A(11) => z1_11_port, A(10) =>
                           z1_10_port, A(9) => z1_9_port, A(8) => z1_8_port, 
                           A(7) => z1_7_port, A(6) => z1_6_port, A(5) => 
                           z1_5_port, A(4) => z1_4_port, A(3) => z1_3_port, 
                           A(2) => z1_2_port, A(1) => z1_1_port, A(0) => 
                           z1_0_port, B(15) => m2_15_port, B(14) => m2_14_port,
                           B(13) => m2_13_port, B(12) => m2_12_port, B(11) => 
                           m2_11_port, B(10) => m2_10_port, B(9) => m2_9_port, 
                           B(8) => m2_8_port, B(7) => m2_7_port, B(6) => 
                           m2_6_port, B(5) => m2_5_port, B(4) => m2_4_port, 
                           B(3) => m2_3_port, B(2) => m2_2_port, B(1) => 
                           m2_1_port, B(0) => m2_0_port, CI => n61, SUM(15) => 
                           z2_temp_15_port, SUM(14) => z2_temp_14_port, SUM(13)
                           => z2_temp_13_port, SUM(12) => z2_temp_12_port, 
                           SUM(11) => z2_temp_11_port, SUM(10) => 
                           z2_temp_10_port, SUM(9) => z2_temp_9_port, SUM(8) =>
                           z2_temp_8_port, SUM(7) => z2_temp_7_port, SUM(6) => 
                           z2_temp_6_port, SUM(5) => z2_temp_5_port, SUM(4) => 
                           z2_temp_4_port, SUM(3) => z2_temp_3_port, SUM(2) => 
                           z2_temp_2_port, SUM(1) => z2_temp_1_port, SUM(0) => 
                           z2_temp_0_port, CO => n_1123);
   mult_28_C92 : siso_gen_DW_mult_tc_10 port map( a(15) => coeff_memory_79_port
                           , a(14) => coeff_memory_78_port, a(13) => 
                           coeff_memory_77_port, a(12) => coeff_memory_76_port,
                           a(11) => coeff_memory_75_port, a(10) => 
                           coeff_memory_74_port, a(9) => coeff_memory_73_port, 
                           a(8) => coeff_memory_72_port, a(7) => 
                           coeff_memory_71_port, a(6) => coeff_memory_70_port, 
                           a(5) => coeff_memory_69_port, a(4) => 
                           coeff_memory_68_port, a(3) => coeff_memory_67_port, 
                           a(2) => coeff_memory_66_port, a(1) => 
                           coeff_memory_65_port, a(0) => coeff_memory_64_port, 
                           b(15) => data_in(15), b(14) => data_in(14), b(13) =>
                           data_in(13), b(12) => data_in(12), b(11) => 
                           data_in(11), b(10) => data_in(10), b(9) => 
                           data_in(9), b(8) => data_in(8), b(7) => data_in(7), 
                           b(6) => data_in(6), b(5) => data_in(5), b(4) => 
                           data_in(4), b(3) => data_in(3), b(2) => data_in(2), 
                           b(1) => data_in(1), b(0) => data_in(0), product(31) 
                           => n_1124, product(30) => n_1125, product(29) => 
                           m1_15_port, product(28) => m1_14_port, product(27) 
                           => m1_13_port, product(26) => m1_12_port, 
                           product(25) => m1_11_port, product(24) => m1_10_port
                           , product(23) => m1_9_port, product(22) => m1_8_port
                           , product(21) => m1_7_port, product(20) => m1_6_port
                           , product(19) => m1_5_port, product(18) => m1_4_port
                           , product(17) => m1_3_port, product(16) => m1_2_port
                           , product(15) => m1_1_port, product(14) => m1_0_port
                           , product(13) => n_1126, product(12) => n_1127, 
                           product(11) => n_1128, product(10) => n_1129, 
                           product(9) => n_1130, product(8) => n_1131, 
                           product(7) => n_1132, product(6) => n_1133, 
                           product(5) => n_1134, product(4) => n_1135, 
                           product(3) => n_1136, product(2) => n_1137, 
                           product(1) => n_1138, product(0) => n_1139);
   add_102 : siso_gen_DW01_add_13 port map( A(15) => z2_15_port, A(14) => 
                           z2_14_port, A(13) => z2_13_port, A(12) => z2_12_port
                           , A(11) => z2_11_port, A(10) => z2_10_port, A(9) => 
                           z2_9_port, A(8) => z2_8_port, A(7) => z2_7_port, 
                           A(6) => z2_6_port, A(5) => z2_5_port, A(4) => 
                           z2_4_port, A(3) => z2_3_port, A(2) => z2_2_port, 
                           A(1) => z2_1_port, A(0) => z2_0_port, B(15) => 
                           m1_15_port, B(14) => m1_14_port, B(13) => m1_13_port
                           , B(12) => m1_12_port, B(11) => m1_11_port, B(10) =>
                           m1_10_port, B(9) => m1_9_port, B(8) => m1_8_port, 
                           B(7) => m1_7_port, B(6) => m1_6_port, B(5) => 
                           m1_5_port, B(4) => m1_4_port, B(3) => m1_3_port, 
                           B(2) => m1_2_port, B(1) => m1_1_port, B(0) => 
                           m1_0_port, CI => n61, SUM(15) => y_15_port, SUM(14) 
                           => y_14_port, SUM(13) => y_13_port, SUM(12) => 
                           y_12_port, SUM(11) => y_11_port, SUM(10) => 
                           y_10_port, SUM(9) => y_9_port, SUM(8) => y_8_port, 
                           SUM(7) => y_7_port, SUM(6) => y_6_port, SUM(5) => 
                           y_5_port, SUM(4) => y_4_port, SUM(3) => y_3_port, 
                           SUM(2) => y_2_port, SUM(1) => y_1_port, SUM(0) => 
                           y_0_port, CO => n_1140);
   add_0_root_add_0_root_add_101 : siso_gen_DW01_add_11 port map( A(15) => 
                           z2_temp_15_port, A(14) => z2_temp_14_port, A(13) => 
                           z2_temp_13_port, A(12) => z2_temp_12_port, A(11) => 
                           z2_temp_11_port, A(10) => z2_temp_10_port, A(9) => 
                           z2_temp_9_port, A(8) => z2_temp_8_port, A(7) => 
                           z2_temp_7_port, A(6) => z2_temp_6_port, A(5) => 
                           z2_temp_5_port, A(4) => z2_temp_4_port, A(3) => 
                           z2_temp_3_port, A(2) => z2_temp_2_port, A(1) => 
                           z2_temp_1_port, A(0) => z2_temp_0_port, B(15) => 
                           m3_15_port, B(14) => m3_14_port, B(13) => m3_13_port
                           , B(12) => m3_12_port, B(11) => m3_11_port, B(10) =>
                           m3_10_port, B(9) => m3_9_port, B(8) => m3_8_port, 
                           B(7) => m3_7_port, B(6) => m3_6_port, B(5) => 
                           m3_5_port, B(4) => m3_4_port, B(3) => m3_3_port, 
                           B(2) => m3_2_port, B(1) => m3_1_port, B(0) => 
                           m3_0_port, CI => n61, SUM(15) => z2_next_15_port, 
                           SUM(14) => z2_next_14_port, SUM(13) => 
                           z2_next_13_port, SUM(12) => z2_next_12_port, SUM(11)
                           => z2_next_11_port, SUM(10) => z2_next_10_port, 
                           SUM(9) => z2_next_9_port, SUM(8) => z2_next_8_port, 
                           SUM(7) => z2_next_7_port, SUM(6) => z2_next_6_port, 
                           SUM(5) => z2_next_5_port, SUM(4) => z2_next_4_port, 
                           SUM(3) => z2_next_3_port, SUM(2) => z2_next_2_port, 
                           SUM(1) => z2_next_1_port, SUM(0) => z2_next_0_port, 
                           CO => n_1141);
   add_99 : siso_gen_DW01_add_12 port map( A(15) => m4_15_port, A(14) => 
                           m4_14_port, A(13) => m4_13_port, A(12) => m4_12_port
                           , A(11) => m4_11_port, A(10) => m4_10_port, A(9) => 
                           m4_9_port, A(8) => m4_8_port, A(7) => m4_7_port, 
                           A(6) => m4_6_port, A(5) => m4_5_port, A(4) => 
                           m4_4_port, A(3) => m4_3_port, A(2) => m4_2_port, 
                           A(1) => m4_1_port, A(0) => m4_0_port, B(15) => 
                           m5_15_port, B(14) => m5_14_port, B(13) => m5_13_port
                           , B(12) => m5_12_port, B(11) => m5_11_port, B(10) =>
                           m5_10_port, B(9) => m5_9_port, B(8) => m5_8_port, 
                           B(7) => m5_7_port, B(6) => m5_6_port, B(5) => 
                           m5_5_port, B(4) => m5_4_port, B(3) => m5_3_port, 
                           B(2) => m5_2_port, B(1) => m5_1_port, B(0) => 
                           m5_0_port, CI => n61, SUM(15) => z1_next_15_port, 
                           SUM(14) => z1_next_14_port, SUM(13) => 
                           z1_next_13_port, SUM(12) => z1_next_12_port, SUM(11)
                           => z1_next_11_port, SUM(10) => z1_next_10_port, 
                           SUM(9) => z1_next_9_port, SUM(8) => z1_next_8_port, 
                           SUM(7) => z1_next_7_port, SUM(6) => z1_next_6_port, 
                           SUM(5) => z1_next_5_port, SUM(4) => z1_next_4_port, 
                           SUM(3) => z1_next_3_port, SUM(2) => z1_next_2_port, 
                           SUM(1) => z1_next_1_port, SUM(0) => z1_next_0_port, 
                           CO => n_1142);
   mult_28_C95 : siso_gen_DW_mult_tc_17 port map( a(15) => coeff_memory_31_port
                           , a(14) => coeff_memory_30_port, a(13) => 
                           coeff_memory_29_port, a(12) => coeff_memory_28_port,
                           a(11) => coeff_memory_27_port, a(10) => 
                           coeff_memory_26_port, a(9) => coeff_memory_25_port, 
                           a(8) => coeff_memory_24_port, a(7) => 
                           coeff_memory_23_port, a(6) => coeff_memory_22_port, 
                           a(5) => coeff_memory_21_port, a(4) => 
                           coeff_memory_20_port, a(3) => coeff_memory_19_port, 
                           a(2) => coeff_memory_18_port, a(1) => 
                           coeff_memory_17_port, a(0) => coeff_memory_16_port, 
                           b(15) => y_15_port, b(14) => y_14_port, b(13) => 
                           y_13_port, b(12) => y_12_port, b(11) => y_11_port, 
                           b(10) => n42, b(9) => y_9_port, b(8) => y_8_port, 
                           b(7) => y_7_port, b(6) => y_6_port, b(5) => n38, 
                           b(4) => y_4_port, b(3) => y_3_port, b(2) => y_2_port
                           , b(1) => n36, b(0) => n39, product(31) => n_1143, 
                           product(30) => n_1144, product(29) => m3_15_port, 
                           product(28) => m3_14_port, product(27) => m3_13_port
                           , product(26) => m3_12_port, product(25) => 
                           m3_11_port, product(24) => m3_10_port, product(23) 
                           => m3_9_port, product(22) => m3_8_port, product(21) 
                           => m3_7_port, product(20) => m3_6_port, product(19) 
                           => m3_5_port, product(18) => m3_4_port, product(17) 
                           => m3_3_port, product(16) => m3_2_port, product(15) 
                           => m3_1_port, product(14) => m3_0_port, product(13) 
                           => n_1145, product(12) => n_1146, product(11) => 
                           n_1147, product(10) => n_1148, product(9) => n_1149,
                           product(8) => n_1150, product(7) => n_1151, 
                           product(6) => n_1152, product(5) => n_1153, 
                           product(4) => n_1154, product(3) => n_1155, 
                           product(2) => n_1156, product(1) => n_1157, 
                           product(0) => n_1158);
   mult_28_C96 : siso_gen_DW_mult_tc_18 port map( a(15) => coeff_memory_15_port
                           , a(14) => coeff_memory_14_port, a(13) => 
                           coeff_memory_13_port, a(12) => coeff_memory_12_port,
                           a(11) => coeff_memory_11_port, a(10) => 
                           coeff_memory_10_port, a(9) => coeff_memory_9_port, 
                           a(8) => coeff_memory_8_port, a(7) => 
                           coeff_memory_7_port, a(6) => coeff_memory_6_port, 
                           a(5) => coeff_memory_5_port, a(4) => 
                           coeff_memory_4_port, a(3) => coeff_memory_3_port, 
                           a(2) => coeff_memory_2_port, a(1) => 
                           coeff_memory_1_port, a(0) => coeff_memory_0_port, 
                           b(15) => y_15_port, b(14) => y_14_port, b(13) => 
                           y_13_port, b(12) => y_12_port, b(11) => y_11_port, 
                           b(10) => n42, b(9) => y_9_port, b(8) => y_8_port, 
                           b(7) => y_7_port, b(6) => y_6_port, b(5) => n33, 
                           b(4) => y_4_port, b(3) => y_3_port, b(2) => n43, 
                           b(1) => n34, b(0) => n39, product(31) => n_1159, 
                           product(30) => n_1160, product(29) => m5_15_port, 
                           product(28) => m5_14_port, product(27) => m5_13_port
                           , product(26) => m5_12_port, product(25) => 
                           m5_11_port, product(24) => m5_10_port, product(23) 
                           => m5_9_port, product(22) => m5_8_port, product(21) 
                           => m5_7_port, product(20) => m5_6_port, product(19) 
                           => m5_5_port, product(18) => m5_4_port, product(17) 
                           => m5_3_port, product(16) => m5_2_port, product(15) 
                           => m5_1_port, product(14) => m5_0_port, product(13) 
                           => n_1161, product(12) => n_1162, product(11) => 
                           n_1163, product(10) => n_1164, product(9) => n_1165,
                           product(8) => n_1166, product(7) => n_1167, 
                           product(6) => n_1168, product(5) => n_1169, 
                           product(4) => n_1170, product(3) => n_1171, 
                           product(2) => n_1172, product(1) => n_1173, 
                           product(0) => n_1174);
   coeff_memory_reg_2_1_inst : DFERPQ1 port map( D => data_in(1), CEB => n27, 
                           CK => clk, RB => n52, Q => coeff_memory_33_port);
   coeff_memory_reg_4_1_inst : DFERPQ1 port map( D => data_in(1), CEB => n26, 
                           CK => clk, RB => n51, Q => coeff_memory_1_port);
   coeff_memory_reg_3_1_inst : DFERPQ1 port map( D => data_in(1), CEB => n28, 
                           CK => clk, RB => n60, Q => coeff_memory_17_port);
   data_out_reg_15_inst : DFERPQL port map( D => y_15_port, CEB => n23, CK => 
                           clk, RB => n45, Q => data_out(15));
   z2_reg_5_inst : DFERPQ1 port map( D => z2_next_5_port, CEB => n23, CK => clk
                           , RB => n47, Q => z2_5_port);
   coeff_counter_reg_0_inst : DFFRPQ1 port map( D => n32, CK => clk, RB => n53,
                           Q => coeff_counter_0_port);
   coeff_counter_reg_2_inst : DFFRPQ1 port map( D => n30, CK => clk, RB => n60,
                           Q => coeff_counter_2_port);
   coeff_counter_reg_1_inst : DFFRPQ1 port map( D => n31, CK => clk, RB => n60,
                           Q => coeff_counter_1_port);
   z1_reg_5_inst : DFERPQ1 port map( D => z1_next_5_port, CEB => n23, CK => clk
                           , RB => n50, Q => z1_5_port);
   z1_reg_4_inst : DFERPQ1 port map( D => z1_next_4_port, CEB => n23, CK => clk
                           , RB => n50, Q => z1_4_port);
   z1_reg_2_inst : DFERPQ1 port map( D => z1_next_2_port, CEB => n23, CK => clk
                           , RB => n50, Q => z1_2_port);
   z1_reg_3_inst : DFERPQ1 port map( D => z1_next_3_port, CEB => n23, CK => clk
                           , RB => n50, Q => z1_3_port);
   z1_reg_1_inst : DFERPQ1 port map( D => z1_next_1_port, CEB => n23, CK => clk
                           , RB => n50, Q => z1_1_port);
   z1_reg_0_inst : DFERPQ1 port map( D => z1_next_0_port, CEB => n23, CK => clk
                           , RB => n50, Q => z1_0_port);
   ready_reg : DFFRPQ1 port map( D => n22, CK => clk, RB => n53, Q => 
                           ready_port);
   coeff_memory_reg_4_0_inst : DFERPQ1 port map( D => data_in(0), CEB => n26, 
                           CK => clk, RB => n51, Q => coeff_memory_0_port);
   coeff_memory_reg_3_0_inst : DFERPQ1 port map( D => data_in(0), CEB => n28, 
                           CK => clk, RB => n60, Q => coeff_memory_16_port);
   coeff_memory_reg_4_2_inst : DFERPQ1 port map( D => data_in(2), CEB => n26, 
                           CK => clk, RB => n51, Q => coeff_memory_2_port);
   coeff_memory_reg_3_2_inst : DFERPQ1 port map( D => data_in(2), CEB => n28, 
                           CK => clk, RB => n60, Q => coeff_memory_18_port);
   coeff_memory_reg_4_4_inst : DFERPQ1 port map( D => data_in(4), CEB => n26, 
                           CK => clk, RB => n51, Q => coeff_memory_4_port);
   coeff_memory_reg_3_4_inst : DFERPQ1 port map( D => data_in(4), CEB => n28, 
                           CK => clk, RB => n48, Q => coeff_memory_20_port);
   coeff_memory_reg_4_6_inst : DFERPQ1 port map( D => data_in(6), CEB => n26, 
                           CK => clk, RB => n51, Q => coeff_memory_6_port);
   coeff_memory_reg_3_6_inst : DFERPQ1 port map( D => data_in(6), CEB => n28, 
                           CK => clk, RB => n48, Q => coeff_memory_22_port);
   coeff_memory_reg_4_8_inst : DFERPQ1 port map( D => data_in(8), CEB => n26, 
                           CK => clk, RB => n52, Q => coeff_memory_8_port);
   coeff_memory_reg_4_3_inst : DFERPQ1 port map( D => data_in(3), CEB => n26, 
                           CK => clk, RB => n51, Q => coeff_memory_3_port);
   z2_reg_4_inst : DFERPQ1 port map( D => z2_next_4_port, CEB => n23, CK => clk
                           , RB => n47, Q => z2_4_port);
   coeff_memory_reg_3_8_inst : DFERPQ1 port map( D => data_in(8), CEB => n28, 
                           CK => clk, RB => n48, Q => coeff_memory_24_port);
   coeff_memory_reg_3_3_inst : DFERPQ1 port map( D => data_in(3), CEB => n28, 
                           CK => clk, RB => n60, Q => coeff_memory_19_port);
   coeff_memory_reg_4_10_inst : DFERPQ1 port map( D => data_in(10), CEB => n26,
                           CK => clk, RB => n52, Q => coeff_memory_10_port);
   coeff_memory_reg_3_10_inst : DFERPQ1 port map( D => data_in(10), CEB => n28,
                           CK => clk, RB => n48, Q => coeff_memory_26_port);
   coeff_memory_reg_4_15_inst : DFERPQ1 port map( D => data_in(15), CEB => n26,
                           CK => clk, RB => n52, Q => coeff_memory_15_port);
   z2_reg_3_inst : DFERPQ1 port map( D => z2_next_3_port, CEB => n23, CK => clk
                           , RB => n47, Q => z2_3_port);
   coeff_memory_reg_4_5_inst : DFERPQ1 port map( D => data_in(5), CEB => n26, 
                           CK => clk, RB => n51, Q => coeff_memory_5_port);
   coeff_memory_reg_4_12_inst : DFERPQ1 port map( D => data_in(12), CEB => n26,
                           CK => clk, RB => n52, Q => coeff_memory_12_port);
   coeff_memory_reg_3_15_inst : DFERPQ1 port map( D => data_in(15), CEB => n28,
                           CK => clk, RB => n48, Q => coeff_memory_31_port);
   z2_reg_2_inst : DFERPQ1 port map( D => z2_next_2_port, CEB => n23, CK => clk
                           , RB => n47, Q => z2_2_port);
   coeff_memory_reg_3_12_inst : DFERPQ1 port map( D => data_in(12), CEB => n28,
                           CK => clk, RB => n48, Q => coeff_memory_28_port);
   coeff_memory_reg_3_5_inst : DFERPQ1 port map( D => data_in(5), CEB => n28, 
                           CK => clk, RB => n48, Q => coeff_memory_21_port);
   coeff_memory_reg_4_14_inst : DFERPQ1 port map( D => data_in(14), CEB => n26,
                           CK => clk, RB => n52, Q => coeff_memory_14_port);
   coeff_memory_reg_3_14_inst : DFERPQ1 port map( D => data_in(14), CEB => n28,
                           CK => clk, RB => n48, Q => coeff_memory_30_port);
   coeff_memory_reg_3_7_inst : DFERPQ1 port map( D => data_in(7), CEB => n28, 
                           CK => clk, RB => n48, Q => coeff_memory_23_port);
   z2_reg_1_inst : DFERPQ1 port map( D => z2_next_1_port, CEB => n23, CK => clk
                           , RB => n47, Q => z2_1_port);
   coeff_memory_reg_4_9_inst : DFERPQ1 port map( D => data_in(9), CEB => n26, 
                           CK => clk, RB => n52, Q => coeff_memory_9_port);
   coeff_memory_reg_3_9_inst : DFERPQ1 port map( D => data_in(9), CEB => n28, 
                           CK => clk, RB => n48, Q => coeff_memory_25_port);
   z2_reg_0_inst : DFERPQ1 port map( D => z2_next_0_port, CEB => n23, CK => clk
                           , RB => n47, Q => z2_0_port);
   coeff_memory_reg_4_11_inst : DFERPQ1 port map( D => data_in(11), CEB => n26,
                           CK => clk, RB => n52, Q => coeff_memory_11_port);
   coeff_memory_reg_2_15_inst : DFERPQ1 port map( D => data_in(15), CEB => n27,
                           CK => clk, RB => n53, Q => coeff_memory_47_port);
   coeff_memory_reg_3_11_inst : DFERPQ1 port map( D => data_in(11), CEB => n28,
                           CK => clk, RB => n48, Q => coeff_memory_27_port);
   coeff_memory_reg_4_13_inst : DFERPQ1 port map( D => data_in(13), CEB => n26,
                           CK => clk, RB => n52, Q => coeff_memory_13_port);
   coeff_memory_reg_3_13_inst : DFERPQ1 port map( D => data_in(13), CEB => n28,
                           CK => clk, RB => n48, Q => coeff_memory_29_port);
   coeff_memory_reg_2_0_inst : DFERPQ1 port map( D => data_in(0), CEB => n27, 
                           CK => clk, RB => n52, Q => coeff_memory_32_port);
   coeff_memory_reg_2_14_inst : DFERPQ1 port map( D => data_in(14), CEB => n27,
                           CK => clk, RB => n53, Q => coeff_memory_46_port);
   coeff_memory_reg_2_12_inst : DFERPQ1 port map( D => data_in(12), CEB => n27,
                           CK => clk, RB => n53, Q => coeff_memory_44_port);
   coeff_memory_reg_2_4_inst : DFERPQ1 port map( D => data_in(4), CEB => n27, 
                           CK => clk, RB => n52, Q => coeff_memory_36_port);
   coeff_memory_reg_2_13_inst : DFERPQ1 port map( D => data_in(13), CEB => n27,
                           CK => clk, RB => n53, Q => coeff_memory_45_port);
   coeff_memory_reg_2_11_inst : DFERPQ1 port map( D => data_in(11), CEB => n27,
                           CK => clk, RB => n53, Q => coeff_memory_43_port);
   coeff_memory_reg_2_8_inst : DFERPQ1 port map( D => data_in(8), CEB => n27, 
                           CK => clk, RB => n53, Q => coeff_memory_40_port);
   coeff_memory_reg_2_2_inst : DFERPQ1 port map( D => data_in(2), CEB => n27, 
                           CK => clk, RB => n52, Q => coeff_memory_34_port);
   coeff_memory_reg_2_10_inst : DFERPQ1 port map( D => data_in(10), CEB => n27,
                           CK => clk, RB => n53, Q => coeff_memory_42_port);
   coeff_memory_reg_2_6_inst : DFERPQ1 port map( D => data_in(6), CEB => n27, 
                           CK => clk, RB => n53, Q => coeff_memory_38_port);
   coeff_memory_reg_2_7_inst : DFERPQ1 port map( D => data_in(7), CEB => n27, 
                           CK => clk, RB => n53, Q => coeff_memory_39_port);
   coeff_memory_reg_2_3_inst : DFERPQ1 port map( D => data_in(3), CEB => n27, 
                           CK => clk, RB => n52, Q => coeff_memory_35_port);
   coeff_memory_reg_2_9_inst : DFERPQ1 port map( D => data_in(9), CEB => n27, 
                           CK => clk, RB => n53, Q => coeff_memory_41_port);
   coeff_memory_reg_2_5_inst : DFERPQ1 port map( D => data_in(5), CEB => n27, 
                           CK => clk, RB => n53, Q => coeff_memory_37_port);
   coeff_memory_reg_1_15_inst : DFERPQ1 port map( D => data_in(15), CEB => n29,
                           CK => clk, RB => n50, Q => coeff_memory_63_port);
   coeff_memory_reg_1_0_inst : DFERPQ1 port map( D => data_in(0), CEB => n29, 
                           CK => clk, RB => n48, Q => coeff_memory_48_port);
   coeff_memory_reg_1_14_inst : DFERPQ1 port map( D => data_in(14), CEB => n29,
                           CK => clk, RB => n50, Q => coeff_memory_62_port);
   coeff_memory_reg_1_12_inst : DFERPQ1 port map( D => data_in(12), CEB => n29,
                           CK => clk, RB => n49, Q => coeff_memory_60_port);
   coeff_memory_reg_1_4_inst : DFERPQ1 port map( D => data_in(4), CEB => n29, 
                           CK => clk, RB => n49, Q => coeff_memory_52_port);
   coeff_memory_reg_1_13_inst : DFERPQ1 port map( D => data_in(13), CEB => n29,
                           CK => clk, RB => n49, Q => coeff_memory_61_port);
   coeff_memory_reg_1_11_inst : DFERPQ1 port map( D => data_in(11), CEB => n29,
                           CK => clk, RB => n49, Q => coeff_memory_59_port);
   coeff_memory_reg_1_8_inst : DFERPQ1 port map( D => data_in(8), CEB => n29, 
                           CK => clk, RB => n49, Q => coeff_memory_56_port);
   coeff_memory_reg_1_2_inst : DFERPQ1 port map( D => data_in(2), CEB => n29, 
                           CK => clk, RB => n49, Q => coeff_memory_50_port);
   coeff_memory_reg_1_10_inst : DFERPQ1 port map( D => data_in(10), CEB => n29,
                           CK => clk, RB => n49, Q => coeff_memory_58_port);
   coeff_memory_reg_1_6_inst : DFERPQ1 port map( D => data_in(6), CEB => n29, 
                           CK => clk, RB => n49, Q => coeff_memory_54_port);
   coeff_memory_reg_1_7_inst : DFERPQ1 port map( D => data_in(7), CEB => n29, 
                           CK => clk, RB => n49, Q => coeff_memory_55_port);
   coeff_memory_reg_1_1_inst : DFERPQ1 port map( D => data_in(1), CEB => n29, 
                           CK => clk, RB => n49, Q => coeff_memory_49_port);
   coeff_memory_reg_1_3_inst : DFERPQ1 port map( D => data_in(3), CEB => n29, 
                           CK => clk, RB => n49, Q => coeff_memory_51_port);
   coeff_memory_reg_1_9_inst : DFERPQ1 port map( D => data_in(9), CEB => n29, 
                           CK => clk, RB => n49, Q => coeff_memory_57_port);
   coeff_memory_reg_1_5_inst : DFERPQ1 port map( D => data_in(5), CEB => n29, 
                           CK => clk, RB => n49, Q => coeff_memory_53_port);
   coeff_memory_reg_0_0_inst : DFERPQ1 port map( D => data_in(0), CEB => n25, 
                           CK => clk, RB => n46, Q => coeff_memory_64_port);
   coeff_memory_reg_0_14_inst : DFERPQ1 port map( D => data_in(14), CEB => n25,
                           CK => clk, RB => n47, Q => coeff_memory_78_port);
   coeff_memory_reg_0_10_inst : DFERPQ1 port map( D => data_in(10), CEB => n25,
                           CK => clk, RB => n47, Q => coeff_memory_74_port);
   coeff_memory_reg_0_8_inst : DFERPQ1 port map( D => data_in(8), CEB => n25, 
                           CK => clk, RB => n46, Q => coeff_memory_72_port);
   coeff_memory_reg_0_6_inst : DFERPQ1 port map( D => data_in(6), CEB => n25, 
                           CK => clk, RB => n46, Q => coeff_memory_70_port);
   coeff_memory_reg_0_4_inst : DFERPQ1 port map( D => data_in(4), CEB => n25, 
                           CK => clk, RB => n46, Q => coeff_memory_68_port);
   coeff_memory_reg_0_2_inst : DFERPQ1 port map( D => data_in(2), CEB => n25, 
                           CK => clk, RB => n46, Q => coeff_memory_66_port);
   coeff_memory_reg_0_12_inst : DFERPQ1 port map( D => data_in(12), CEB => n25,
                           CK => clk, RB => n47, Q => coeff_memory_76_port);
   data_out_reg_14_inst : DFERPQL port map( D => y_14_port, CEB => n23, CK => 
                           clk, RB => n45, Q => data_out(14));
   data_out_reg_13_inst : DFERPQL port map( D => y_13_port, CEB => n23, CK => 
                           clk, RB => n45, Q => data_out(13));
   data_out_reg_12_inst : DFERPQL port map( D => y_12_port, CEB => n23, CK => 
                           clk, RB => n45, Q => data_out(12));
   data_out_reg_11_inst : DFERPQL port map( D => y_11_port, CEB => n23, CK => 
                           clk, RB => n45, Q => data_out(11));
   data_out_reg_10_inst : DFERPQL port map( D => n42, CEB => n23, CK => clk, RB
                           => n45, Q => data_out(10));
   data_out_reg_9_inst : DFERPQL port map( D => y_9_port, CEB => n23, CK => clk
                           , RB => n45, Q => data_out(9));
   data_out_reg_8_inst : DFERPQL port map( D => y_8_port, CEB => n23, CK => clk
                           , RB => n45, Q => data_out(8));
   data_out_reg_7_inst : DFERPQL port map( D => y_7_port, CEB => n23, CK => clk
                           , RB => n45, Q => data_out(7));
   data_out_reg_6_inst : DFERPQL port map( D => y_6_port, CEB => n23, CK => clk
                           , RB => n45, Q => data_out(6));
   data_out_reg_5_inst : DFERPQL port map( D => n38, CEB => n23, CK => clk, RB 
                           => n45, Q => data_out(5));
   data_out_reg_3_inst : DFERPQL port map( D => y_3_port, CEB => n23, CK => clk
                           , RB => n45, Q => data_out(3));
   data_out_reg_1_inst : DFERPQL port map( D => n36, CEB => n23, CK => clk, RB 
                           => n46, Q => data_out(1));
   data_out_reg_0_inst : DFERPQ1 port map( D => n39, CEB => n23, CK => clk, RB 
                           => n46, Q => data_out(0));
   data_out_reg_4_inst : DFERPQ1 port map( D => n44, CEB => n23, CK => clk, RB 
                           => n45, Q => data_out(4));
   data_out_reg_2_inst : DFERPQL port map( D => n43, CEB => n23, CK => clk, RB 
                           => n46, Q => data_out(2));
   z1_reg_15_inst : DFERPQ1 port map( D => z1_next_15_port, CEB => n23, CK => 
                           clk, RB => n60, Q => z1_15_port);
   z1_reg_14_inst : DFERPQ1 port map( D => z1_next_14_port, CEB => n23, CK => 
                           clk, RB => n60, Q => z1_14_port);
   z1_reg_13_inst : DFERPQ1 port map( D => z1_next_13_port, CEB => n23, CK => 
                           clk, RB => n60, Q => z1_13_port);
   z1_reg_12_inst : DFERPQ1 port map( D => z1_next_12_port, CEB => n23, CK => 
                           clk, RB => n60, Q => z1_12_port);
   z1_reg_8_inst : DFERPQ1 port map( D => z1_next_8_port, CEB => n23, CK => clk
                           , RB => n60, Q => z1_8_port);
   z1_reg_11_inst : DFERPQ1 port map( D => z1_next_11_port, CEB => n23, CK => 
                           clk, RB => n60, Q => z1_11_port);
   z1_reg_10_inst : DFERPQ1 port map( D => z1_next_10_port, CEB => n23, CK => 
                           clk, RB => n60, Q => z1_10_port);
   z1_reg_9_inst : DFERPQ1 port map( D => z1_next_9_port, CEB => n23, CK => clk
                           , RB => n60, Q => z1_9_port);
   z1_reg_7_inst : DFERPQ1 port map( D => z1_next_7_port, CEB => n23, CK => clk
                           , RB => n60, Q => z1_7_port);
   z1_reg_6_inst : DFERPQ1 port map( D => z1_next_6_port, CEB => n23, CK => clk
                           , RB => n60, Q => z1_6_port);
   z2_reg_15_inst : DFERPQ1 port map( D => z2_next_15_port, CEB => n23, CK => 
                           clk, RB => n60, Q => z2_15_port);
   z2_reg_14_inst : DFERPQ1 port map( D => z2_next_14_port, CEB => n23, CK => 
                           clk, RB => n60, Q => z2_14_port);
   z2_reg_10_inst : DFERPQ1 port map( D => z2_next_10_port, CEB => n23, CK => 
                           clk, RB => n60, Q => z2_10_port);
   z2_reg_12_inst : DFERPQ1 port map( D => z2_next_12_port, CEB => n23, CK => 
                           clk, RB => n60, Q => z2_12_port);
   z2_reg_11_inst : DFERPQ1 port map( D => z2_next_11_port, CEB => n23, CK => 
                           clk, RB => n60, Q => z2_11_port);
   z2_reg_13_inst : DFERPQ1 port map( D => z2_next_13_port, CEB => n23, CK => 
                           clk, RB => n60, Q => z2_13_port);
   z2_reg_8_inst : DFERPQ1 port map( D => z2_next_8_port, CEB => n23, CK => clk
                           , RB => n60, Q => z2_8_port);
   z2_reg_7_inst : DFERPQ1 port map( D => z2_next_7_port, CEB => n23, CK => clk
                           , RB => n60, Q => z2_7_port);
   z2_reg_9_inst : DFERPQ1 port map( D => z2_next_9_port, CEB => n23, CK => clk
                           , RB => n60, Q => z2_9_port);
   z2_reg_6_inst : DFERPQ1 port map( D => z2_next_6_port, CEB => n23, CK => clk
                           , RB => n60, Q => z2_6_port);
   coeff_memory_reg_0_1_inst : DFERPQ4 port map( D => data_in(1), CEB => n25, 
                           CK => clk, RB => n46, Q => coeff_memory_65_port);
   coeff_memory_reg_0_11_inst : DFERPQ2 port map( D => data_in(11), CEB => n25,
                           CK => clk, RB => n47, Q => coeff_memory_75_port);
   coeff_memory_reg_0_5_inst : DFERPQ4 port map( D => data_in(5), CEB => n25, 
                           CK => clk, RB => n46, Q => coeff_memory_69_port);
   coeff_memory_reg_0_7_inst : DFERPQ4 port map( D => data_in(7), CEB => n25, 
                           CK => clk, RB => n46, Q => coeff_memory_71_port);
   coeff_memory_reg_0_3_inst : DFERPQ4 port map( D => data_in(3), CEB => n25, 
                           CK => clk, RB => n46, Q => coeff_memory_67_port);
   coeff_memory_reg_0_13_inst : DFERPQ2 port map( D => data_in(13), CEB => n25,
                           CK => clk, RB => n47, Q => coeff_memory_77_port);
   coeff_memory_reg_4_7_inst : DFERPQL port map( D => data_in(7), CEB => n26, 
                           CK => clk, RB => n60, Q => coeff_memory_7_port);
   coeff_memory_reg_0_9_inst : DFERPQ4 port map( D => data_in(9), CEB => n25, 
                           CK => clk, RB => n46, Q => coeff_memory_73_port);
   coeff_memory_reg_0_15_inst : DFERPQ1 port map( D => data_in(15), CEB => n25,
                           CK => clk, RB => n60, Q => coeff_memory_79_port);
   U21 : INVD4 port map( A => n35, Z => n36);
   U22 : INVD4 port map( A => n35, Z => n34);
   U23 : INVD4 port map( A => n37, Z => n33);
   U24 : INVBD4 port map( A => y_5_port, Z => n37);
   U25 : INVD4 port map( A => y_1_port, Z => n35);
   U26 : BUFD4 port map( A => y_10_port, Z => n42);
   U27 : INVD4 port map( A => n37, Z => n38);
   U28 : BUFD8 port map( A => y_0_port, Z => n39);
   U29 : INVD1 port map( A => n56, Z => n59);
   U30 : INVD1 port map( A => reset, Z => n46);
   U31 : INVD1 port map( A => reset, Z => n52);
   U32 : INVD1 port map( A => n54, Z => n48);
   U33 : INVD1 port map( A => reset, Z => n49);
   U34 : INVD1 port map( A => n54, Z => n53);
   U35 : INVD1 port map( A => n54, Z => n45);
   U36 : INVD1 port map( A => n54, Z => n47);
   U37 : INVD1 port map( A => n54, Z => n51);
   U38 : INVD1 port map( A => reset, Z => n50);
   U39 : NAN3D1 port map( A1 => n59, A2 => n58, A3 => n57, Z => n25);
   U40 : OA21D1 port map( A1 => n57, A2 => n58, B => n23, Z => n40);
   U41 : NAN2D1 port map( A1 => n41, A2 => n58, Z => n29);
   U42 : INVD1 port map( A => n60, Z => n54);
   U43 : INVD1 port map( A => coeff_counter_1_port, Z => n58);
   U44 : NAN2D1 port map( A1 => coeff_counter_2_port, A2 => n59, Z => n26);
   U45 : NAN2D1 port map( A1 => coeff_counter_1_port, A2 => n59, Z => n27);
   U46 : NAN2D1 port map( A1 => n41, A2 => coeff_counter_1_port, Z => n28);
   U47 : AND2D1 port map( A1 => n40, A2 => coeff_counter_0_port, Z => n41);
   U48 : INVD1 port map( A => coeff_counter_2_port, Z => n57);
   U49 : NAN2M1D1 port map( A1 => ready_port, A2 => n23, Z => n22);
   U50 : INVD1 port map( A => coeff_counter_0_port, Z => n55);
   U51 : INVD1 port map( A => reset, Z => n60);
   U52 : TIEHI port map( Z => req);
   U53 : TIELO port map( Z => n61);
   U54 : BUFD4 port map( A => y_2_port, Z => n43);
   U55 : BUFDL port map( A => y_4_port, Z => n44);
   U56 : NAN3D1 port map( A1 => coeff_counter_2_port, A2 => 
                           coeff_counter_0_port, A3 => n58, Z => n23);
   U57 : OAI21D1 port map( A1 => n41, A2 => n58, B => n29, Z => n31);
   U58 : NAN2D1 port map( A1 => n57, A2 => n28, Z => n30);
   U59 : NAN2D1 port map( A1 => n40, A2 => n55, Z => n56);
   U60 : OAI21D1 port map( A1 => n40, A2 => n55, B => n56, Z => n32);

end hier_sec_par_16_5;
