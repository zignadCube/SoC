
library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

package CONV_PACK_siso_gen is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_siso_gen;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_siso_gen.all;

architecture flat_dpctrl_gcd_16_10 of siso_gen is

   component AOI211D1
      port( A1, A2, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211D1
      port( A1, A2, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN3M1D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFRPQ1
      port( D, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFSPQ1
      port( D, CK, SB : in std_logic;  Q : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AO211D1
      port( A1, A2, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN4D1
      port( A1, A2, A3, A4 : in std_logic;  Z : out std_logic);
   end component;
   
   component TIELO
      port( Z : out std_logic);
   end component;
   
   component TIEHI
      port( Z : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component EXOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component DFERPQ1
      port( D, CEB, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component BUFD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4D1
      port( A1, A2, A3, A4 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI32D1
      port( A1, A2, A3, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AO32D1
      port( A1, A2, A3, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI32D1
      port( A1, A2, A3, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22M10D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3M1D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4M1D1
      port( A1, A2, A3, A4 : in std_logic;  Z : out std_logic);
   end component;
   
   signal data_out_15_port, data_out_14_port, data_out_13_port, 
      data_out_12_port, data_out_11_port, data_out_10_port, data_out_9_port, 
      data_out_8_port, data_out_7_port, data_out_6_port, data_out_5_port, 
      data_out_4_port, data_out_3_port, data_out_2_port, data_out_1_port, 
      data_out_0_port, add_l_sel, add_r_sel, add_l_en, add_r_en, sub, cmp_r_sel
      , cmp_l_en, cmp_r_en, rd_addr_1_port, rd_addr_0_port, wr_addr_0, 
      wr_sel_en_1_port, wr_sel_en_0_port, equal, greater, n1, dp_n_1001, 
      dp_n2020, dp_n2010, dp_n200, dp_n199, dp_n198, dp_n197, dp_n196, dp_n195,
      dp_n194, dp_n193, dp_n192, dp_n191, dp_n1901, dp_n189, dp_n188, dp_n187, 
      dp_n186, dp_n185, dp_n184, dp_n183, dp_n182, dp_n181, dp_n1801, dp_n179, 
      dp_n178, dp_n177, dp_n176, dp_n175, dp_n174, dp_n173, dp_n172, dp_n171, 
      dp_n170, dp_n169, dp_n168, dp_n1670, dp_n1660, dp_n1650, dp_n1640, 
      dp_n1630, dp_n1620, dp_n1610, dp_n1600, dp_n1590, dp_n1580, dp_n1570, 
      dp_n1560, dp_n1550, dp_n1540, dp_n1530, dp_n1520, dp_n151, dp_n1500, 
      dp_n1490, dp_n1480, dp_n1470, dp_n1460, dp_n1450, dp_n1440, dp_n1430, 
      dp_n1420, dp_n1410, dp_n1400, dp_n1390, dp_n1380, dp_n1370, dp_n1360, 
      dp_n1350, dp_n134, dp_n1330, dp_n1320, dp_n1310, dp_n1300, dp_n1290, 
      dp_n1280, dp_n1270, dp_n1260, dp_n1250, dp_n1240, dp_n1230, dp_n1220, 
      dp_n1210, dp_n1200, dp_n1190, dp_n58, dp_n57, dp_n56, dp_n55, dp_n54, 
      dp_n53, dp_n52, dp_n51, dp_n50, dp_n49, dp_n48, dp_n47, dp_n46, dp_n45, 
      dp_n44, dp_n43, dp_n42, dp_n41, dp_n40, dp_n39, dp_n38, dp_n37, dp_n36, 
      dp_n35, dp_n34, dp_n33, dp_n32, dp_n31, dp_n30, dp_n29, dp_n28, dp_n27, 
      dp_n26, dp_n25, dp_n24, dp_n23, dp_n22, dp_n21, dp_n20, dp_n1900, 
      dp_n1800, dp_n17, dp_n16, dp_n15, dp_n14, dp_n13, dp_n12, dp_n11, dp_n10,
      dp_n9, dp_n8, dp_n7, dp_n6, dp_n5, dp_n4, dp_n3, dp_n2, dp_n1, dp_n1180, 
      dp_n117, dp_n1160, dp_n1150, dp_n1140, dp_n1130, dp_n1120, dp_n1110, 
      dp_n1100, dp_n1090, dp_n1080, dp_n1070, dp_n1060, dp_n1050, dp_n1040, 
      dp_n1030, dp_n1020, dp_n1010, dp_n100, dp_n99, dp_n98, dp_n97, dp_n96, 
      dp_n95, dp_n94, dp_n93, dp_n92, dp_n91, dp_n90, dp_n89, dp_n88, dp_n87, 
      dp_n86, dp_n85, dp_n84, dp_n83, dp_n82, dp_n81, dp_n80, dp_n79, dp_n78, 
      dp_n77, dp_n76, dp_n75, dp_n74, dp_n73, dp_n72, dp_n71, dp_n70, dp_n69, 
      dp_n68, dp_n67, dp_n66, dp_n65, dp_n64, dp_n63, dp_n62, dp_n61, dp_n60, 
      dp_n59, dp_add_r_in_0, dp_add_r_in_1, dp_add_r_in_2, dp_add_r_in_3, 
      dp_add_r_in_4, dp_add_r_in_5, dp_add_r_in_6, dp_add_r_in_7, dp_add_r_in_8
      , dp_add_r_in_9, dp_add_r_in_10, dp_add_r_in_11, dp_add_r_in_12, 
      dp_add_r_in_13, dp_add_r_in_14, dp_add_r_in_15, dp_N167, dp_N166, dp_N165
      , dp_N164, dp_N163, dp_N162, dp_N161, dp_N160, dp_N159, dp_N158, dp_N157,
      dp_N156, dp_N155, dp_N154, dp_N153, dp_N152, dp_N150, dp_N149, dp_N148, 
      dp_N147, dp_N146, dp_N145, dp_N144, dp_N143, dp_N142, dp_N141, dp_N140, 
      dp_N139, dp_N138, dp_N137, dp_N136, dp_N135, dp_N133, dp_N132, dp_N131, 
      dp_N130, dp_N129, dp_N128, dp_N127, dp_N126, dp_N125, dp_N124, dp_N123, 
      dp_N122, dp_N121, dp_N120, dp_N119, dp_N118, dp_N116, dp_N115, dp_N114, 
      dp_N113, dp_N112, dp_N111, dp_N110, dp_N109, dp_N108, dp_N107, dp_N106, 
      dp_N105, dp_N104, dp_N103, dp_N102, dp_N101, dp_add_out_0_port, 
      dp_add_out_1_port, dp_add_out_2_port, dp_add_out_3_port, 
      dp_add_out_4_port, dp_add_out_5_port, dp_add_out_6_port, 
      dp_add_out_7_port, dp_add_out_8_port, dp_add_out_9_port, 
      dp_add_out_10_port, dp_add_out_11_port, dp_add_out_12_port, 
      dp_add_out_13_port, dp_add_out_14_port, dp_add_out_15_port, 
      dp_cmp_r_0_port, dp_cmp_r_1_port, dp_cmp_r_2_port, dp_cmp_r_3_port, 
      dp_cmp_r_4_port, dp_cmp_r_5_port, dp_cmp_r_6_port, dp_cmp_r_7_port, 
      dp_cmp_r_8_port, dp_cmp_r_9_port, dp_cmp_r_10_port, dp_cmp_r_11_port, 
      dp_cmp_r_12_port, dp_cmp_r_13_port, dp_cmp_r_14_port, dp_cmp_r_15_port, 
      dp_cmp_l_0_port, dp_cmp_l_1_port, dp_cmp_l_2_port, dp_cmp_l_3_port, 
      dp_cmp_l_4_port, dp_cmp_l_5_port, dp_cmp_l_6_port, dp_cmp_l_7_port, 
      dp_cmp_l_8_port, dp_cmp_l_9_port, dp_cmp_l_10_port, dp_cmp_l_11_port, 
      dp_cmp_l_12_port, dp_cmp_l_13_port, dp_cmp_l_14_port, dp_cmp_l_15_port, 
      dp_add_r_0_port, dp_add_r_1_port, dp_add_r_2_port, dp_add_r_3_port, 
      dp_add_r_4_port, dp_add_r_5_port, dp_add_r_6_port, dp_add_r_7_port, 
      dp_add_r_8_port, dp_add_r_9_port, dp_add_r_10_port, dp_add_r_11_port, 
      dp_add_r_12_port, dp_add_r_13_port, dp_add_r_14_port, dp_add_r_15_port, 
      dp_add_l_0_port, dp_add_l_1_port, dp_add_l_2_port, dp_add_l_3_port, 
      dp_add_l_4_port, dp_add_l_5_port, dp_add_l_6_port, dp_add_l_7_port, 
      dp_add_l_8_port, dp_add_l_9_port, dp_add_l_10_port, dp_add_l_11_port, 
      dp_add_l_12_port, dp_add_l_13_port, dp_add_l_14_port, dp_add_l_15_port, 
      dp_mem_0_port, dp_mem_1_port, dp_mem_2_port, dp_mem_3_port, dp_mem_4_port
      , dp_mem_5_port, dp_mem_6_port, dp_mem_7_port, dp_mem_8_port, 
      dp_mem_9_port, dp_mem_10_port, dp_mem_11_port, dp_mem_12_port, 
      dp_mem_13_port, dp_mem_14_port, dp_mem_15_port, dp_mem_16_port, 
      dp_mem_17_port, dp_mem_18_port, dp_mem_19_port, dp_mem_20_port, 
      dp_mem_21_port, dp_mem_22_port, dp_mem_23_port, dp_mem_24_port, 
      dp_mem_25_port, dp_mem_26_port, dp_mem_27_port, dp_mem_28_port, 
      dp_mem_29_port, dp_mem_30_port, dp_mem_31_port, dp_mem_32_port, 
      dp_mem_33_port, dp_mem_34_port, dp_mem_35_port, dp_mem_36_port, 
      dp_mem_37_port, dp_mem_38_port, dp_mem_39_port, dp_mem_40_port, 
      dp_mem_41_port, dp_mem_42_port, dp_mem_43_port, dp_mem_44_port, 
      dp_mem_45_port, dp_mem_46_port, dp_mem_47_port, dp_mem_48_port, 
      dp_mem_49_port, dp_mem_50_port, dp_mem_51_port, dp_mem_52_port, 
      dp_mem_53_port, dp_mem_54_port, dp_mem_55_port, dp_mem_56_port, 
      dp_mem_57_port, dp_mem_58_port, dp_mem_59_port, dp_mem_60_port, 
      dp_mem_61_port, dp_mem_62_port, dp_mem_63_port, 
      dp_add_1_root_add_129_2_carry_1_port, 
      dp_add_1_root_add_129_2_carry_2_port, 
      dp_add_1_root_add_129_2_carry_3_port, 
      dp_add_1_root_add_129_2_carry_4_port, 
      dp_add_1_root_add_129_2_carry_5_port, 
      dp_add_1_root_add_129_2_carry_6_port, 
      dp_add_1_root_add_129_2_carry_7_port, 
      dp_add_1_root_add_129_2_carry_8_port, 
      dp_add_1_root_add_129_2_carry_9_port, 
      dp_add_1_root_add_129_2_carry_10_port, 
      dp_add_1_root_add_129_2_carry_11_port, 
      dp_add_1_root_add_129_2_carry_12_port, 
      dp_add_1_root_add_129_2_carry_13_port, 
      dp_add_1_root_add_129_2_carry_14_port, 
      dp_add_1_root_add_129_2_carry_15_port, cn_n32, cn_n31, cn_n14, cn_n13, 
      cn_n12, cn_n11, cn_n9, cn_n8, cn_n7, cn_n6, cn_n3, cn_n2, cn_sub, 
      cn_wr_addr_1, cn_n30, cn_n29, cn_n28, cn_n27, cn_n26, cn_n25, cn_n24, 
      cn_n23, cn_n22, cn_n210, cn_n20, cn_n19, cn_n18, cn_n17, cn_n16, cn_n15, 
      cn_N21, cn_next_state_0_port, cn_next_state_1_port, cn_next_state_2_port,
      cn_current_state_0_port, cn_current_state_1_port, cn_current_state_2_port
      , cn_current_state_3_port, cn_cmp_l_sel : std_logic;

begin
   data_out <= ( data_out_15_port, data_out_14_port, data_out_13_port, 
      data_out_12_port, data_out_11_port, data_out_10_port, data_out_9_port, 
      data_out_8_port, data_out_7_port, data_out_6_port, data_out_5_port, 
      data_out_4_port, data_out_3_port, data_out_2_port, data_out_1_port, 
      data_out_0_port );
   
   U1 : TIELO port map( Z => n1);
   U2 : TIEHI port map( Z => sub);
   dp_U301 : OAI32D1 port map( A1 => dp_n1450, A2 => dp_n1440, A3 => dp_n1430, 
                           B1 => dp_n1420, B2 => dp_n1450, Z => greater);
   dp_U300 : NOR4M1D1 port map( A1 => dp_n1410, A2 => dp_n1400, A3 => dp_n1390,
                           A4 => dp_n1380, Z => dp_n1420);
   dp_U299 : AND2D1 port map( A1 => dp_cmp_l_8_port, A2 => dp_n1470, Z => 
                           dp_n1400);
   dp_U298 : NOR3M1D1 port map( A1 => dp_n1370, A2 => dp_n1360, A3 => dp_n1350,
                           Z => dp_n1430);
   dp_U297 : OAI211D1 port map( A1 => dp_cmp_r_4_port, A2 => dp_n1550, B => 
                           dp_n134, C => dp_n1330, Z => dp_n1360);
   dp_U296 : NAN2D1 port map( A1 => dp_n1320, A2 => dp_n1310, Z => dp_n1330);
   dp_U295 : OAI21D1 port map( A1 => dp_cmp_r_2_port, A2 => dp_n1530, B => 
                           dp_n1300, Z => dp_n1310);
   dp_U294 : OAI211D1 port map( A1 => dp_n1460, A2 => dp_cmp_l_1_port, B => 
                           dp_n1320, C => dp_n1290, Z => dp_n1370);
   dp_U293 : OAI22M10D1 port map( A1 => dp_cmp_l_0_port, A2 => dp_cmp_r_0_port,
                           B1 => dp_n1520, B2 => dp_cmp_r_1_port, Z => dp_n1290
                           );
   dp_U292 : AOI32D1 port map( A1 => dp_cmp_r_2_port, A2 => dp_n1530, A3 => 
                           dp_n1300, B1 => dp_n1540, B2 => dp_cmp_r_3_port, Z 
                           => dp_n1320);
   dp_U291 : OR2D1 port map( A1 => dp_cmp_r_3_port, A2 => dp_n1540, Z => 
                           dp_n1300);
   dp_U290 : AOI22D1 port map( A1 => dp_n1280, A2 => dp_n1270, B1 => dp_n1270, 
                           B2 => dp_n1350, Z => dp_n1440);
   dp_U289 : OAI21D1 port map( A1 => dp_cmp_r_6_port, A2 => dp_n1570, B => 
                           dp_n1260, Z => dp_n1350);
   dp_U288 : AOI32D1 port map( A1 => dp_cmp_r_6_port, A2 => dp_n1570, A3 => 
                           dp_n1260, B1 => dp_n1580, B2 => dp_cmp_r_7_port, Z 
                           => dp_n1270);
   dp_U287 : OR2D1 port map( A1 => dp_cmp_r_7_port, A2 => dp_n1580, Z => 
                           dp_n1260);
   dp_U286 : AOI32D1 port map( A1 => dp_n134, A2 => dp_n1550, A3 => 
                           dp_cmp_r_4_port, B1 => dp_cmp_r_5_port, B2 => 
                           dp_n1560, Z => dp_n1280);
   dp_U285 : NAN2M1D1 port map( A1 => dp_cmp_r_5_port, A2 => dp_cmp_l_5_port, Z
                           => dp_n134);
   dp_U284 : OAI21D1 port map( A1 => dp_n1380, A2 => dp_n1250, B => dp_n1240, Z
                           => dp_n1450);
   dp_U283 : OAI22D1 port map( A1 => dp_n1230, A2 => dp_n1220, B1 => dp_n1220, 
                           B2 => dp_n1210, Z => dp_n1240);
   dp_U282 : AO32D1 port map( A1 => dp_cmp_r_12_port, A2 => dp_n1590, A3 => 
                           dp_n1200, B1 => dp_n1600, B2 => dp_cmp_r_13_port, Z 
                           => dp_n1210);
   dp_U281 : OAI32D1 port map( A1 => dp_n151, A2 => dp_cmp_l_14_port, A3 => 
                           dp_n1190, B1 => dp_cmp_r_15_port, B2 => dp_n1610, Z 
                           => dp_n1220);
   dp_U280 : OAI22D1 port map( A1 => dp_n1410, A2 => dp_n58, B1 => dp_n58, B2 
                           => dp_n57, Z => dp_n1250);
   dp_U279 : OAI32D1 port map( A1 => dp_n1470, A2 => dp_cmp_l_8_port, A3 => 
                           dp_n1390, B1 => dp_cmp_l_9_port, B2 => dp_n1480, Z 
                           => dp_n57);
   dp_U278 : AND2D1 port map( A1 => dp_cmp_l_9_port, A2 => dp_n1480, Z => 
                           dp_n1390);
   dp_U277 : OAI32D1 port map( A1 => dp_n1490, A2 => dp_cmp_l_10_port, A3 => 
                           dp_n56, B1 => dp_cmp_l_11_port, B2 => dp_n1500, Z =>
                           dp_n58);
   dp_U276 : AOI21D1 port map( A1 => dp_n1490, A2 => dp_cmp_l_10_port, B => 
                           dp_n56, Z => dp_n1410);
   dp_U275 : NOR2M1D1 port map( A1 => dp_cmp_l_11_port, A2 => dp_cmp_r_11_port,
                           Z => dp_n56);
   dp_U274 : OAI211D1 port map( A1 => dp_cmp_r_12_port, A2 => dp_n1590, B => 
                           dp_n1200, C => dp_n1230, Z => dp_n1380);
   dp_U273 : AOI21D1 port map( A1 => dp_n151, A2 => dp_cmp_l_14_port, B => 
                           dp_n1190, Z => dp_n1230);
   dp_U272 : NOR2M1D1 port map( A1 => dp_cmp_r_15_port, A2 => dp_cmp_l_15_port,
                           Z => dp_n1190);
   dp_U271 : OR2D1 port map( A1 => dp_cmp_r_13_port, A2 => dp_n1600, Z => 
                           dp_n1200);
   dp_U270 : NAN2D1 port map( A1 => dp_n36, A2 => dp_n35, Z => data_out_15_port
                           );
   dp_U269 : AOI22D1 port map( A1 => dp_mem_63_port, A2 => dp_n34, B1 => 
                           dp_mem_47_port, B2 => dp_n33, Z => dp_n35);
   dp_U268 : AOI22D1 port map( A1 => dp_mem_31_port, A2 => dp_n32, B1 => 
                           dp_mem_15_port, B2 => dp_n31, Z => dp_n36);
   dp_U267 : NAN2D1 port map( A1 => dp_n30, A2 => dp_n29, Z => data_out_14_port
                           );
   dp_U266 : AOI22D1 port map( A1 => dp_mem_62_port, A2 => dp_n34, B1 => 
                           dp_mem_46_port, B2 => dp_n33, Z => dp_n29);
   dp_U265 : AOI22D1 port map( A1 => dp_mem_30_port, A2 => dp_n32, B1 => 
                           dp_mem_14_port, B2 => dp_n31, Z => dp_n30);
   dp_U264 : NAN2D1 port map( A1 => dp_n28, A2 => dp_n27, Z => data_out_13_port
                           );
   dp_U263 : AOI22D1 port map( A1 => dp_mem_61_port, A2 => dp_n34, B1 => 
                           dp_mem_45_port, B2 => dp_n33, Z => dp_n27);
   dp_U262 : AOI22D1 port map( A1 => dp_mem_29_port, A2 => dp_n32, B1 => 
                           dp_mem_13_port, B2 => dp_n31, Z => dp_n28);
   dp_U261 : NAN2D1 port map( A1 => dp_n26, A2 => dp_n25, Z => data_out_12_port
                           );
   dp_U260 : AOI22D1 port map( A1 => dp_mem_60_port, A2 => dp_n34, B1 => 
                           dp_mem_44_port, B2 => dp_n33, Z => dp_n25);
   dp_U259 : AOI22D1 port map( A1 => dp_mem_28_port, A2 => dp_n32, B1 => 
                           dp_mem_12_port, B2 => dp_n31, Z => dp_n26);
   dp_U258 : NAN2D1 port map( A1 => dp_n24, A2 => dp_n23, Z => data_out_11_port
                           );
   dp_U257 : AOI22D1 port map( A1 => dp_mem_59_port, A2 => dp_n34, B1 => 
                           dp_mem_43_port, B2 => dp_n33, Z => dp_n23);
   dp_U256 : AOI22D1 port map( A1 => dp_mem_27_port, A2 => dp_n32, B1 => 
                           dp_mem_11_port, B2 => dp_n31, Z => dp_n24);
   dp_U255 : NAN2D1 port map( A1 => dp_n22, A2 => dp_n21, Z => data_out_10_port
                           );
   dp_U254 : AOI22D1 port map( A1 => dp_mem_58_port, A2 => dp_n34, B1 => 
                           dp_mem_42_port, B2 => dp_n33, Z => dp_n21);
   dp_U253 : AOI22D1 port map( A1 => dp_mem_26_port, A2 => dp_n32, B1 => 
                           dp_mem_10_port, B2 => dp_n31, Z => dp_n22);
   dp_U252 : NAN2D1 port map( A1 => dp_n20, A2 => dp_n1900, Z => 
                           data_out_9_port);
   dp_U251 : AOI22D1 port map( A1 => dp_mem_57_port, A2 => dp_n34, B1 => 
                           dp_mem_41_port, B2 => dp_n33, Z => dp_n1900);
   dp_U250 : AOI22D1 port map( A1 => dp_mem_25_port, A2 => dp_n32, B1 => 
                           dp_mem_9_port, B2 => dp_n31, Z => dp_n20);
   dp_U249 : NAN2D1 port map( A1 => dp_n1800, A2 => dp_n17, Z => 
                           data_out_8_port);
   dp_U248 : AOI22D1 port map( A1 => dp_mem_56_port, A2 => dp_n34, B1 => 
                           dp_mem_40_port, B2 => dp_n33, Z => dp_n17);
   dp_U247 : AOI22D1 port map( A1 => dp_mem_24_port, A2 => dp_n32, B1 => 
                           dp_mem_8_port, B2 => dp_n31, Z => dp_n1800);
   dp_U246 : NAN2D1 port map( A1 => dp_n16, A2 => dp_n15, Z => data_out_7_port)
                           ;
   dp_U245 : AOI22D1 port map( A1 => dp_mem_55_port, A2 => dp_n34, B1 => 
                           dp_mem_39_port, B2 => dp_n33, Z => dp_n15);
   dp_U244 : AOI22D1 port map( A1 => dp_mem_23_port, A2 => dp_n32, B1 => 
                           dp_mem_7_port, B2 => dp_n31, Z => dp_n16);
   dp_U243 : NAN2D1 port map( A1 => dp_n14, A2 => dp_n13, Z => data_out_6_port)
                           ;
   dp_U242 : AOI22D1 port map( A1 => dp_mem_54_port, A2 => dp_n34, B1 => 
                           dp_mem_38_port, B2 => dp_n33, Z => dp_n13);
   dp_U241 : AOI22D1 port map( A1 => dp_mem_22_port, A2 => dp_n32, B1 => 
                           dp_mem_6_port, B2 => dp_n31, Z => dp_n14);
   dp_U240 : NAN2D1 port map( A1 => dp_n12, A2 => dp_n11, Z => data_out_5_port)
                           ;
   dp_U239 : AOI22D1 port map( A1 => dp_mem_53_port, A2 => dp_n34, B1 => 
                           dp_mem_37_port, B2 => dp_n33, Z => dp_n11);
   dp_U238 : AOI22D1 port map( A1 => dp_mem_21_port, A2 => dp_n32, B1 => 
                           dp_mem_5_port, B2 => dp_n31, Z => dp_n12);
   dp_U237 : NAN2D1 port map( A1 => dp_n10, A2 => dp_n9, Z => data_out_4_port);
   dp_U236 : AOI22D1 port map( A1 => dp_mem_52_port, A2 => dp_n34, B1 => 
                           dp_mem_36_port, B2 => dp_n33, Z => dp_n9);
   dp_U235 : AOI22D1 port map( A1 => dp_mem_20_port, A2 => dp_n32, B1 => 
                           dp_mem_4_port, B2 => dp_n31, Z => dp_n10);
   dp_U234 : NAN2D1 port map( A1 => dp_n8, A2 => dp_n7, Z => data_out_3_port);
   dp_U233 : AOI22D1 port map( A1 => dp_mem_51_port, A2 => dp_n34, B1 => 
                           dp_mem_35_port, B2 => dp_n33, Z => dp_n7);
   dp_U232 : AOI22D1 port map( A1 => dp_mem_19_port, A2 => dp_n32, B1 => 
                           dp_mem_3_port, B2 => dp_n31, Z => dp_n8);
   dp_U231 : NAN2D1 port map( A1 => dp_n6, A2 => dp_n5, Z => data_out_2_port);
   dp_U230 : AOI22D1 port map( A1 => dp_mem_50_port, A2 => dp_n34, B1 => 
                           dp_mem_34_port, B2 => dp_n33, Z => dp_n5);
   dp_U229 : AOI22D1 port map( A1 => dp_mem_18_port, A2 => dp_n32, B1 => 
                           dp_mem_2_port, B2 => dp_n31, Z => dp_n6);
   dp_U228 : NAN2D1 port map( A1 => dp_n4, A2 => dp_n3, Z => data_out_1_port);
   dp_U227 : AOI22D1 port map( A1 => dp_mem_49_port, A2 => dp_n34, B1 => 
                           dp_mem_33_port, B2 => dp_n33, Z => dp_n3);
   dp_U226 : AOI22D1 port map( A1 => dp_mem_17_port, A2 => dp_n32, B1 => 
                           dp_mem_1_port, B2 => dp_n31, Z => dp_n4);
   dp_U225 : NAN2D1 port map( A1 => dp_n2, A2 => dp_n1, Z => data_out_0_port);
   dp_U224 : AOI22D1 port map( A1 => dp_mem_48_port, A2 => dp_n34, B1 => 
                           dp_mem_32_port, B2 => dp_n33, Z => dp_n1);
   dp_U223 : AOI22D1 port map( A1 => dp_mem_16_port, A2 => dp_n32, B1 => 
                           dp_mem_0_port, B2 => dp_n31, Z => dp_n2);
   dp_U222 : INVD1 port map( A => n1, Z => dp_n186);
   dp_U221 : NAN3D1 port map( A1 => wr_addr_0, A2 => dp_n76, A3 => n1, Z => 
                           dp_n79);
   dp_U220 : NAN3D1 port map( A1 => dp_n76, A2 => dp_n1620, A3 => n1, Z => 
                           dp_n78);
   dp_U219 : INVD1 port map( A => dp_add_out_15_port, Z => dp_n187);
   dp_U218 : INVD1 port map( A => dp_cmp_r_1_port, Z => dp_n1460);
   dp_U217 : INVD1 port map( A => dp_cmp_l_4_port, Z => dp_n1550);
   dp_U216 : INVD1 port map( A => dp_cmp_r_8_port, Z => dp_n1470);
   dp_U215 : INVD1 port map( A => dp_cmp_l_6_port, Z => dp_n1570);
   dp_U214 : INVD1 port map( A => dp_cmp_r_14_port, Z => dp_n151);
   dp_U213 : NAN4D1 port map( A1 => dp_n1030, A2 => dp_n1040, A3 => dp_n1050, 
                           A4 => dp_n1060, Z => dp_n1020);
   dp_U212 : INVD1 port map( A => dp_cmp_l_1_port, Z => dp_n1520);
   dp_U211 : INVD1 port map( A => dp_cmp_r_10_port, Z => dp_n1490);
   dp_U210 : INVD1 port map( A => dp_cmp_l_5_port, Z => dp_n1560);
   dp_U209 : INVD1 port map( A => dp_cmp_l_12_port, Z => dp_n1590);
   dp_U208 : INVD1 port map( A => dp_cmp_l_2_port, Z => dp_n1530);
   dp_U207 : INVD1 port map( A => dp_cmp_r_9_port, Z => dp_n1480);
   dp_U206 : INVD1 port map( A => dp_cmp_l_7_port, Z => dp_n1580);
   dp_U205 : INVD1 port map( A => dp_cmp_r_11_port, Z => dp_n1500);
   dp_U204 : INVD1 port map( A => dp_cmp_l_13_port, Z => dp_n1600);
   dp_U203 : INVD1 port map( A => dp_cmp_l_15_port, Z => dp_n1610);
   dp_U202 : INVD1 port map( A => dp_cmp_l_3_port, Z => dp_n1540);
   dp_U201 : INVD1 port map( A => reset, Z => dp_n40);
   dp_U200 : INVD1 port map( A => dp_add_out_0_port, Z => dp_n2020);
   dp_U199 : INVD1 port map( A => dp_add_out_1_port, Z => dp_n2010);
   dp_U198 : INVD1 port map( A => dp_add_out_2_port, Z => dp_n200);
   dp_U197 : INVD1 port map( A => dp_add_out_3_port, Z => dp_n199);
   dp_U196 : INVD1 port map( A => dp_add_out_4_port, Z => dp_n198);
   dp_U195 : INVD1 port map( A => dp_add_out_5_port, Z => dp_n197);
   dp_U194 : INVD1 port map( A => dp_add_out_6_port, Z => dp_n196);
   dp_U193 : INVD1 port map( A => data_out_0_port, Z => dp_n170);
   dp_U192 : INVD1 port map( A => data_out_1_port, Z => dp_n171);
   dp_U191 : INVD1 port map( A => data_out_2_port, Z => dp_n172);
   dp_U190 : INVD1 port map( A => data_out_3_port, Z => dp_n173);
   dp_U189 : INVD1 port map( A => data_out_4_port, Z => dp_n174);
   dp_U59 : INVD1 port map( A => data_out_5_port, Z => dp_n175);
   dp_U58 : INVD1 port map( A => data_out_6_port, Z => dp_n176);
   dp_U57 : INVD1 port map( A => data_out_7_port, Z => dp_n177);
   dp_U56 : INVD1 port map( A => data_out_8_port, Z => dp_n178);
   dp_U55 : INVD1 port map( A => data_out_9_port, Z => dp_n179);
   dp_U54 : INVD1 port map( A => data_out_10_port, Z => dp_n1801);
   dp_U53 : INVD1 port map( A => data_out_11_port, Z => dp_n181);
   dp_U52 : INVD1 port map( A => data_out_12_port, Z => dp_n182);
   dp_U51 : INVD1 port map( A => data_out_13_port, Z => dp_n183);
   dp_U50 : INVD1 port map( A => data_out_14_port, Z => dp_n184);
   dp_U49 : INVD1 port map( A => data_out_15_port, Z => dp_n185);
   dp_U48 : INVD1 port map( A => dp_add_out_7_port, Z => dp_n195);
   dp_U47 : INVD1 port map( A => dp_add_out_8_port, Z => dp_n194);
   dp_U46 : NAN2D1 port map( A1 => wr_sel_en_1_port, A2 => wr_sel_en_0_port, Z 
                           => dp_n98);
   dp_U45 : INVD1 port map( A => dp_add_out_9_port, Z => dp_n193);
   dp_U44 : NAN2M1D1 port map( A1 => wr_sel_en_1_port, A2 => wr_sel_en_0_port, 
                           Z => dp_n80);
   dp_U43 : NAN3D1 port map( A1 => dp_n76, A2 => dp_n186, A3 => wr_addr_0, Z =>
                           dp_n77);
   dp_U42 : NOR2M1D1 port map( A1 => wr_sel_en_1_port, A2 => wr_sel_en_0_port, 
                           Z => dp_n82);
   dp_U41 : NAN3D1 port map( A1 => dp_n1620, A2 => dp_n186, A3 => dp_n76, Z => 
                           dp_n59);
   dp_U40 : INVD1 port map( A => dp_add_out_10_port, Z => dp_n192);
   dp_U39 : INVD1 port map( A => dp_add_out_11_port, Z => dp_n191);
   dp_U38 : INVD1 port map( A => dp_add_out_12_port, Z => dp_n1901);
   dp_U37 : INVD1 port map( A => dp_add_out_13_port, Z => dp_n189);
   dp_U36 : INVD1 port map( A => dp_add_out_14_port, Z => dp_n188);
   dp_U35 : NAN4D1 port map( A1 => dp_n1070, A2 => dp_n1080, A3 => dp_n1090, A4
                           => dp_n1100, Z => dp_n1010);
   dp_U34 : NAN4D1 port map( A1 => dp_n1110, A2 => dp_n1120, A3 => dp_n1130, A4
                           => dp_n1140, Z => dp_n100);
   dp_U33 : NAN4D1 port map( A1 => dp_n1150, A2 => dp_n1160, A3 => dp_n117, A4 
                           => dp_n1180, Z => dp_n99);
   dp_U32 : NOR4D1 port map( A1 => dp_n99, A2 => dp_n100, A3 => dp_n1010, A4 =>
                           dp_n1020, Z => equal);
   dp_U31 : INVD1 port map( A => reset, Z => dp_n49);
   dp_U30 : INVD1 port map( A => reset, Z => dp_n48);
   dp_U29 : INVD1 port map( A => reset, Z => dp_n47);
   dp_U28 : INVD1 port map( A => reset, Z => dp_n46);
   dp_U27 : INVD1 port map( A => reset, Z => dp_n45);
   dp_U26 : INVD1 port map( A => reset, Z => dp_n44);
   dp_U25 : INVD1 port map( A => reset, Z => dp_n43);
   dp_U24 : INVD1 port map( A => reset, Z => dp_n42);
   dp_U23 : INVD1 port map( A => reset, Z => dp_n41);
   dp_U22 : INVD1 port map( A => cmp_l_en, Z => dp_n168);
   dp_U21 : INVD1 port map( A => add_l_en, Z => dp_n169);
   dp_U20 : INVD1 port map( A => add_l_sel, Z => dp_n55);
   dp_U19 : INVD1 port map( A => add_l_sel, Z => dp_n52);
   dp_U18 : INVD1 port map( A => dp_n98, Z => dp_n1630);
   dp_U17 : NOR2D1 port map( A1 => rd_addr_0_port, A2 => rd_addr_1_port, Z => 
                           dp_n34);
   dp_U16 : NOR2D1 port map( A1 => dp_n37, A2 => rd_addr_0_port, Z => dp_n32);
   dp_U15 : INVD1 port map( A => rd_addr_0_port, Z => dp_n38);
   dp_U14 : INVD1 port map( A => cmp_r_en, Z => dp_n1660);
   dp_U13 : INVD1 port map( A => add_r_en, Z => dp_n1670);
   dp_U12 : BUFD1 port map( A => cmp_r_sel, Z => dp_n39);
   dp_U11 : INVD1 port map( A => wr_addr_0, Z => dp_n1620);
   dp_U10 : INVD1 port map( A => dp_n55, Z => dp_n54);
   dp_U9 : INVD1 port map( A => dp_n52, Z => dp_n51);
   dp_U8 : INVD1 port map( A => dp_n52, Z => dp_n50);
   dp_U7 : NOR2D1 port map( A1 => dp_n38, A2 => rd_addr_1_port, Z => dp_n33);
   dp_U6 : NOR2D1 port map( A1 => dp_n37, A2 => dp_n38, Z => dp_n31);
   dp_U5 : INVD1 port map( A => dp_n39, Z => dp_n1640);
   dp_U4 : INVD1 port map( A => dp_n50, Z => dp_n53);
   dp_U3 : INVD1 port map( A => add_r_sel, Z => dp_n1650);
   dp_U2 : INVD1 port map( A => rd_addr_1_port, Z => dp_n37);
   dp_cmp_l_reg_3 : DFERPQ1 port map( D => dp_N138, CEB => dp_n168, CK => clk, 
                           RB => dp_n41, Q => dp_cmp_l_3_port);
   dp_cmp_l_reg_13 : DFERPQ1 port map( D => dp_N148, CEB => dp_n168, CK => clk,
                           RB => dp_n42, Q => dp_cmp_l_13_port);
   dp_cmp_r_reg_3 : DFERPQ1 port map( D => dp_N155, CEB => dp_n1660, CK => clk,
                           RB => dp_n40, Q => dp_cmp_r_3_port);
   dp_cmp_l_reg_11 : DFERPQ1 port map( D => dp_N146, CEB => dp_n168, CK => clk,
                           RB => dp_n42, Q => dp_cmp_l_11_port);
   dp_cmp_r_reg_15 : DFERPQ1 port map( D => dp_N167, CEB => dp_n1660, CK => clk
                           , RB => dp_n41, Q => dp_cmp_r_15_port);
   dp_cmp_r_reg_13 : DFERPQ1 port map( D => dp_N165, CEB => dp_n1660, CK => clk
                           , RB => dp_n41, Q => dp_cmp_r_13_port);
   dp_cmp_l_reg_7 : DFERPQ1 port map( D => dp_N142, CEB => dp_n168, CK => clk, 
                           RB => dp_n41, Q => dp_cmp_l_7_port);
   dp_cmp_r_reg_11 : DFERPQ1 port map( D => dp_N163, CEB => dp_n1660, CK => clk
                           , RB => dp_n40, Q => dp_cmp_r_11_port);
   dp_cmp_r_reg_9 : DFERPQ1 port map( D => dp_N161, CEB => dp_n1660, CK => clk,
                           RB => dp_n40, Q => dp_cmp_r_9_port);
   dp_cmp_l_reg_15 : DFERPQ1 port map( D => dp_N150, CEB => dp_n168, CK => clk,
                           RB => dp_n42, Q => dp_cmp_l_15_port);
   dp_cmp_l_reg_2 : DFERPQ1 port map( D => dp_N137, CEB => dp_n168, CK => clk, 
                           RB => dp_n41, Q => dp_cmp_l_2_port);
   dp_cmp_r_reg_7 : DFERPQ1 port map( D => dp_N159, CEB => dp_n1660, CK => clk,
                           RB => dp_n40, Q => dp_cmp_r_7_port);
   dp_cmp_l_reg_9 : DFERPQ1 port map( D => dp_N144, CEB => dp_n168, CK => clk, 
                           RB => dp_n41, Q => dp_cmp_l_9_port);
   dp_cmp_l_reg_12 : DFERPQ1 port map( D => dp_N147, CEB => dp_n168, CK => clk,
                           RB => dp_n42, Q => dp_cmp_l_12_port);
   dp_cmp_r_reg_2 : DFERPQ1 port map( D => dp_N154, CEB => dp_n1660, CK => clk,
                           RB => dp_n40, Q => dp_cmp_r_2_port);
   dp_cmp_r_reg_5 : DFERPQ1 port map( D => dp_N157, CEB => dp_n1660, CK => clk,
                           RB => dp_n40, Q => dp_cmp_r_5_port);
   dp_cmp_r_reg_10 : DFERPQ1 port map( D => dp_N162, CEB => dp_n1660, CK => clk
                           , RB => dp_n40, Q => dp_cmp_r_10_port);
   dp_cmp_l_reg_0 : DFERPQ1 port map( D => dp_N135, CEB => dp_n168, CK => clk, 
                           RB => dp_n41, Q => dp_cmp_l_0_port);
   dp_cmp_l_reg_1 : DFERPQ1 port map( D => dp_N136, CEB => dp_n168, CK => clk, 
                           RB => dp_n41, Q => dp_cmp_l_1_port);
   dp_cmp_l_reg_10 : DFERPQ1 port map( D => dp_N145, CEB => dp_n168, CK => clk,
                           RB => dp_n42, Q => dp_cmp_l_10_port);
   dp_cmp_r_reg_12 : DFERPQ1 port map( D => dp_N164, CEB => dp_n1660, CK => clk
                           , RB => dp_n40, Q => dp_cmp_r_12_port);
   dp_cmp_r_reg_0 : DFERPQ1 port map( D => dp_N152, CEB => dp_n1660, CK => clk,
                           RB => dp_n40, Q => dp_cmp_r_0_port);
   dp_cmp_r_reg_14 : DFERPQ1 port map( D => dp_N166, CEB => dp_n1660, CK => clk
                           , RB => dp_n41, Q => dp_cmp_r_14_port);
   dp_cmp_r_reg_1 : DFERPQ1 port map( D => dp_N153, CEB => dp_n1660, CK => clk,
                           RB => dp_n40, Q => dp_cmp_r_1_port);
   dp_cmp_l_reg_6 : DFERPQ1 port map( D => dp_N141, CEB => dp_n168, CK => clk, 
                           RB => dp_n41, Q => dp_cmp_l_6_port);
   dp_cmp_l_reg_5 : DFERPQ1 port map( D => dp_N140, CEB => dp_n168, CK => clk, 
                           RB => dp_n41, Q => dp_cmp_l_5_port);
   dp_cmp_l_reg_14 : DFERPQ1 port map( D => dp_N149, CEB => dp_n168, CK => clk,
                           RB => dp_n42, Q => dp_cmp_l_14_port);
   dp_cmp_r_reg_8 : DFERPQ1 port map( D => dp_N160, CEB => dp_n1660, CK => clk,
                           RB => dp_n40, Q => dp_cmp_r_8_port);
   dp_cmp_l_reg_4 : DFERPQ1 port map( D => dp_N139, CEB => dp_n168, CK => clk, 
                           RB => dp_n41, Q => dp_cmp_l_4_port);
   dp_cmp_l_reg_8 : DFERPQ1 port map( D => dp_N143, CEB => dp_n168, CK => clk, 
                           RB => dp_n41, Q => dp_cmp_l_8_port);
   dp_cmp_r_reg_6 : DFERPQ1 port map( D => dp_N158, CEB => dp_n1660, CK => clk,
                           RB => dp_n40, Q => dp_cmp_r_6_port);
   dp_cmp_r_reg_4 : DFERPQ1 port map( D => dp_N156, CEB => dp_n1660, CK => clk,
                           RB => dp_n40, Q => dp_cmp_r_4_port);
   dp_mem_reg_0_15 : DFERPQ1 port map( D => dp_n60, CEB => dp_n59, CK => clk, 
                           RB => dp_n42, Q => dp_mem_63_port);
   dp_mem_reg_0_14 : DFERPQ1 port map( D => dp_n61, CEB => dp_n59, CK => clk, 
                           RB => dp_n43, Q => dp_mem_62_port);
   dp_mem_reg_0_13 : DFERPQ1 port map( D => dp_n62, CEB => dp_n59, CK => clk, 
                           RB => dp_n43, Q => dp_mem_61_port);
   dp_mem_reg_0_12 : DFERPQ1 port map( D => dp_n63, CEB => dp_n59, CK => clk, 
                           RB => dp_n44, Q => dp_mem_60_port);
   dp_mem_reg_0_11 : DFERPQ1 port map( D => dp_n64, CEB => dp_n59, CK => clk, 
                           RB => dp_n44, Q => dp_mem_59_port);
   dp_mem_reg_0_10 : DFERPQ1 port map( D => dp_n65, CEB => dp_n59, CK => clk, 
                           RB => dp_n45, Q => dp_mem_58_port);
   dp_mem_reg_0_9 : DFERPQ1 port map( D => dp_n66, CEB => dp_n59, CK => clk, RB
                           => dp_n45, Q => dp_mem_57_port);
   dp_mem_reg_0_8 : DFERPQ1 port map( D => dp_n67, CEB => dp_n59, CK => clk, RB
                           => dp_n45, Q => dp_mem_56_port);
   dp_mem_reg_0_7 : DFERPQ1 port map( D => dp_n68, CEB => dp_n59, CK => clk, RB
                           => dp_n46, Q => dp_mem_55_port);
   dp_mem_reg_0_6 : DFERPQ1 port map( D => dp_n69, CEB => dp_n59, CK => clk, RB
                           => dp_n46, Q => dp_mem_54_port);
   dp_mem_reg_0_5 : DFERPQ1 port map( D => dp_n70, CEB => dp_n59, CK => clk, RB
                           => dp_n47, Q => dp_mem_53_port);
   dp_mem_reg_0_4 : DFERPQ1 port map( D => dp_n71, CEB => dp_n59, CK => clk, RB
                           => dp_n47, Q => dp_mem_52_port);
   dp_mem_reg_0_3 : DFERPQ1 port map( D => dp_n72, CEB => dp_n59, CK => clk, RB
                           => dp_n48, Q => dp_mem_51_port);
   dp_mem_reg_0_2 : DFERPQ1 port map( D => dp_n73, CEB => dp_n59, CK => clk, RB
                           => dp_n48, Q => dp_mem_50_port);
   dp_mem_reg_0_1 : DFERPQ1 port map( D => dp_n74, CEB => dp_n59, CK => clk, RB
                           => dp_n49, Q => dp_mem_49_port);
   dp_mem_reg_0_0 : DFERPQ1 port map( D => dp_n75, CEB => dp_n59, CK => clk, RB
                           => dp_n49, Q => dp_mem_48_port);
   dp_mem_reg_2_15 : DFERPQ1 port map( D => dp_n60, CEB => dp_n78, CK => clk, 
                           RB => dp_n42, Q => dp_mem_31_port);
   dp_mem_reg_2_14 : DFERPQ1 port map( D => dp_n61, CEB => dp_n78, CK => clk, 
                           RB => dp_n43, Q => dp_mem_30_port);
   dp_mem_reg_2_13 : DFERPQ1 port map( D => dp_n62, CEB => dp_n78, CK => clk, 
                           RB => dp_n43, Q => dp_mem_29_port);
   dp_mem_reg_2_12 : DFERPQ1 port map( D => dp_n63, CEB => dp_n78, CK => clk, 
                           RB => dp_n43, Q => dp_mem_28_port);
   dp_mem_reg_2_11 : DFERPQ1 port map( D => dp_n64, CEB => dp_n78, CK => clk, 
                           RB => dp_n44, Q => dp_mem_27_port);
   dp_mem_reg_2_10 : DFERPQ1 port map( D => dp_n65, CEB => dp_n78, CK => clk, 
                           RB => dp_n44, Q => dp_mem_26_port);
   dp_mem_reg_2_9 : DFERPQ1 port map( D => dp_n66, CEB => dp_n78, CK => clk, RB
                           => dp_n45, Q => dp_mem_25_port);
   dp_mem_reg_2_8 : DFERPQ1 port map( D => dp_n67, CEB => dp_n78, CK => clk, RB
                           => dp_n45, Q => dp_mem_24_port);
   dp_mem_reg_2_7 : DFERPQ1 port map( D => dp_n68, CEB => dp_n78, CK => clk, RB
                           => dp_n46, Q => dp_mem_23_port);
   dp_mem_reg_2_6 : DFERPQ1 port map( D => dp_n69, CEB => dp_n78, CK => clk, RB
                           => dp_n46, Q => dp_mem_22_port);
   dp_mem_reg_2_5 : DFERPQ1 port map( D => dp_n70, CEB => dp_n78, CK => clk, RB
                           => dp_n47, Q => dp_mem_21_port);
   dp_mem_reg_2_4 : DFERPQ1 port map( D => dp_n71, CEB => dp_n78, CK => clk, RB
                           => dp_n47, Q => dp_mem_20_port);
   dp_mem_reg_2_3 : DFERPQ1 port map( D => dp_n72, CEB => dp_n78, CK => clk, RB
                           => dp_n48, Q => dp_mem_19_port);
   dp_mem_reg_2_2 : DFERPQ1 port map( D => dp_n73, CEB => dp_n78, CK => clk, RB
                           => dp_n48, Q => dp_mem_18_port);
   dp_mem_reg_2_1 : DFERPQ1 port map( D => dp_n74, CEB => dp_n78, CK => clk, RB
                           => dp_n49, Q => dp_mem_17_port);
   dp_mem_reg_2_0 : DFERPQ1 port map( D => dp_n75, CEB => dp_n78, CK => clk, RB
                           => dp_n49, Q => dp_mem_16_port);
   dp_mem_reg_1_15 : DFERPQ1 port map( D => dp_n60, CEB => dp_n77, CK => clk, 
                           RB => dp_n42, Q => dp_mem_47_port);
   dp_mem_reg_1_14 : DFERPQ1 port map( D => dp_n61, CEB => dp_n77, CK => clk, 
                           RB => dp_n43, Q => dp_mem_46_port);
   dp_mem_reg_1_13 : DFERPQ1 port map( D => dp_n62, CEB => dp_n77, CK => clk, 
                           RB => dp_n43, Q => dp_mem_45_port);
   dp_mem_reg_1_12 : DFERPQ1 port map( D => dp_n63, CEB => dp_n77, CK => clk, 
                           RB => dp_n44, Q => dp_mem_44_port);
   dp_mem_reg_1_11 : DFERPQ1 port map( D => dp_n64, CEB => dp_n77, CK => clk, 
                           RB => dp_n44, Q => dp_mem_43_port);
   dp_mem_reg_1_10 : DFERPQ1 port map( D => dp_n65, CEB => dp_n77, CK => clk, 
                           RB => dp_n44, Q => dp_mem_42_port);
   dp_mem_reg_1_9 : DFERPQ1 port map( D => dp_n66, CEB => dp_n77, CK => clk, RB
                           => dp_n45, Q => dp_mem_41_port);
   dp_mem_reg_1_8 : DFERPQ1 port map( D => dp_n67, CEB => dp_n77, CK => clk, RB
                           => dp_n45, Q => dp_mem_40_port);
   dp_mem_reg_1_7 : DFERPQ1 port map( D => dp_n68, CEB => dp_n77, CK => clk, RB
                           => dp_n46, Q => dp_mem_39_port);
   dp_mem_reg_1_6 : DFERPQ1 port map( D => dp_n69, CEB => dp_n77, CK => clk, RB
                           => dp_n46, Q => dp_mem_38_port);
   dp_mem_reg_1_5 : DFERPQ1 port map( D => dp_n70, CEB => dp_n77, CK => clk, RB
                           => dp_n47, Q => dp_mem_37_port);
   dp_mem_reg_1_4 : DFERPQ1 port map( D => dp_n71, CEB => dp_n77, CK => clk, RB
                           => dp_n47, Q => dp_mem_36_port);
   dp_mem_reg_1_3 : DFERPQ1 port map( D => dp_n72, CEB => dp_n77, CK => clk, RB
                           => dp_n48, Q => dp_mem_35_port);
   dp_mem_reg_1_2 : DFERPQ1 port map( D => dp_n73, CEB => dp_n77, CK => clk, RB
                           => dp_n48, Q => dp_mem_34_port);
   dp_mem_reg_1_1 : DFERPQ1 port map( D => dp_n74, CEB => dp_n77, CK => clk, RB
                           => dp_n49, Q => dp_mem_33_port);
   dp_mem_reg_1_0 : DFERPQ1 port map( D => dp_n75, CEB => dp_n77, CK => clk, RB
                           => dp_n49, Q => dp_mem_32_port);
   dp_mem_reg_3_15 : DFERPQ1 port map( D => dp_n60, CEB => dp_n79, CK => clk, 
                           RB => dp_n42, Q => dp_mem_15_port);
   dp_mem_reg_3_14 : DFERPQ1 port map( D => dp_n61, CEB => dp_n79, CK => clk, 
                           RB => dp_n42, Q => dp_mem_14_port);
   dp_mem_reg_3_13 : DFERPQ1 port map( D => dp_n62, CEB => dp_n79, CK => clk, 
                           RB => dp_n43, Q => dp_mem_13_port);
   dp_mem_reg_3_12 : DFERPQ1 port map( D => dp_n63, CEB => dp_n79, CK => clk, 
                           RB => dp_n43, Q => dp_mem_12_port);
   dp_mem_reg_3_11 : DFERPQ1 port map( D => dp_n64, CEB => dp_n79, CK => clk, 
                           RB => dp_n44, Q => dp_mem_11_port);
   dp_mem_reg_3_10 : DFERPQ1 port map( D => dp_n65, CEB => dp_n79, CK => clk, 
                           RB => dp_n44, Q => dp_mem_10_port);
   dp_mem_reg_3_9 : DFERPQ1 port map( D => dp_n66, CEB => dp_n79, CK => clk, RB
                           => dp_n45, Q => dp_mem_9_port);
   dp_mem_reg_3_8 : DFERPQ1 port map( D => dp_n67, CEB => dp_n79, CK => clk, RB
                           => dp_n45, Q => dp_mem_8_port);
   dp_mem_reg_3_7 : DFERPQ1 port map( D => dp_n68, CEB => dp_n79, CK => clk, RB
                           => dp_n46, Q => dp_mem_7_port);
   dp_mem_reg_3_6 : DFERPQ1 port map( D => dp_n69, CEB => dp_n79, CK => clk, RB
                           => dp_n46, Q => dp_mem_6_port);
   dp_mem_reg_3_5 : DFERPQ1 port map( D => dp_n70, CEB => dp_n79, CK => clk, RB
                           => dp_n47, Q => dp_mem_5_port);
   dp_mem_reg_3_4 : DFERPQ1 port map( D => dp_n71, CEB => dp_n79, CK => clk, RB
                           => dp_n47, Q => dp_mem_4_port);
   dp_mem_reg_3_3 : DFERPQ1 port map( D => dp_n72, CEB => dp_n79, CK => clk, RB
                           => dp_n48, Q => dp_mem_3_port);
   dp_mem_reg_3_2 : DFERPQ1 port map( D => dp_n73, CEB => dp_n79, CK => clk, RB
                           => dp_n48, Q => dp_mem_2_port);
   dp_mem_reg_3_1 : DFERPQ1 port map( D => dp_n74, CEB => dp_n79, CK => clk, RB
                           => dp_n48, Q => dp_mem_1_port);
   dp_mem_reg_3_0 : DFERPQ1 port map( D => dp_n75, CEB => dp_n79, CK => clk, RB
                           => dp_n49, Q => dp_mem_0_port);
   dp_add_r_reg_0 : DFERPQ1 port map( D => dp_N118, CEB => dp_n1670, CK => clk,
                           RB => dp_n49, Q => dp_add_r_0_port);
   dp_add_r_reg_1 : DFERPQ1 port map( D => dp_N119, CEB => dp_n1670, CK => clk,
                           RB => dp_n49, Q => dp_add_r_1_port);
   dp_add_l_reg_0 : DFERPQ1 port map( D => dp_N101, CEB => dp_n169, CK => clk, 
                           RB => dp_n49, Q => dp_add_l_0_port);
   dp_add_r_reg_2 : DFERPQ1 port map( D => dp_N120, CEB => dp_n1670, CK => clk,
                           RB => dp_n48, Q => dp_add_r_2_port);
   dp_add_l_reg_1 : DFERPQ1 port map( D => dp_N102, CEB => dp_n169, CK => clk, 
                           RB => dp_n49, Q => dp_add_l_1_port);
   dp_add_r_reg_3 : DFERPQ1 port map( D => dp_N121, CEB => dp_n1670, CK => clk,
                           RB => dp_n48, Q => dp_add_r_3_port);
   dp_add_l_reg_2 : DFERPQ1 port map( D => dp_N103, CEB => dp_n169, CK => clk, 
                           RB => dp_n48, Q => dp_add_l_2_port);
   dp_add_r_reg_4 : DFERPQ1 port map( D => dp_N122, CEB => dp_n1670, CK => clk,
                           RB => dp_n47, Q => dp_add_r_4_port);
   dp_add_l_reg_3 : DFERPQ1 port map( D => dp_N104, CEB => dp_n169, CK => clk, 
                           RB => dp_n48, Q => dp_add_l_3_port);
   dp_add_r_reg_5 : DFERPQ1 port map( D => dp_N123, CEB => dp_n1670, CK => clk,
                           RB => dp_n47, Q => dp_add_r_5_port);
   dp_add_l_reg_4 : DFERPQ1 port map( D => dp_N105, CEB => dp_n169, CK => clk, 
                           RB => dp_n47, Q => dp_add_l_4_port);
   dp_add_r_reg_6 : DFERPQ1 port map( D => dp_N124, CEB => dp_n1670, CK => clk,
                           RB => dp_n46, Q => dp_add_r_6_port);
   dp_add_l_reg_5 : DFERPQ1 port map( D => dp_N106, CEB => dp_n169, CK => clk, 
                           RB => dp_n47, Q => dp_add_l_5_port);
   dp_add_r_reg_7 : DFERPQ1 port map( D => dp_N125, CEB => dp_n1670, CK => clk,
                           RB => dp_n46, Q => dp_add_r_7_port);
   dp_add_l_reg_6 : DFERPQ1 port map( D => dp_N107, CEB => dp_n169, CK => clk, 
                           RB => dp_n47, Q => dp_add_l_6_port);
   dp_add_r_reg_8 : DFERPQ1 port map( D => dp_N126, CEB => dp_n1670, CK => clk,
                           RB => dp_n46, Q => dp_add_r_8_port);
   dp_add_l_reg_7 : DFERPQ1 port map( D => dp_N108, CEB => dp_n169, CK => clk, 
                           RB => dp_n46, Q => dp_add_l_7_port);
   dp_add_r_reg_9 : DFERPQ1 port map( D => dp_N127, CEB => dp_n1670, CK => clk,
                           RB => dp_n45, Q => dp_add_r_9_port);
   dp_add_l_reg_8 : DFERPQ1 port map( D => dp_N109, CEB => dp_n169, CK => clk, 
                           RB => dp_n46, Q => dp_add_l_8_port);
   dp_add_r_reg_10 : DFERPQ1 port map( D => dp_N128, CEB => dp_n1670, CK => clk
                           , RB => dp_n45, Q => dp_add_r_10_port);
   dp_add_l_reg_9 : DFERPQ1 port map( D => dp_N110, CEB => dp_n169, CK => clk, 
                           RB => dp_n45, Q => dp_add_l_9_port);
   dp_add_r_reg_11 : DFERPQ1 port map( D => dp_N129, CEB => dp_n1670, CK => clk
                           , RB => dp_n44, Q => dp_add_r_11_port);
   dp_add_l_reg_10 : DFERPQ1 port map( D => dp_N111, CEB => dp_n169, CK => clk,
                           RB => dp_n45, Q => dp_add_l_10_port);
   dp_add_r_reg_12 : DFERPQ1 port map( D => dp_N130, CEB => dp_n1670, CK => clk
                           , RB => dp_n44, Q => dp_add_r_12_port);
   dp_add_l_reg_11 : DFERPQ1 port map( D => dp_N112, CEB => dp_n169, CK => clk,
                           RB => dp_n44, Q => dp_add_l_11_port);
   dp_add_r_reg_13 : DFERPQ1 port map( D => dp_N131, CEB => dp_n1670, CK => clk
                           , RB => dp_n43, Q => dp_add_r_13_port);
   dp_add_l_reg_12 : DFERPQ1 port map( D => dp_N113, CEB => dp_n169, CK => clk,
                           RB => dp_n44, Q => dp_add_l_12_port);
   dp_add_r_reg_14 : DFERPQ1 port map( D => dp_N132, CEB => dp_n1670, CK => clk
                           , RB => dp_n43, Q => dp_add_r_14_port);
   dp_add_l_reg_13 : DFERPQ1 port map( D => dp_N114, CEB => dp_n169, CK => clk,
                           RB => dp_n43, Q => dp_add_l_13_port);
   dp_add_r_reg_15 : DFERPQ1 port map( D => dp_N133, CEB => dp_n1670, CK => clk
                           , RB => dp_n42, Q => dp_add_r_15_port);
   dp_add_l_reg_14 : DFERPQ1 port map( D => dp_N115, CEB => dp_n169, CK => clk,
                           RB => dp_n43, Q => dp_add_l_14_port);
   dp_add_l_reg_15 : DFERPQ1 port map( D => dp_N116, CEB => dp_n169, CK => clk,
                           RB => dp_n42, Q => dp_add_l_15_port);
   dp_U188 : OAI22D1 port map( A1 => dp_n2020, A2 => dp_n55, B1 => dp_n54, B2 
                           => dp_n170, Z => dp_N101);
   dp_U187 : OAI22D1 port map( A1 => dp_n2010, A2 => dp_n55, B1 => add_l_sel, 
                           B2 => dp_n171, Z => dp_N102);
   dp_U186 : OAI22D1 port map( A1 => dp_n200, A2 => dp_n55, B1 => add_l_sel, B2
                           => dp_n172, Z => dp_N103);
   dp_U185 : OAI22D1 port map( A1 => dp_n199, A2 => dp_n55, B1 => add_l_sel, B2
                           => dp_n173, Z => dp_N104);
   dp_U184 : OAI22D1 port map( A1 => dp_n198, A2 => dp_n55, B1 => dp_n54, B2 =>
                           dp_n174, Z => dp_N105);
   dp_U183 : OAI22D1 port map( A1 => dp_n197, A2 => dp_n55, B1 => dp_n54, B2 =>
                           dp_n175, Z => dp_N106);
   dp_U182 : OAI22D1 port map( A1 => dp_n196, A2 => dp_n55, B1 => dp_n54, B2 =>
                           dp_n176, Z => dp_N107);
   dp_U181 : OAI22D1 port map( A1 => dp_n195, A2 => dp_n55, B1 => dp_n54, B2 =>
                           dp_n177, Z => dp_N108);
   dp_U180 : OAI22D1 port map( A1 => dp_n194, A2 => dp_n55, B1 => dp_n54, B2 =>
                           dp_n178, Z => dp_N109);
   dp_U179 : OAI22D1 port map( A1 => dp_n193, A2 => dp_n55, B1 => dp_n54, B2 =>
                           dp_n179, Z => dp_N110);
   dp_U178 : OAI22D1 port map( A1 => dp_n192, A2 => dp_n55, B1 => dp_n54, B2 =>
                           dp_n1801, Z => dp_N111);
   dp_U177 : OAI22D1 port map( A1 => dp_n191, A2 => dp_n55, B1 => dp_n54, B2 =>
                           dp_n181, Z => dp_N112);
   dp_U176 : OAI22D1 port map( A1 => dp_n1901, A2 => dp_n55, B1 => dp_n54, B2 
                           => dp_n182, Z => dp_N113);
   dp_U175 : OAI22D1 port map( A1 => dp_n189, A2 => dp_n55, B1 => dp_n54, B2 =>
                           dp_n183, Z => dp_N114);
   dp_U174 : OAI22D1 port map( A1 => dp_n188, A2 => dp_n55, B1 => dp_n54, B2 =>
                           dp_n184, Z => dp_N115);
   dp_U173 : OAI22D1 port map( A1 => dp_n187, A2 => dp_n55, B1 => dp_n54, B2 =>
                           dp_n185, Z => dp_N116);
   dp_U172 : OAI22D1 port map( A1 => add_r_sel, A2 => dp_n170, B1 => dp_n2020, 
                           B2 => dp_n1650, Z => dp_N118);
   dp_U171 : OAI22D1 port map( A1 => add_r_sel, A2 => dp_n171, B1 => dp_n2010, 
                           B2 => dp_n1650, Z => dp_N119);
   dp_U170 : OAI22D1 port map( A1 => add_r_sel, A2 => dp_n172, B1 => dp_n200, 
                           B2 => dp_n1650, Z => dp_N120);
   dp_U169 : OAI22D1 port map( A1 => add_r_sel, A2 => dp_n173, B1 => dp_n199, 
                           B2 => dp_n1650, Z => dp_N121);
   dp_U168 : OAI22D1 port map( A1 => add_r_sel, A2 => dp_n174, B1 => dp_n198, 
                           B2 => dp_n1650, Z => dp_N122);
   dp_U167 : OAI22D1 port map( A1 => add_r_sel, A2 => dp_n175, B1 => dp_n197, 
                           B2 => dp_n1650, Z => dp_N123);
   dp_U166 : OAI22D1 port map( A1 => add_r_sel, A2 => dp_n176, B1 => dp_n196, 
                           B2 => dp_n1650, Z => dp_N124);
   dp_U165 : OAI22D1 port map( A1 => add_r_sel, A2 => dp_n177, B1 => dp_n195, 
                           B2 => dp_n1650, Z => dp_N125);
   dp_U164 : OAI22D1 port map( A1 => add_r_sel, A2 => dp_n178, B1 => dp_n194, 
                           B2 => dp_n1650, Z => dp_N126);
   dp_U163 : OAI22D1 port map( A1 => add_r_sel, A2 => dp_n179, B1 => dp_n193, 
                           B2 => dp_n1650, Z => dp_N127);
   dp_U162 : OAI22D1 port map( A1 => add_r_sel, A2 => dp_n1801, B1 => dp_n192, 
                           B2 => dp_n1650, Z => dp_N128);
   dp_U161 : OAI22D1 port map( A1 => add_r_sel, A2 => dp_n181, B1 => dp_n191, 
                           B2 => dp_n1650, Z => dp_N129);
   dp_U160 : OAI22D1 port map( A1 => add_r_sel, A2 => dp_n182, B1 => dp_n1901, 
                           B2 => dp_n1650, Z => dp_N130);
   dp_U159 : OAI22D1 port map( A1 => add_r_sel, A2 => dp_n183, B1 => dp_n189, 
                           B2 => dp_n1650, Z => dp_N131);
   dp_U158 : OAI22D1 port map( A1 => add_r_sel, A2 => dp_n184, B1 => dp_n188, 
                           B2 => dp_n1650, Z => dp_N132);
   dp_U157 : OAI22D1 port map( A1 => add_r_sel, A2 => dp_n185, B1 => dp_n187, 
                           B2 => dp_n1650, Z => dp_N133);
   dp_U156 : OAI22D1 port map( A1 => dp_n51, A2 => dp_n170, B1 => dp_n2020, B2 
                           => dp_n53, Z => dp_N135);
   dp_U155 : OAI22D1 port map( A1 => dp_n51, A2 => dp_n171, B1 => dp_n2010, B2 
                           => dp_n52, Z => dp_N136);
   dp_U154 : OAI22D1 port map( A1 => dp_n51, A2 => dp_n172, B1 => dp_n200, B2 
                           => dp_n52, Z => dp_N137);
   dp_U153 : OAI22D1 port map( A1 => dp_n51, A2 => dp_n173, B1 => dp_n199, B2 
                           => dp_n53, Z => dp_N138);
   dp_U152 : OAI22D1 port map( A1 => dp_n51, A2 => dp_n174, B1 => dp_n198, B2 
                           => dp_n53, Z => dp_N139);
   dp_U151 : OAI22D1 port map( A1 => dp_n51, A2 => dp_n175, B1 => dp_n197, B2 
                           => dp_n53, Z => dp_N140);
   dp_U150 : OAI22D1 port map( A1 => dp_n51, A2 => dp_n176, B1 => dp_n196, B2 
                           => dp_n53, Z => dp_N141);
   dp_U149 : OAI22D1 port map( A1 => dp_n51, A2 => dp_n177, B1 => dp_n195, B2 
                           => dp_n53, Z => dp_N142);
   dp_U148 : OAI22D1 port map( A1 => dp_n51, A2 => dp_n178, B1 => dp_n194, B2 
                           => dp_n53, Z => dp_N143);
   dp_U147 : OAI22D1 port map( A1 => dp_n51, A2 => dp_n179, B1 => dp_n193, B2 
                           => dp_n53, Z => dp_N144);
   dp_U146 : OAI22D1 port map( A1 => dp_n51, A2 => dp_n1801, B1 => dp_n192, B2 
                           => dp_n53, Z => dp_N145);
   dp_U145 : OAI22D1 port map( A1 => dp_n51, A2 => dp_n181, B1 => dp_n191, B2 
                           => dp_n53, Z => dp_N146);
   dp_U144 : OAI22D1 port map( A1 => dp_n51, A2 => dp_n182, B1 => dp_n1901, B2 
                           => dp_n53, Z => dp_N147);
   dp_U143 : OAI22D1 port map( A1 => dp_n50, A2 => dp_n183, B1 => dp_n189, B2 
                           => dp_n53, Z => dp_N148);
   dp_U142 : OAI22D1 port map( A1 => dp_n50, A2 => dp_n184, B1 => dp_n188, B2 
                           => dp_n53, Z => dp_N149);
   dp_U141 : OAI22D1 port map( A1 => dp_n50, A2 => dp_n185, B1 => dp_n187, B2 
                           => dp_n53, Z => dp_N150);
   dp_U140 : OAI22D1 port map( A1 => dp_n39, A2 => dp_n170, B1 => dp_n2020, B2 
                           => dp_n1640, Z => dp_N152);
   dp_U139 : OAI22D1 port map( A1 => dp_n39, A2 => dp_n171, B1 => dp_n2010, B2 
                           => dp_n1640, Z => dp_N153);
   dp_U138 : OAI22D1 port map( A1 => dp_n39, A2 => dp_n172, B1 => dp_n200, B2 
                           => dp_n1640, Z => dp_N154);
   dp_U137 : OAI22D1 port map( A1 => dp_n39, A2 => dp_n173, B1 => dp_n199, B2 
                           => dp_n1640, Z => dp_N155);
   dp_U136 : OAI22D1 port map( A1 => dp_n39, A2 => dp_n174, B1 => dp_n198, B2 
                           => dp_n1640, Z => dp_N156);
   dp_U135 : OAI22D1 port map( A1 => dp_n39, A2 => dp_n175, B1 => dp_n197, B2 
                           => dp_n1640, Z => dp_N157);
   dp_U134 : OAI22D1 port map( A1 => dp_n39, A2 => dp_n176, B1 => dp_n196, B2 
                           => dp_n1640, Z => dp_N158);
   dp_U133 : OAI22D1 port map( A1 => dp_n39, A2 => dp_n177, B1 => dp_n195, B2 
                           => dp_n1640, Z => dp_N159);
   dp_U132 : OAI22D1 port map( A1 => dp_n39, A2 => dp_n178, B1 => dp_n194, B2 
                           => dp_n1640, Z => dp_N160);
   dp_U131 : OAI22D1 port map( A1 => dp_n39, A2 => dp_n179, B1 => dp_n193, B2 
                           => dp_n1640, Z => dp_N161);
   dp_U130 : OAI22D1 port map( A1 => dp_n39, A2 => dp_n1801, B1 => dp_n192, B2 
                           => dp_n1640, Z => dp_N162);
   dp_U129 : OAI22D1 port map( A1 => dp_n39, A2 => dp_n181, B1 => dp_n191, B2 
                           => dp_n1640, Z => dp_N163);
   dp_U128 : OAI22D1 port map( A1 => dp_n39, A2 => dp_n182, B1 => dp_n1901, B2 
                           => dp_n1640, Z => dp_N164);
   dp_U127 : OAI22D1 port map( A1 => dp_n39, A2 => dp_n183, B1 => dp_n189, B2 
                           => dp_n1640, Z => dp_N165);
   dp_U126 : OAI22D1 port map( A1 => dp_n39, A2 => dp_n184, B1 => dp_n188, B2 
                           => dp_n1640, Z => dp_N166);
   dp_U125 : OAI22D1 port map( A1 => dp_n39, A2 => dp_n185, B1 => dp_n187, B2 
                           => dp_n1640, Z => dp_N167);
   dp_U124 : EXNOR2D1 port map( A1 => dp_cmp_r_0_port, A2 => dp_cmp_l_0_port, Z
                           => dp_n1150);
   dp_U123 : EXNOR2D1 port map( A1 => dp_cmp_r_1_port, A2 => dp_cmp_l_1_port, Z
                           => dp_n1160);
   dp_U122 : EXNOR2D1 port map( A1 => dp_cmp_r_2_port, A2 => dp_cmp_l_2_port, Z
                           => dp_n117);
   dp_U121 : EXNOR2D1 port map( A1 => dp_cmp_r_3_port, A2 => dp_cmp_l_3_port, Z
                           => dp_n1180);
   dp_U120 : EXNOR2D1 port map( A1 => dp_cmp_r_4_port, A2 => dp_cmp_l_4_port, Z
                           => dp_n1110);
   dp_U119 : EXNOR2D1 port map( A1 => dp_cmp_r_5_port, A2 => dp_cmp_l_5_port, Z
                           => dp_n1120);
   dp_U118 : EXNOR2D1 port map( A1 => dp_cmp_r_6_port, A2 => dp_cmp_l_6_port, Z
                           => dp_n1130);
   dp_U117 : EXNOR2D1 port map( A1 => dp_cmp_r_7_port, A2 => dp_cmp_l_7_port, Z
                           => dp_n1140);
   dp_U116 : EXNOR2D1 port map( A1 => dp_cmp_r_8_port, A2 => dp_cmp_l_8_port, Z
                           => dp_n1070);
   dp_U115 : EXNOR2D1 port map( A1 => dp_cmp_r_9_port, A2 => dp_cmp_l_9_port, Z
                           => dp_n1080);
   dp_U114 : EXNOR2D1 port map( A1 => dp_cmp_r_10_port, A2 => dp_cmp_l_10_port,
                           Z => dp_n1090);
   dp_U113 : EXNOR2D1 port map( A1 => dp_cmp_r_11_port, A2 => dp_cmp_l_11_port,
                           Z => dp_n1100);
   dp_U112 : EXNOR2D1 port map( A1 => dp_cmp_r_12_port, A2 => dp_cmp_l_12_port,
                           Z => dp_n1030);
   dp_U111 : EXNOR2D1 port map( A1 => dp_cmp_r_13_port, A2 => dp_cmp_l_13_port,
                           Z => dp_n1040);
   dp_U110 : EXNOR2D1 port map( A1 => dp_cmp_r_14_port, A2 => dp_cmp_l_14_port,
                           Z => dp_n1050);
   dp_U109 : EXNOR2D1 port map( A1 => dp_cmp_r_15_port, A2 => dp_cmp_l_15_port,
                           Z => dp_n1060);
   dp_U108 : EXOR2D1 port map( A1 => sub, A2 => dp_add_r_0_port, Z => 
                           dp_add_r_in_0);
   dp_U107 : EXOR2D1 port map( A1 => sub, A2 => dp_add_r_10_port, Z => 
                           dp_add_r_in_10);
   dp_U106 : EXOR2D1 port map( A1 => sub, A2 => dp_add_r_11_port, Z => 
                           dp_add_r_in_11);
   dp_U105 : EXOR2D1 port map( A1 => sub, A2 => dp_add_r_12_port, Z => 
                           dp_add_r_in_12);
   dp_U104 : EXOR2D1 port map( A1 => sub, A2 => dp_add_r_13_port, Z => 
                           dp_add_r_in_13);
   dp_U103 : EXOR2D1 port map( A1 => sub, A2 => dp_add_r_14_port, Z => 
                           dp_add_r_in_14);
   dp_U102 : EXOR2D1 port map( A1 => sub, A2 => dp_add_r_15_port, Z => 
                           dp_add_r_in_15);
   dp_U101 : EXOR2D1 port map( A1 => sub, A2 => dp_add_r_1_port, Z => 
                           dp_add_r_in_1);
   dp_U100 : EXOR2D1 port map( A1 => sub, A2 => dp_add_r_2_port, Z => 
                           dp_add_r_in_2);
   dp_U99 : EXOR2D1 port map( A1 => sub, A2 => dp_add_r_3_port, Z => 
                           dp_add_r_in_3);
   dp_U98 : EXOR2D1 port map( A1 => sub, A2 => dp_add_r_4_port, Z => 
                           dp_add_r_in_4);
   dp_U97 : EXOR2D1 port map( A1 => sub, A2 => dp_add_r_5_port, Z => 
                           dp_add_r_in_5);
   dp_U96 : EXOR2D1 port map( A1 => sub, A2 => dp_add_r_6_port, Z => 
                           dp_add_r_in_6);
   dp_U95 : EXOR2D1 port map( A1 => sub, A2 => dp_add_r_7_port, Z => 
                           dp_add_r_in_7);
   dp_U94 : EXOR2D1 port map( A1 => sub, A2 => dp_add_r_8_port, Z => 
                           dp_add_r_in_8);
   dp_U93 : EXOR2D1 port map( A1 => sub, A2 => dp_add_r_9_port, Z => 
                           dp_add_r_in_9);
   dp_U92 : NAN3M1D1 port map( A1 => dp_n82, A2 => dp_n80, A3 => dp_n98, Z => 
                           dp_n76);
   dp_U91 : AOI22D1 port map( A1 => data_in(0), A2 => dp_n1630, B1 => 
                           data_out_0_port, B2 => dp_n82, Z => dp_n97);
   dp_U90 : OAI21D1 port map( A1 => dp_n80, A2 => dp_n2020, B => dp_n97, Z => 
                           dp_n75);
   dp_U89 : AOI22D1 port map( A1 => data_in(1), A2 => dp_n1630, B1 => 
                           data_out_1_port, B2 => dp_n82, Z => dp_n96);
   dp_U88 : OAI21D1 port map( A1 => dp_n80, A2 => dp_n2010, B => dp_n96, Z => 
                           dp_n74);
   dp_U87 : AOI22D1 port map( A1 => data_in(2), A2 => dp_n1630, B1 => 
                           data_out_2_port, B2 => dp_n82, Z => dp_n95);
   dp_U86 : OAI21D1 port map( A1 => dp_n80, A2 => dp_n200, B => dp_n95, Z => 
                           dp_n73);
   dp_U85 : AOI22D1 port map( A1 => data_in(3), A2 => dp_n1630, B1 => 
                           data_out_3_port, B2 => dp_n82, Z => dp_n94);
   dp_U84 : OAI21D1 port map( A1 => dp_n80, A2 => dp_n199, B => dp_n94, Z => 
                           dp_n72);
   dp_U83 : AOI22D1 port map( A1 => data_in(4), A2 => dp_n1630, B1 => 
                           data_out_4_port, B2 => dp_n82, Z => dp_n93);
   dp_U82 : OAI21D1 port map( A1 => dp_n80, A2 => dp_n198, B => dp_n93, Z => 
                           dp_n71);
   dp_U81 : AOI22D1 port map( A1 => data_in(5), A2 => dp_n1630, B1 => 
                           data_out_5_port, B2 => dp_n82, Z => dp_n92);
   dp_U80 : OAI21D1 port map( A1 => dp_n80, A2 => dp_n197, B => dp_n92, Z => 
                           dp_n70);
   dp_U79 : AOI22D1 port map( A1 => data_in(6), A2 => dp_n1630, B1 => 
                           data_out_6_port, B2 => dp_n82, Z => dp_n91);
   dp_U78 : OAI21D1 port map( A1 => dp_n80, A2 => dp_n196, B => dp_n91, Z => 
                           dp_n69);
   dp_U77 : AOI22D1 port map( A1 => data_in(7), A2 => dp_n1630, B1 => 
                           data_out_7_port, B2 => dp_n82, Z => dp_n90);
   dp_U76 : OAI21D1 port map( A1 => dp_n80, A2 => dp_n195, B => dp_n90, Z => 
                           dp_n68);
   dp_U75 : AOI22D1 port map( A1 => data_in(8), A2 => dp_n1630, B1 => 
                           data_out_8_port, B2 => dp_n82, Z => dp_n89);
   dp_U74 : OAI21D1 port map( A1 => dp_n80, A2 => dp_n194, B => dp_n89, Z => 
                           dp_n67);
   dp_U73 : AOI22D1 port map( A1 => data_in(9), A2 => dp_n1630, B1 => 
                           data_out_9_port, B2 => dp_n82, Z => dp_n88);
   dp_U72 : OAI21D1 port map( A1 => dp_n80, A2 => dp_n193, B => dp_n88, Z => 
                           dp_n66);
   dp_U71 : AOI22D1 port map( A1 => data_in(10), A2 => dp_n1630, B1 => 
                           data_out_10_port, B2 => dp_n82, Z => dp_n87);
   dp_U70 : OAI21D1 port map( A1 => dp_n80, A2 => dp_n192, B => dp_n87, Z => 
                           dp_n65);
   dp_U69 : AOI22D1 port map( A1 => data_in(11), A2 => dp_n1630, B1 => 
                           data_out_11_port, B2 => dp_n82, Z => dp_n86);
   dp_U68 : OAI21D1 port map( A1 => dp_n80, A2 => dp_n191, B => dp_n86, Z => 
                           dp_n64);
   dp_U67 : AOI22D1 port map( A1 => data_in(12), A2 => dp_n1630, B1 => 
                           data_out_12_port, B2 => dp_n82, Z => dp_n85);
   dp_U66 : OAI21D1 port map( A1 => dp_n80, A2 => dp_n1901, B => dp_n85, Z => 
                           dp_n63);
   dp_U65 : AOI22D1 port map( A1 => data_in(13), A2 => dp_n1630, B1 => 
                           data_out_13_port, B2 => dp_n82, Z => dp_n84);
   dp_U64 : OAI21D1 port map( A1 => dp_n80, A2 => dp_n189, B => dp_n84, Z => 
                           dp_n62);
   dp_U63 : AOI22D1 port map( A1 => data_in(14), A2 => dp_n1630, B1 => 
                           data_out_14_port, B2 => dp_n82, Z => dp_n83);
   dp_U62 : OAI21D1 port map( A1 => dp_n80, A2 => dp_n188, B => dp_n83, Z => 
                           dp_n61);
   dp_U61 : AOI22D1 port map( A1 => data_in(15), A2 => dp_n1630, B1 => 
                           data_out_15_port, B2 => dp_n82, Z => dp_n81);
   dp_U60 : OAI21D1 port map( A1 => dp_n80, A2 => dp_n187, B => dp_n81, Z => 
                           dp_n60);
   dp_add_1_root_add_129_2_U1_15 : EXOR3D1 port map( A1 => dp_add_l_15_port, A2
                           => dp_add_r_in_15, A3 => 
                           dp_add_1_root_add_129_2_carry_15_port, Z => 
                           dp_add_out_15_port);
   dp_add_1_root_add_129_2_U1_0 : ADFULD1 port map( A => dp_add_l_0_port, B => 
                           dp_add_r_in_0, CI => sub, CO => 
                           dp_add_1_root_add_129_2_carry_1_port, S => 
                           dp_add_out_0_port);
   dp_add_1_root_add_129_2_U1_1 : ADFULD1 port map( A => dp_add_l_1_port, B => 
                           dp_add_r_in_1, CI => 
                           dp_add_1_root_add_129_2_carry_1_port, CO => 
                           dp_add_1_root_add_129_2_carry_2_port, S => 
                           dp_add_out_1_port);
   dp_add_1_root_add_129_2_U1_2 : ADFULD1 port map( A => dp_add_l_2_port, B => 
                           dp_add_r_in_2, CI => 
                           dp_add_1_root_add_129_2_carry_2_port, CO => 
                           dp_add_1_root_add_129_2_carry_3_port, S => 
                           dp_add_out_2_port);
   dp_add_1_root_add_129_2_U1_3 : ADFULD1 port map( A => dp_add_l_3_port, B => 
                           dp_add_r_in_3, CI => 
                           dp_add_1_root_add_129_2_carry_3_port, CO => 
                           dp_add_1_root_add_129_2_carry_4_port, S => 
                           dp_add_out_3_port);
   dp_add_1_root_add_129_2_U1_4 : ADFULD1 port map( A => dp_add_l_4_port, B => 
                           dp_add_r_in_4, CI => 
                           dp_add_1_root_add_129_2_carry_4_port, CO => 
                           dp_add_1_root_add_129_2_carry_5_port, S => 
                           dp_add_out_4_port);
   dp_add_1_root_add_129_2_U1_5 : ADFULD1 port map( A => dp_add_l_5_port, B => 
                           dp_add_r_in_5, CI => 
                           dp_add_1_root_add_129_2_carry_5_port, CO => 
                           dp_add_1_root_add_129_2_carry_6_port, S => 
                           dp_add_out_5_port);
   dp_add_1_root_add_129_2_U1_6 : ADFULD1 port map( A => dp_add_l_6_port, B => 
                           dp_add_r_in_6, CI => 
                           dp_add_1_root_add_129_2_carry_6_port, CO => 
                           dp_add_1_root_add_129_2_carry_7_port, S => 
                           dp_add_out_6_port);
   dp_add_1_root_add_129_2_U1_7 : ADFULD1 port map( A => dp_add_l_7_port, B => 
                           dp_add_r_in_7, CI => 
                           dp_add_1_root_add_129_2_carry_7_port, CO => 
                           dp_add_1_root_add_129_2_carry_8_port, S => 
                           dp_add_out_7_port);
   dp_add_1_root_add_129_2_U1_8 : ADFULD1 port map( A => dp_add_l_8_port, B => 
                           dp_add_r_in_8, CI => 
                           dp_add_1_root_add_129_2_carry_8_port, CO => 
                           dp_add_1_root_add_129_2_carry_9_port, S => 
                           dp_add_out_8_port);
   dp_add_1_root_add_129_2_U1_9 : ADFULD1 port map( A => dp_add_l_9_port, B => 
                           dp_add_r_in_9, CI => 
                           dp_add_1_root_add_129_2_carry_9_port, CO => 
                           dp_add_1_root_add_129_2_carry_10_port, S => 
                           dp_add_out_9_port);
   dp_add_1_root_add_129_2_U1_10 : ADFULD1 port map( A => dp_add_l_10_port, B 
                           => dp_add_r_in_10, CI => 
                           dp_add_1_root_add_129_2_carry_10_port, CO => 
                           dp_add_1_root_add_129_2_carry_11_port, S => 
                           dp_add_out_10_port);
   dp_add_1_root_add_129_2_U1_11 : ADFULD1 port map( A => dp_add_l_11_port, B 
                           => dp_add_r_in_11, CI => 
                           dp_add_1_root_add_129_2_carry_11_port, CO => 
                           dp_add_1_root_add_129_2_carry_12_port, S => 
                           dp_add_out_11_port);
   dp_add_1_root_add_129_2_U1_12 : ADFULD1 port map( A => dp_add_l_12_port, B 
                           => dp_add_r_in_12, CI => 
                           dp_add_1_root_add_129_2_carry_12_port, CO => 
                           dp_add_1_root_add_129_2_carry_13_port, S => 
                           dp_add_out_12_port);
   dp_add_1_root_add_129_2_U1_13 : ADFULD1 port map( A => dp_add_l_13_port, B 
                           => dp_add_r_in_13, CI => 
                           dp_add_1_root_add_129_2_carry_13_port, CO => 
                           dp_add_1_root_add_129_2_carry_14_port, S => 
                           dp_add_out_13_port);
   dp_add_1_root_add_129_2_U1_14 : ADFULD1 port map( A => dp_add_l_14_port, B 
                           => dp_add_r_in_14, CI => 
                           dp_add_1_root_add_129_2_carry_14_port, CO => 
                           dp_add_1_root_add_129_2_carry_15_port, S => 
                           dp_add_out_14_port);
   cn_U49 : TIEHI port map( Z => cn_sub);
   cn_U48 : TIELO port map( Z => cn_wr_addr_1);
   cn_U47 : INVD1 port map( A => reset, Z => cn_n32);
   cn_U46 : NOR3D1 port map( A1 => cn_n15, A2 => cn_current_state_3_port, A3 =>
                           cn_current_state_1_port, Z => wr_sel_en_1_port);
   cn_U38 : NOR2D1 port map( A1 => cn_current_state_2_port, A2 => 
                           cn_current_state_3_port, Z => cn_n24);
   cn_U37 : INVD1 port map( A => cn_current_state_0_port, Z => cn_n9);
   cn_U36 : NAN4D1 port map( A1 => cn_current_state_3_port, A2 => cn_n9, A3 => 
                           cn_n14, A4 => cn_n31, Z => cn_n23);
   cn_U35 : INVD1 port map( A => cn_current_state_3_port, Z => cn_n12);
   cn_U34 : NAN4D1 port map( A1 => cn_current_state_0_port, A2 => 
                           cn_current_state_2_port, A3 => cn_n14, A4 => cn_n12,
                           Z => cn_n27);
   cn_U33 : NAN3D1 port map( A1 => cn_n27, A2 => cn_n23, A3 => cn_n28, Z => 
                           cn_next_state_0_port);
   cn_U32 : INVD1 port map( A => cn_current_state_2_port, Z => cn_n31);
   cn_U31 : NOR2D1 port map( A1 => cn_n31, A2 => cn_current_state_0_port, Z => 
                           cn_n15);
   cn_U30 : INVD1 port map( A => cn_current_state_1_port, Z => cn_n14);
   cn_U29 : INVD1 port map( A => cn_n24, Z => cn_n13);
   cn_U28 : NAN3D1 port map( A1 => cn_current_state_0_port, A2 => cn_n24, A3 =>
                           cn_current_state_1_port, Z => cn_n22);
   cn_U27 : AND2D1 port map( A1 => cn_N21, A2 => cn_next_state_2_port, Z => 
                           cn_n30);
   cn_U26 : NOR2D1 port map( A1 => cn_n6, A2 => cn_next_state_1_port, Z => 
                           cn_N21);
   cn_U25 : INVD1 port map( A => cn_next_state_0_port, Z => cn_n6);
   cn_U24 : NOR2D1 port map( A1 => cn_n7, A2 => cn_next_state_2_port, Z => 
                           cn_n16);
   cn_U23 : NOR3D1 port map( A1 => cn_n8, A2 => cn_next_state_0_port, A3 => 
                           cn_n7, Z => cn_cmp_l_sel);
   cn_U22 : INVD1 port map( A => cn_cmp_l_sel, Z => cn_n2);
   cn_U21 : INVD1 port map( A => cn_n2, Z => add_l_sel);
   cn_U20 : INVD1 port map( A => cn_next_state_1_port, Z => cn_n7);
   cn_U19 : NOR2D1 port map( A1 => cn_n31, A2 => cn_n14, Z => cn_n29);
   cn_U18 : INVD1 port map( A => cn_next_state_2_port, Z => cn_n8);
   cn_U17 : NOR3D1 port map( A1 => cn_next_state_0_port, A2 => 
                           cn_next_state_1_port, A3 => cn_n8, Z => 
                           rd_addr_0_port);
   cn_U16 : NOR2D1 port map( A1 => cmp_r_sel, A2 => rd_addr_0_port, Z => cn_n18
                           );
   cn_U15 : INVD1 port map( A => cn_n19, Z => cmp_l_en);
   cn_U14 : NAN2D1 port map( A1 => cn_n19, A2 => cn_n17, Z => add_l_en);
   cn_U13 : AO211D1 port map( A1 => cn_n8, A2 => cn_N21, B => add_l_sel, C => 
                           wr_addr_0, Z => wr_sel_en_0_port);
   cn_U12 : OAI21M20D1 port map( A1 => cn_n6, A2 => cn_n16, B => cn_n3, Z => 
                           wr_addr_0);
   cn_U11 : NOR3D1 port map( A1 => cn_n7, A2 => cn_n8, A3 => cn_n6, Z => 
                           cmp_r_sel);
   cn_U10 : INVD1 port map( A => cn_n210, Z => cn_n11);
   cn_U9 : NOR2D1 port map( A1 => greater, A2 => equal, Z => cn_n20);
   cn_U8 : INVD1 port map( A => cn_n18, Z => cmp_r_en);
   cn_U7 : NAN2D1 port map( A1 => cn_n18, A2 => cn_n17, Z => add_r_en);
   cn_U6 : INVD1 port map( A => cmp_r_sel, Z => cn_n3);
   cn_U5 : NAN2D1 port map( A1 => cn_n20, A2 => cn_n11, Z => cn_n17);
   cn_U4 : NAN2D1 port map( A1 => cn_n3, A2 => cn_n17, Z => add_r_sel);
   cn_U3 : INVD1 port map( A => cn_n17, Z => rd_addr_1_port);
   cn_ready_reg : DFFRPQ1 port map( D => cn_n30, CK => clk, RB => cn_n32, Q => 
                           ready);
   cn_req_reg : DFFSPQ1 port map( D => cn_N21, CK => clk, SB => cn_n32, Q => 
                           req);
   cn_current_state_reg_1 : DFFRPQ1 port map( D => cn_next_state_1_port, CK => 
                           clk, RB => cn_n32, Q => cn_current_state_1_port);
   cn_current_state_reg_2 : DFFRPQ1 port map( D => cn_next_state_2_port, CK => 
                           clk, RB => cn_n32, Q => cn_current_state_2_port);
   cn_current_state_reg_0 : DFFRPQ1 port map( D => cn_next_state_0_port, CK => 
                           clk, RB => cn_n32, Q => cn_current_state_0_port);
   cn_current_state_reg_3 : DFFRPQ1 port map( D => rd_addr_1_port, CK => clk, 
                           RB => cn_n32, Q => cn_current_state_3_port);
   cn_U45 : OAI21D1 port map( A1 => cn_n15, A2 => cn_n29, B => cn_n12, Z => 
                           cn_n210);
   cn_U44 : AOI22D1 port map( A1 => cn_n24, A2 => cn_n9, B1 => equal, B2 => 
                           cn_n11, Z => cn_n28);
   cn_U43 : EXNOR2D1 port map( A1 => cn_current_state_0_port, A2 => 
                           cn_current_state_1_port, Z => cn_n25);
   cn_U42 : NAN3M1D1 port map( A1 => equal, A2 => cn_n11, A3 => greater, Z => 
                           cn_n26);
   cn_U41 : OAI211D1 port map( A1 => cn_n25, A2 => cn_n13, B => cn_n26, C => 
                           cn_n23, Z => cn_next_state_1_port);
   cn_U40 : OAI211D1 port map( A1 => cn_n20, A2 => cn_n210, B => cn_n22, C => 
                           cn_n23, Z => cn_next_state_2_port);
   cn_U39 : AOI211D1 port map( A1 => cn_next_state_0_port, A2 => cn_n16, B => 
                           cmp_r_sel, C => add_l_sel, Z => cn_n19);

end flat_dpctrl_gcd_16_10;
