
library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

package CONV_PACK_gp_custom is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_gp_custom;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_gp_custom.all;

architecture flat_filter_none_20 of gp_custom is

   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component MUXB2DL
      port( A0, A1, SL : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN4D1
      port( A1, A2, A3, A4 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AO22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AO31D1
      port( A1, A2, A3, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22M10D1
      port( B1, B2, A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3M1D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211D1
      port( A1, A2, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFBD2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFRPQ1
      port( D, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component DFERPQ1
      port( D, CEB, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFSPQ1
      port( D, CK, SB : in std_logic;  Q : out std_logic);
   end component;
   
   component OA21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI32D1
      port( A1, A2, A3, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   signal N62, N63, N64, avs_readdata_31_port, avs_readdata_30_port, 
      avs_readdata_29_port, avs_readdata_28_port, avs_readdata_27_port, 
      avs_readdata_26_port, avs_readdata_25_port, avs_readdata_24_port, 
      avs_readdata_23_port, avs_readdata_22_port, avs_readdata_21_port, 
      avs_readdata_20_port, avs_readdata_19_port, avs_readdata_18_port, 
      avs_readdata_17_port, avs_readdata_16_port, avs_readdata_15_port, 
      avs_readdata_14_port, avs_readdata_13_port, avs_readdata_12_port, 
      avs_readdata_11_port, avs_readdata_10_port, avs_readdata_9_port, 
      avs_readdata_8_port, avs_readdata_7_port, avs_readdata_6_port, 
      avs_readdata_5_port, avs_readdata_4_port, avs_readdata_3_port, 
      avs_readdata_2_port, avs_readdata_1_port, avs_readdata_0_port, 
      stop_sim_port, out_buf_255_port, out_buf_254_port, out_buf_253_port, 
      out_buf_252_port, out_buf_251_port, out_buf_250_port, out_buf_249_port, 
      out_buf_248_port, out_buf_247_port, out_buf_246_port, out_buf_245_port, 
      out_buf_244_port, out_buf_243_port, out_buf_242_port, out_buf_241_port, 
      out_buf_240_port, out_buf_239_port, out_buf_238_port, out_buf_237_port, 
      out_buf_236_port, out_buf_235_port, out_buf_234_port, out_buf_233_port, 
      out_buf_232_port, out_buf_231_port, out_buf_230_port, out_buf_229_port, 
      out_buf_228_port, out_buf_227_port, out_buf_226_port, out_buf_225_port, 
      out_buf_224_port, out_buf_223_port, out_buf_222_port, out_buf_221_port, 
      out_buf_220_port, out_buf_219_port, out_buf_218_port, out_buf_217_port, 
      out_buf_216_port, out_buf_215_port, out_buf_214_port, out_buf_213_port, 
      out_buf_212_port, out_buf_211_port, out_buf_210_port, out_buf_209_port, 
      out_buf_208_port, out_buf_207_port, out_buf_206_port, out_buf_205_port, 
      out_buf_204_port, out_buf_203_port, out_buf_202_port, out_buf_201_port, 
      out_buf_200_port, out_buf_199_port, out_buf_198_port, out_buf_197_port, 
      out_buf_196_port, out_buf_195_port, out_buf_194_port, out_buf_193_port, 
      out_buf_192_port, out_buf_191_port, out_buf_190_port, out_buf_189_port, 
      out_buf_188_port, out_buf_187_port, out_buf_186_port, out_buf_185_port, 
      out_buf_184_port, out_buf_183_port, out_buf_182_port, out_buf_181_port, 
      out_buf_180_port, out_buf_179_port, out_buf_178_port, out_buf_177_port, 
      out_buf_176_port, out_buf_175_port, out_buf_174_port, out_buf_173_port, 
      out_buf_172_port, out_buf_171_port, out_buf_170_port, out_buf_169_port, 
      out_buf_168_port, out_buf_167_port, out_buf_166_port, out_buf_165_port, 
      out_buf_164_port, out_buf_163_port, out_buf_162_port, out_buf_161_port, 
      out_buf_160_port, out_buf_159_port, out_buf_158_port, out_buf_157_port, 
      out_buf_156_port, out_buf_155_port, out_buf_154_port, out_buf_153_port, 
      out_buf_152_port, out_buf_151_port, out_buf_150_port, out_buf_149_port, 
      out_buf_148_port, out_buf_147_port, out_buf_146_port, out_buf_145_port, 
      out_buf_144_port, out_buf_143_port, out_buf_142_port, out_buf_141_port, 
      out_buf_140_port, out_buf_139_port, out_buf_138_port, out_buf_137_port, 
      out_buf_136_port, out_buf_135_port, out_buf_134_port, out_buf_133_port, 
      out_buf_132_port, out_buf_131_port, out_buf_130_port, out_buf_129_port, 
      out_buf_128_port, out_buf_127_port, out_buf_126_port, out_buf_125_port, 
      out_buf_124_port, out_buf_123_port, out_buf_122_port, out_buf_121_port, 
      out_buf_120_port, out_buf_119_port, out_buf_118_port, out_buf_117_port, 
      out_buf_116_port, out_buf_115_port, out_buf_114_port, out_buf_113_port, 
      out_buf_112_port, out_buf_111_port, out_buf_110_port, out_buf_109_port, 
      out_buf_108_port, out_buf_107_port, out_buf_106_port, out_buf_105_port, 
      out_buf_104_port, out_buf_103_port, out_buf_102_port, out_buf_101_port, 
      out_buf_100_port, out_buf_99_port, out_buf_98_port, out_buf_97_port, 
      out_buf_96_port, out_buf_95_port, out_buf_94_port, out_buf_93_port, 
      out_buf_92_port, out_buf_91_port, out_buf_90_port, out_buf_89_port, 
      out_buf_88_port, out_buf_87_port, out_buf_86_port, out_buf_85_port, 
      out_buf_84_port, out_buf_83_port, out_buf_82_port, out_buf_81_port, 
      out_buf_80_port, out_buf_79_port, out_buf_78_port, out_buf_77_port, 
      out_buf_76_port, out_buf_75_port, out_buf_74_port, out_buf_73_port, 
      out_buf_72_port, out_buf_71_port, out_buf_70_port, out_buf_69_port, 
      out_buf_68_port, out_buf_67_port, out_buf_66_port, out_buf_65_port, 
      out_buf_64_port, out_buf_63_port, out_buf_62_port, out_buf_61_port, 
      out_buf_60_port, out_buf_59_port, out_buf_58_port, out_buf_57_port, 
      out_buf_56_port, out_buf_55_port, out_buf_54_port, out_buf_53_port, 
      out_buf_52_port, out_buf_51_port, out_buf_50_port, out_buf_49_port, 
      out_buf_48_port, out_buf_47_port, out_buf_46_port, out_buf_45_port, 
      out_buf_44_port, out_buf_43_port, out_buf_42_port, out_buf_41_port, 
      out_buf_40_port, out_buf_39_port, out_buf_38_port, out_buf_37_port, 
      out_buf_36_port, out_buf_35_port, out_buf_34_port, out_buf_33_port, 
      out_buf_32_port, out_buf_31_port, out_buf_30_port, out_buf_29_port, 
      out_buf_28_port, out_buf_27_port, out_buf_26_port, out_buf_25_port, 
      out_buf_24_port, out_buf_23_port, out_buf_22_port, out_buf_21_port, 
      out_buf_20_port, out_buf_19_port, out_buf_18_port, out_buf_17_port, 
      out_buf_16_port, out_buf_15_port, out_buf_14_port, out_buf_13_port, 
      out_buf_12_port, out_buf_11_port, out_buf_10_port, out_buf_9_port, 
      out_buf_8_port, out_buf_7_port, out_buf_6_port, out_buf_5_port, 
      out_buf_4_port, out_buf_3_port, out_buf_2_port, out_buf_1_port, 
      out_buf_0_port, coeff_memory_0_31, coeff_memory_0_30, coeff_memory_0_29, 
      coeff_memory_0_28, coeff_memory_0_27, coeff_memory_0_26, 
      coeff_memory_0_25, coeff_memory_0_24, coeff_memory_0_23, 
      coeff_memory_0_22, coeff_memory_0_21, coeff_memory_0_20, 
      coeff_memory_0_19, coeff_memory_0_18, coeff_memory_0_17, 
      coeff_memory_0_16, coeff_memory_0_15, coeff_memory_0_14, 
      coeff_memory_0_13, coeff_memory_0_12, coeff_memory_0_11, 
      coeff_memory_0_10, coeff_memory_0_9, coeff_memory_0_8, coeff_memory_0_7, 
      coeff_memory_0_6, coeff_memory_0_5, coeff_memory_0_4, coeff_memory_0_3, 
      coeff_memory_0_2, coeff_memory_0_1, coeff_memory_0_0, coeff_memory_1_31, 
      coeff_memory_1_30, coeff_memory_1_29, coeff_memory_1_28, 
      coeff_memory_1_27, coeff_memory_1_26, coeff_memory_1_25, 
      coeff_memory_1_24, coeff_memory_1_23, coeff_memory_1_22, 
      coeff_memory_1_21, coeff_memory_1_20, coeff_memory_1_19, 
      coeff_memory_1_18, coeff_memory_1_17, coeff_memory_1_16, 
      coeff_memory_1_15, coeff_memory_1_14, coeff_memory_1_13, 
      coeff_memory_1_12, coeff_memory_1_11, coeff_memory_1_10, coeff_memory_1_9
      , coeff_memory_1_8, coeff_memory_1_7, coeff_memory_1_6, coeff_memory_1_5,
      coeff_memory_1_4, coeff_memory_1_3, coeff_memory_1_2, coeff_memory_1_1, 
      coeff_memory_1_0, coeff_memory_2_31, coeff_memory_2_30, coeff_memory_2_29
      , coeff_memory_2_28, coeff_memory_2_27, coeff_memory_2_26, 
      coeff_memory_2_25, coeff_memory_2_24, coeff_memory_2_23, 
      coeff_memory_2_22, coeff_memory_2_21, coeff_memory_2_20, 
      coeff_memory_2_19, coeff_memory_2_18, coeff_memory_2_17, 
      coeff_memory_2_16, coeff_memory_2_15, coeff_memory_2_14, 
      coeff_memory_2_13, coeff_memory_2_12, coeff_memory_2_11, 
      coeff_memory_2_10, coeff_memory_2_9, coeff_memory_2_8, coeff_memory_2_7, 
      coeff_memory_2_6, coeff_memory_2_5, coeff_memory_2_4, coeff_memory_2_3, 
      coeff_memory_2_2, coeff_memory_2_1, coeff_memory_2_0, coeff_memory_3_31, 
      coeff_memory_3_30, coeff_memory_3_29, coeff_memory_3_28, 
      coeff_memory_3_27, coeff_memory_3_26, coeff_memory_3_25, 
      coeff_memory_3_24, coeff_memory_3_23, coeff_memory_3_22, 
      coeff_memory_3_21, coeff_memory_3_20, coeff_memory_3_19, 
      coeff_memory_3_18, coeff_memory_3_17, coeff_memory_3_16, 
      coeff_memory_3_15, coeff_memory_3_14, coeff_memory_3_13, 
      coeff_memory_3_12, coeff_memory_3_11, coeff_memory_3_10, coeff_memory_3_9
      , coeff_memory_3_8, coeff_memory_3_7, coeff_memory_3_6, coeff_memory_3_5,
      coeff_memory_3_4, coeff_memory_3_3, coeff_memory_3_2, coeff_memory_3_1, 
      coeff_memory_3_0, coeff_memory_4_31, coeff_memory_4_30, coeff_memory_4_29
      , coeff_memory_4_28, coeff_memory_4_27, coeff_memory_4_26, 
      coeff_memory_4_25, coeff_memory_4_24, coeff_memory_4_23, 
      coeff_memory_4_22, coeff_memory_4_21, coeff_memory_4_20, 
      coeff_memory_4_19, coeff_memory_4_18, coeff_memory_4_17, 
      coeff_memory_4_16, coeff_memory_4_15, coeff_memory_4_14, 
      coeff_memory_4_13, coeff_memory_4_12, coeff_memory_4_11, 
      coeff_memory_4_10, coeff_memory_4_9, coeff_memory_4_8, coeff_memory_4_7, 
      coeff_memory_4_6, coeff_memory_4_5, coeff_memory_4_4, coeff_memory_4_3, 
      coeff_memory_4_2, coeff_memory_4_1, coeff_memory_4_0, 
      operand_regs_255_port, operand_regs_254_port, operand_regs_253_port, 
      operand_regs_252_port, operand_regs_251_port, operand_regs_250_port, 
      operand_regs_249_port, operand_regs_248_port, operand_regs_247_port, 
      operand_regs_246_port, operand_regs_245_port, operand_regs_244_port, 
      operand_regs_243_port, operand_regs_242_port, operand_regs_241_port, 
      operand_regs_240_port, operand_regs_239_port, operand_regs_238_port, 
      operand_regs_237_port, operand_regs_236_port, operand_regs_235_port, 
      operand_regs_234_port, operand_regs_233_port, operand_regs_232_port, 
      operand_regs_231_port, operand_regs_230_port, operand_regs_229_port, 
      operand_regs_228_port, operand_regs_227_port, operand_regs_226_port, 
      operand_regs_225_port, operand_regs_224_port, operand_regs_223_port, 
      operand_regs_222_port, operand_regs_221_port, operand_regs_220_port, 
      operand_regs_219_port, operand_regs_218_port, operand_regs_217_port, 
      operand_regs_216_port, operand_regs_215_port, operand_regs_214_port, 
      operand_regs_213_port, operand_regs_212_port, operand_regs_211_port, 
      operand_regs_210_port, operand_regs_209_port, operand_regs_208_port, 
      operand_regs_207_port, operand_regs_206_port, operand_regs_205_port, 
      operand_regs_204_port, operand_regs_203_port, operand_regs_202_port, 
      operand_regs_201_port, operand_regs_200_port, operand_regs_199_port, 
      operand_regs_198_port, operand_regs_197_port, operand_regs_196_port, 
      operand_regs_195_port, operand_regs_194_port, operand_regs_193_port, 
      operand_regs_192_port, operand_regs_191_port, operand_regs_190_port, 
      operand_regs_189_port, operand_regs_188_port, operand_regs_187_port, 
      operand_regs_186_port, operand_regs_185_port, operand_regs_184_port, 
      operand_regs_183_port, operand_regs_182_port, operand_regs_181_port, 
      operand_regs_180_port, operand_regs_179_port, operand_regs_178_port, 
      operand_regs_177_port, operand_regs_176_port, operand_regs_175_port, 
      operand_regs_174_port, operand_regs_173_port, operand_regs_172_port, 
      operand_regs_171_port, operand_regs_170_port, operand_regs_169_port, 
      operand_regs_168_port, operand_regs_167_port, operand_regs_166_port, 
      operand_regs_165_port, operand_regs_164_port, operand_regs_163_port, 
      operand_regs_162_port, operand_regs_161_port, operand_regs_160_port, 
      operand_regs_159_port, operand_regs_158_port, operand_regs_157_port, 
      operand_regs_156_port, operand_regs_155_port, operand_regs_154_port, 
      operand_regs_153_port, operand_regs_152_port, operand_regs_151_port, 
      operand_regs_150_port, operand_regs_149_port, operand_regs_148_port, 
      operand_regs_147_port, operand_regs_146_port, operand_regs_145_port, 
      operand_regs_144_port, operand_regs_143_port, operand_regs_142_port, 
      operand_regs_141_port, operand_regs_140_port, operand_regs_139_port, 
      operand_regs_138_port, operand_regs_137_port, operand_regs_136_port, 
      operand_regs_135_port, operand_regs_134_port, operand_regs_133_port, 
      operand_regs_132_port, operand_regs_131_port, operand_regs_130_port, 
      operand_regs_129_port, operand_regs_128_port, operand_regs_127_port, 
      operand_regs_126_port, operand_regs_125_port, operand_regs_124_port, 
      operand_regs_123_port, operand_regs_122_port, operand_regs_121_port, 
      operand_regs_120_port, operand_regs_119_port, operand_regs_118_port, 
      operand_regs_117_port, operand_regs_116_port, operand_regs_115_port, 
      operand_regs_114_port, operand_regs_113_port, operand_regs_112_port, 
      operand_regs_111_port, operand_regs_110_port, operand_regs_109_port, 
      operand_regs_108_port, operand_regs_107_port, operand_regs_106_port, 
      operand_regs_105_port, operand_regs_104_port, operand_regs_103_port, 
      operand_regs_102_port, operand_regs_101_port, operand_regs_100_port, 
      operand_regs_99_port, operand_regs_98_port, operand_regs_97_port, 
      operand_regs_96_port, operand_regs_95_port, operand_regs_94_port, 
      operand_regs_93_port, operand_regs_92_port, operand_regs_91_port, 
      operand_regs_90_port, operand_regs_89_port, operand_regs_88_port, 
      operand_regs_87_port, operand_regs_86_port, operand_regs_85_port, 
      operand_regs_84_port, operand_regs_83_port, operand_regs_82_port, 
      operand_regs_81_port, operand_regs_80_port, operand_regs_79_port, 
      operand_regs_78_port, operand_regs_77_port, operand_regs_76_port, 
      operand_regs_75_port, operand_regs_74_port, operand_regs_73_port, 
      operand_regs_72_port, operand_regs_71_port, operand_regs_70_port, 
      operand_regs_69_port, operand_regs_68_port, operand_regs_67_port, 
      operand_regs_66_port, operand_regs_65_port, operand_regs_64_port, 
      operand_regs_63_port, operand_regs_62_port, operand_regs_61_port, 
      operand_regs_60_port, operand_regs_59_port, operand_regs_58_port, 
      operand_regs_57_port, operand_regs_56_port, operand_regs_55_port, 
      operand_regs_54_port, operand_regs_53_port, operand_regs_52_port, 
      operand_regs_51_port, operand_regs_50_port, operand_regs_49_port, 
      operand_regs_48_port, operand_regs_47_port, operand_regs_46_port, 
      operand_regs_45_port, operand_regs_44_port, operand_regs_43_port, 
      operand_regs_42_port, operand_regs_41_port, operand_regs_40_port, 
      operand_regs_39_port, operand_regs_38_port, operand_regs_37_port, 
      operand_regs_36_port, operand_regs_35_port, operand_regs_34_port, 
      operand_regs_33_port, operand_regs_32_port, operand_regs_31_port, 
      operand_regs_30_port, operand_regs_29_port, operand_regs_28_port, 
      operand_regs_27_port, operand_regs_26_port, operand_regs_25_port, 
      operand_regs_24_port, operand_regs_23_port, operand_regs_22_port, 
      operand_regs_21_port, operand_regs_20_port, operand_regs_19_port, 
      operand_regs_18_port, operand_regs_17_port, operand_regs_16_port, 
      operand_regs_15_port, operand_regs_14_port, operand_regs_13_port, 
      operand_regs_12_port, operand_regs_11_port, operand_regs_10_port, 
      operand_regs_9_port, operand_regs_8_port, operand_regs_7_port, 
      operand_regs_6_port, operand_regs_5_port, operand_regs_4_port, 
      operand_regs_3_port, operand_regs_2_port, operand_regs_1_port, 
      operand_regs_0_port, in_trigger, out_trigger, coeff_load, operand_load, 
      read_comp_res, filt_mult_inputs, N66, comp_res_159_port, 
      comp_res_158_port, comp_res_157_port, comp_res_156_port, 
      comp_res_155_port, comp_res_154_port, comp_res_153_port, 
      comp_res_152_port, comp_res_151_port, comp_res_150_port, 
      comp_res_149_port, comp_res_148_port, comp_res_147_port, 
      comp_res_146_port, comp_res_145_port, comp_res_144_port, 
      comp_res_143_port, comp_res_142_port, comp_res_141_port, 
      comp_res_140_port, comp_res_139_port, comp_res_138_port, 
      comp_res_137_port, comp_res_136_port, comp_res_135_port, 
      comp_res_134_port, comp_res_133_port, comp_res_132_port, 
      comp_res_131_port, comp_res_130_port, comp_res_129_port, 
      comp_res_128_port, comp_res_127_port, comp_res_126_port, 
      comp_res_125_port, comp_res_124_port, comp_res_123_port, 
      comp_res_122_port, comp_res_121_port, comp_res_120_port, 
      comp_res_119_port, comp_res_118_port, comp_res_117_port, 
      comp_res_116_port, comp_res_115_port, comp_res_114_port, 
      comp_res_113_port, comp_res_112_port, comp_res_111_port, 
      comp_res_110_port, comp_res_109_port, comp_res_108_port, 
      comp_res_107_port, comp_res_106_port, comp_res_105_port, 
      comp_res_104_port, comp_res_103_port, comp_res_102_port, 
      comp_res_101_port, comp_res_100_port, comp_res_99_port, comp_res_98_port,
      comp_res_97_port, comp_res_96_port, comp_res_95_port, comp_res_94_port, 
      comp_res_93_port, comp_res_92_port, comp_res_91_port, comp_res_90_port, 
      comp_res_89_port, comp_res_88_port, comp_res_87_port, comp_res_86_port, 
      comp_res_85_port, comp_res_84_port, comp_res_83_port, comp_res_82_port, 
      comp_res_81_port, comp_res_80_port, comp_res_79_port, comp_res_78_port, 
      comp_res_77_port, comp_res_76_port, comp_res_75_port, comp_res_74_port, 
      comp_res_73_port, comp_res_72_port, comp_res_71_port, comp_res_70_port, 
      comp_res_69_port, comp_res_68_port, comp_res_67_port, comp_res_66_port, 
      comp_res_65_port, comp_res_64_port, comp_res_63_port, comp_res_62_port, 
      comp_res_61_port, comp_res_60_port, comp_res_59_port, comp_res_58_port, 
      comp_res_57_port, comp_res_56_port, comp_res_55_port, comp_res_54_port, 
      comp_res_53_port, comp_res_52_port, comp_res_51_port, comp_res_50_port, 
      comp_res_49_port, comp_res_48_port, comp_res_47_port, comp_res_46_port, 
      comp_res_45_port, comp_res_44_port, comp_res_43_port, comp_res_42_port, 
      comp_res_41_port, comp_res_40_port, comp_res_39_port, comp_res_38_port, 
      comp_res_37_port, comp_res_36_port, comp_res_35_port, comp_res_34_port, 
      comp_res_33_port, comp_res_32_port, comp_res_31_port, comp_res_30_port, 
      comp_res_29_port, comp_res_28_port, comp_res_27_port, comp_res_26_port, 
      comp_res_25_port, comp_res_24_port, comp_res_23_port, comp_res_22_port, 
      comp_res_21_port, comp_res_20_port, comp_res_19_port, comp_res_18_port, 
      comp_res_17_port, comp_res_16_port, comp_res_15_port, comp_res_14_port, 
      comp_res_13_port, comp_res_12_port, comp_res_11_port, comp_res_10_port, 
      comp_res_9_port, comp_res_8_port, comp_res_7_port, comp_res_6_port, 
      comp_res_5_port, comp_res_4_port, comp_res_3_port, comp_res_2_port, 
      comp_res_1_port, comp_res_0_port, N1978, N1979, N1980, N1981, N1982, 
      N1983, N1984, N1985, N1986, N1987, N1988, N1989, N1990, N1991, N1992, 
      N1993, N1994, N1995, N1996, N1997, N1998, N1999, N2000, N2001, N2002, 
      N2003, N2004, N2005, N2006, N2007, N2008, N2009, in_buf_255_port, 
      in_buf_254_port, in_buf_253_port, in_buf_252_port, in_buf_251_port, 
      in_buf_250_port, in_buf_249_port, in_buf_248_port, in_buf_247_port, 
      in_buf_246_port, in_buf_245_port, in_buf_244_port, in_buf_243_port, 
      in_buf_242_port, in_buf_241_port, in_buf_240_port, in_buf_239_port, 
      in_buf_238_port, in_buf_237_port, in_buf_236_port, in_buf_235_port, 
      in_buf_234_port, in_buf_233_port, in_buf_232_port, in_buf_231_port, 
      in_buf_230_port, in_buf_229_port, in_buf_228_port, in_buf_227_port, 
      in_buf_226_port, in_buf_225_port, in_buf_224_port, in_buf_223_port, 
      in_buf_222_port, in_buf_221_port, in_buf_220_port, in_buf_219_port, 
      in_buf_218_port, in_buf_217_port, in_buf_216_port, in_buf_215_port, 
      in_buf_214_port, in_buf_213_port, in_buf_212_port, in_buf_211_port, 
      in_buf_210_port, in_buf_209_port, in_buf_208_port, in_buf_207_port, 
      in_buf_206_port, in_buf_205_port, in_buf_204_port, in_buf_203_port, 
      in_buf_202_port, in_buf_201_port, in_buf_200_port, in_buf_199_port, 
      in_buf_198_port, in_buf_197_port, in_buf_196_port, in_buf_195_port, 
      in_buf_194_port, in_buf_193_port, in_buf_192_port, in_buf_191_port, 
      in_buf_190_port, in_buf_189_port, in_buf_188_port, in_buf_187_port, 
      in_buf_186_port, in_buf_185_port, in_buf_184_port, in_buf_183_port, 
      in_buf_182_port, in_buf_181_port, in_buf_180_port, in_buf_179_port, 
      in_buf_178_port, in_buf_177_port, in_buf_176_port, in_buf_175_port, 
      in_buf_174_port, in_buf_173_port, in_buf_172_port, in_buf_171_port, 
      in_buf_170_port, in_buf_169_port, in_buf_168_port, in_buf_167_port, 
      in_buf_166_port, in_buf_165_port, in_buf_164_port, in_buf_163_port, 
      in_buf_162_port, in_buf_161_port, in_buf_160_port, in_buf_159_port, 
      in_buf_158_port, in_buf_157_port, in_buf_156_port, in_buf_155_port, 
      in_buf_154_port, in_buf_153_port, in_buf_152_port, in_buf_151_port, 
      in_buf_150_port, in_buf_149_port, in_buf_148_port, in_buf_147_port, 
      in_buf_146_port, in_buf_145_port, in_buf_144_port, in_buf_143_port, 
      in_buf_142_port, in_buf_141_port, in_buf_140_port, in_buf_139_port, 
      in_buf_138_port, in_buf_137_port, in_buf_136_port, in_buf_135_port, 
      in_buf_134_port, in_buf_133_port, in_buf_132_port, in_buf_131_port, 
      in_buf_130_port, in_buf_129_port, in_buf_128_port, in_buf_127_port, 
      in_buf_126_port, in_buf_125_port, in_buf_124_port, in_buf_123_port, 
      in_buf_122_port, in_buf_121_port, in_buf_120_port, in_buf_119_port, 
      in_buf_118_port, in_buf_117_port, in_buf_116_port, in_buf_115_port, 
      in_buf_114_port, in_buf_113_port, in_buf_112_port, in_buf_111_port, 
      in_buf_110_port, in_buf_109_port, in_buf_108_port, in_buf_107_port, 
      in_buf_106_port, in_buf_105_port, in_buf_104_port, in_buf_103_port, 
      in_buf_102_port, in_buf_101_port, in_buf_100_port, in_buf_99_port, 
      in_buf_98_port, in_buf_97_port, in_buf_96_port, in_buf_95_port, 
      in_buf_94_port, in_buf_93_port, in_buf_92_port, in_buf_91_port, 
      in_buf_90_port, in_buf_89_port, in_buf_88_port, in_buf_87_port, 
      in_buf_86_port, in_buf_85_port, in_buf_84_port, in_buf_83_port, 
      in_buf_82_port, in_buf_81_port, in_buf_80_port, in_buf_79_port, 
      in_buf_78_port, in_buf_77_port, in_buf_76_port, in_buf_75_port, 
      in_buf_74_port, in_buf_73_port, in_buf_72_port, in_buf_71_port, 
      in_buf_70_port, in_buf_69_port, in_buf_68_port, in_buf_67_port, 
      in_buf_66_port, in_buf_65_port, in_buf_64_port, in_buf_63_port, 
      in_buf_62_port, in_buf_61_port, in_buf_60_port, in_buf_59_port, 
      in_buf_58_port, in_buf_57_port, in_buf_56_port, in_buf_55_port, 
      in_buf_54_port, in_buf_53_port, in_buf_52_port, in_buf_51_port, 
      in_buf_50_port, in_buf_49_port, in_buf_48_port, in_buf_47_port, 
      in_buf_46_port, in_buf_45_port, in_buf_44_port, in_buf_43_port, 
      in_buf_42_port, in_buf_41_port, in_buf_40_port, in_buf_39_port, 
      in_buf_38_port, in_buf_37_port, in_buf_36_port, in_buf_35_port, 
      in_buf_34_port, in_buf_33_port, in_buf_32_port, in_buf_31_port, 
      in_buf_30_port, in_buf_29_port, in_buf_28_port, in_buf_27_port, 
      in_buf_26_port, in_buf_25_port, in_buf_24_port, in_buf_23_port, 
      in_buf_22_port, in_buf_21_port, in_buf_20_port, in_buf_19_port, 
      in_buf_18_port, in_buf_17_port, in_buf_16_port, in_buf_15_port, 
      in_buf_14_port, in_buf_13_port, in_buf_12_port, in_buf_11_port, 
      in_buf_10_port, in_buf_9_port, in_buf_8_port, in_buf_7_port, 
      in_buf_6_port, in_buf_5_port, in_buf_4_port, in_buf_3_port, in_buf_2_port
      , in_buf_1_port, in_buf_0_port, N2010, N2011, N2012, N2013, N2014, N2015,
      N2016, N2017, N2018, N2019, N2020, N2021, N2022, N2023, N2024, N2025, 
      N2026, N2027, N2028, N2029, N2030, N2031, N2032, N2033, N2034, N2035, 
      N2036, N2037, N2038, N2039, N2040, N2041, in_busy, out_busy, 
      in_counter_2_port, in_counter_1_port, in_counter_0_port, odd, odd1, N2850
      , N2851, N2852, N2853, N2854, N2855, N2856, N2857, N2858, N2859, N2860, 
      N2861, N2862, N2863, N2864, N2865, N2867, N2868, N2869, N2870, N2871, 
      N2872, N2873, N2874, N2875, N2876, N2877, N2878, N2879, N2880, N2881, 
      N2882, N2888, N2889, N2890, N2891, N2892, N2893, N2894, N2895, N2896, 
      N2897, N2898, N2899, N2900, N2901, N2902, N2903, N2913, N2914, N2915, 
      N2916, N2917, N2918, N2919, N2920, N2921, N2922, N2923, N2924, N2925, 
      N2926, N2927, N2928, N2929, N2930, N2931, N2932, N2933, N2934, N2935, 
      N2936, N2937, N2938, N2939, N2940, N2941, N2942, N2943, N2944, N2945, 
      N2946, N2947, N2948, N2949, N2950, N2951, N2952, N2953, N2954, N2955, 
      N2956, N2957, N2958, N2959, N2960, N2961, N2962, N2963, N2964, N2965, 
      N2966, N2967, N2968, N2969, N2970, N2971, N2972, N2973, N2974, N2975, 
      N2976, N2977, N2978, N2979, N2980, N2981, N2982, N2983, N2984, N2985, 
      N2986, N2987, N2988, N2989, N2990, N2991, N2992, N2993, N2994, N2995, 
      N2996, N2997, N2998, N2999, N3000, N3001, N3002, N3003, N3004, N3005, 
      N3006, N3007, N3008, N3009, N3010, N3011, N3012, N3013, N3014, N3015, 
      N3016, N3017, N3018, N3019, N3020, N3021, N3022, N3023, N3024, N3025, 
      N3026, N3027, N3028, N3029, N3030, N3031, N3032, N3033, N3034, N3035, 
      N3036, N3037, N3038, N3039, N3040, N3041, N3042, N3043, N3044, N3045, 
      N3046, N3047, N3048, N3049, N3050, N3051, N3052, N3053, N3054, N3055, 
      N3056, N3057, N3058, N3059, N3060, N3061, N3062, N3063, N3064, N3065, 
      N3066, N3067, N3068, N3069, N3070, N3071, N3072, N3073, N3074, N3075, 
      N3076, N3077, N3078, N3079, N3080, N3081, N3082, N3083, N3084, N3085, 
      N3086, N3087, N3088, N3089, N3090, N3091, N3092, N3093, N3094, N3095, 
      N3096, N3097, N3098, N3099, N3100, N3101, N3102, N3103, N3104, N3105, 
      N3106, N3107, N3108, N3109, N3110, N3111, N3112, N3113, N3114, N3115, 
      N3116, N3117, N3118, N3119, N3120, N3121, N3122, N3123, N3124, N3125, 
      N3126, N3127, N3128, N3129, N3130, N3131, N3132, N3133, N3134, N3135, 
      N3136, N3137, N3138, N3139, N3140, N3141, N3142, N3143, N3144, N3145, 
      N3146, N3147, N3148, N3149, N3150, N3151, N3152, N3153, N3154, N3155, 
      N3156, N3157, N3158, N3159, N3160, N3161, N3162, N3163, N3164, N3165, 
      N3166, N3167, N3168, N3201, N3202, N3203, N3204, N3205, N3206, N3207, 
      N3208, N3209, N3210, N3211, N3212, N3213, N3214, N3215, N3216, N3217, 
      N3218, N3219, N3220, N3221, N3222, N3223, N3224, N3225, N3226, N3227, 
      N3228, N3229, N3230, N3231, N3232, N3233, N3234, N3235, N3236, N3237, 
      N3238, N3239, N3240, N3241, N3242, N3243, N3244, N3245, N3246, N3247, 
      N3248, N3249, N3250, N3251, N3252, N3253, N3254, N3255, N3256, N3257, 
      N3258, N3259, N3260, N3261, N3262, N3263, N3264, N3265, N3266, N3267, 
      N3268, N3269, N3270, N3271, N3272, N3273, N3274, N3275, N3276, N3277, 
      N3278, N3279, N3280, N3281, N3282, N3283, N3284, N3285, N3286, N3287, 
      N3288, N3289, N3290, N3291, N3292, N3293, N3294, N3295, N3296, N3297, 
      N3298, N3299, N3300, N3301, N3302, N3303, N3304, N3305, N3306, N3307, 
      N3308, N3309, N3310, N3311, N3312, N3313, N3314, N3315, N3316, N3317, 
      N3318, N3319, N3320, N3321, N3322, N3323, N3324, N3325, N3326, N3327, 
      N3328, N3329, N3330, N3331, N3332, N3333, N3334, N3335, N3336, N3337, 
      N3338, N3339, N3340, N3341, N3342, N3343, N3344, N3345, N3346, N3347, 
      N3348, N3349, N3350, N3351, N3352, N3353, N3354, N3355, N3356, N3357, 
      N3358, N3359, N3360, N3361, N3362, N3363, N3364, N3365, N3366, N3367, 
      N3368, N3369, N3370, N3371, N3372, N3373, N3374, N3375, N3376, N3377, 
      N3378, N3379, N3380, N3381, N3382, N3383, N3384, N3385, N3386, N3387, 
      N3388, N3389, N3390, N3391, N3392, n4, n5, n10, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n5900, 
      n6000, n6100, n6300, n6400, n65, n68, n69, n70, n72, n73, n74, n76, n77, 
      n78, n79, n81, n84, n85, n86, n87, n88, n89, n91, n92, n93, n95, n96, n97
      , n99, n100, n101, n103, n104, n106, n107, n108, n109, n110, n111, n114, 
      n115, n118, n119, n120, n122, n123, n124, n125, n126, n127, n128, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n201, 
      n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, 
      n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, 
      n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, 
      n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, 
      n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, 
      n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, 
      n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, 
      n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, 
      n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, 
      n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, 
      n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, 
      n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, 
      n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, 
      n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, 
      n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, 
      n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, 
      n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, 
      n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, 
      n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, 
      n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, 
      n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, 
      n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, 
      n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, 
      n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, 
      n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, 
      n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, 
      n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, 
      n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, 
      n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, 
      n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, 
      n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, 
      n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, 
      n586, n587, n588, n589, n5901, n591, n592, n593, n594, n595, n596, n597, 
      n598, n599, n6001, n601, n602, n603, n604, n605, n606, n607, n608, n609, 
      n6101, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, 
      n622, n623, n624, n625, n626, n627, n628, n629, n6301, n631, n632, n633, 
      n634, n635, n636, n637, n638, n639, n6401, n641, n642, n643, n644, n645, 
      n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, 
      n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, 
      n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, 
      n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, 
      n694, n695, n696, n697, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, 
      n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, 
      n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, 
      n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, 
      n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, 
      n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, 
      n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, 
      n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, 
      n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, 
      n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, 
      n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, 
      n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, 
      n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, 
      n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, 
      n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, 
      n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, 
      n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, 
      n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, 
      n_1319, mult_21_C241_n1451, mult_21_C241_n1450, mult_21_C241_n1449, 
      mult_21_C241_n1448, mult_21_C241_n1447, mult_21_C241_n1446, 
      mult_21_C241_n1445, mult_21_C241_n1444, mult_21_C241_n1443, 
      mult_21_C241_n1442, mult_21_C241_n1441, mult_21_C241_n1440, 
      mult_21_C241_n1439, mult_21_C241_n1438, mult_21_C241_n1437, 
      mult_21_C241_n1436, mult_21_C241_n1435, mult_21_C241_n1434, 
      mult_21_C241_n1433, mult_21_C241_n1432, mult_21_C241_n1431, 
      mult_21_C241_n1430, mult_21_C241_n1429, mult_21_C241_n1428, 
      mult_21_C241_n1427, mult_21_C241_n1426, mult_21_C241_n1425, 
      mult_21_C241_n1424, mult_21_C241_n1423, mult_21_C241_n1422, 
      mult_21_C241_n1421, mult_21_C241_n1420, mult_21_C241_n1419, 
      mult_21_C241_n1418, mult_21_C241_n1417, mult_21_C241_n1416, 
      mult_21_C241_n1415, mult_21_C241_n1414, mult_21_C241_n1413, 
      mult_21_C241_n1412, mult_21_C241_n1411, mult_21_C241_n1410, 
      mult_21_C241_n1409, mult_21_C241_n1408, mult_21_C241_n1407, 
      mult_21_C241_n1406, mult_21_C241_n1405, mult_21_C241_n1404, 
      mult_21_C241_n1403, mult_21_C241_n1402, mult_21_C241_n1401, 
      mult_21_C241_n1400, mult_21_C241_n1399, mult_21_C241_n1398, 
      mult_21_C241_n1397, mult_21_C241_n1396, mult_21_C241_n1395, 
      mult_21_C241_n1394, mult_21_C241_n1393, mult_21_C241_n1392, 
      mult_21_C241_n1391, mult_21_C241_n1390, mult_21_C241_n1389, 
      mult_21_C241_n1388, mult_21_C241_n1387, mult_21_C241_n1386, 
      mult_21_C241_n1385, mult_21_C241_n1384, mult_21_C241_n1383, 
      mult_21_C241_n1382, mult_21_C241_n1381, mult_21_C241_n1380, 
      mult_21_C241_n1379, mult_21_C241_n1378, mult_21_C241_n1377, 
      mult_21_C241_n1376, mult_21_C241_n1375, mult_21_C241_n1226, 
      mult_21_C241_n1225, mult_21_C241_n1224, mult_21_C241_n1223, 
      mult_21_C241_n1222, mult_21_C241_n1221, mult_21_C241_n1220, 
      mult_21_C241_n1219, mult_21_C241_n1218, mult_21_C241_n1217, 
      mult_21_C241_n1216, mult_21_C241_n1215, mult_21_C241_n1214, 
      mult_21_C241_n1213, mult_21_C241_n1212, mult_21_C241_n1211, 
      mult_21_C241_n1210, mult_21_C241_n1209, mult_21_C241_n1208, 
      mult_21_C241_n1207, mult_21_C241_n1206, mult_21_C241_n1205, 
      mult_21_C241_n1204, mult_21_C241_n1203, mult_21_C241_n1202, 
      mult_21_C241_n1201, mult_21_C241_n1200, mult_21_C241_n1199, 
      mult_21_C241_n1198, mult_21_C241_n1197, mult_21_C241_n1196, 
      mult_21_C241_n1195, mult_21_C241_n1194, mult_21_C241_n1193, 
      mult_21_C241_n1192, mult_21_C241_n1191, mult_21_C241_n1190, 
      mult_21_C241_n1189, mult_21_C241_n1188, mult_21_C241_n1187, 
      mult_21_C241_n1186, mult_21_C241_n1185, mult_21_C241_n1184, 
      mult_21_C241_n1183, mult_21_C241_n1182, mult_21_C241_n1181, 
      mult_21_C241_n1180, mult_21_C241_n1179, mult_21_C241_n1178, 
      mult_21_C241_n1177, mult_21_C241_n1176, mult_21_C241_n1175, 
      mult_21_C241_n1174, mult_21_C241_n1173, mult_21_C241_n1172, 
      mult_21_C241_n1171, mult_21_C241_n1170, mult_21_C241_n1169, 
      mult_21_C241_n1168, mult_21_C241_n1167, mult_21_C241_n1166, 
      mult_21_C241_n1165, mult_21_C241_n1164, mult_21_C241_n1163, 
      mult_21_C241_n1162, mult_21_C241_n1161, mult_21_C241_n1160, 
      mult_21_C241_n1159, mult_21_C241_n1158, mult_21_C241_n1157, 
      mult_21_C241_n1156, mult_21_C241_n1155, mult_21_C241_n1154, 
      mult_21_C241_n1153, mult_21_C241_n1152, mult_21_C241_n1151, 
      mult_21_C241_n1150, mult_21_C241_n1149, mult_21_C241_n1148, 
      mult_21_C241_n1147, mult_21_C241_n1146, mult_21_C241_n1145, 
      mult_21_C241_n1144, mult_21_C241_n1143, mult_21_C241_n1142, 
      mult_21_C241_n1141, mult_21_C241_n1140, mult_21_C241_n1139, 
      mult_21_C241_n1138, mult_21_C241_n1137, mult_21_C241_n1136, 
      mult_21_C241_n1135, mult_21_C241_n1134, mult_21_C241_n1133, 
      mult_21_C241_n1132, mult_21_C241_n1131, mult_21_C241_n1130, 
      mult_21_C241_n1129, mult_21_C241_n1128, mult_21_C241_n1127, 
      mult_21_C241_n1126, mult_21_C241_n1125, mult_21_C241_n1124, 
      mult_21_C241_n1123, mult_21_C241_n1122, mult_21_C241_n1121, 
      mult_21_C241_n1120, mult_21_C241_n1119, mult_21_C241_n1118, 
      mult_21_C241_n1117, mult_21_C241_n1116, mult_21_C241_n1115, 
      mult_21_C241_n1114, mult_21_C241_n1113, mult_21_C241_n1112, 
      mult_21_C241_n1111, mult_21_C241_n1110, mult_21_C241_n1109, 
      mult_21_C241_n1108, mult_21_C241_n1107, mult_21_C241_n1106, 
      mult_21_C241_n1105, mult_21_C241_n1104, mult_21_C241_n1103, 
      mult_21_C241_n1102, mult_21_C241_n1101, mult_21_C241_n1100, 
      mult_21_C241_n1099, mult_21_C241_n1098, mult_21_C241_n1097, 
      mult_21_C241_n1096, mult_21_C241_n1095, mult_21_C241_n1094, 
      mult_21_C241_n1093, mult_21_C241_n1092, mult_21_C241_n1091, 
      mult_21_C241_n1090, mult_21_C241_n1089, mult_21_C241_n1088, 
      mult_21_C241_n1087, mult_21_C241_n1086, mult_21_C241_n1085, 
      mult_21_C241_n1084, mult_21_C241_n1083, mult_21_C241_n1082, 
      mult_21_C241_n1081, mult_21_C241_n1080, mult_21_C241_n1079, 
      mult_21_C241_n1078, mult_21_C241_n1077, mult_21_C241_n1076, 
      mult_21_C241_n1075, mult_21_C241_n1074, mult_21_C241_n1073, 
      mult_21_C241_n1072, mult_21_C241_n1071, mult_21_C241_n1070, 
      mult_21_C241_n1069, mult_21_C241_n1068, mult_21_C241_n1067, 
      mult_21_C241_n1066, mult_21_C241_n1065, mult_21_C241_n1064, 
      mult_21_C241_n1063, mult_21_C241_n1062, mult_21_C241_n1061, 
      mult_21_C241_n1060, mult_21_C241_n1059, mult_21_C241_n1058, 
      mult_21_C241_n1057, mult_21_C241_n1056, mult_21_C241_n1055, 
      mult_21_C241_n1054, mult_21_C241_n1053, mult_21_C241_n1052, 
      mult_21_C241_n1051, mult_21_C241_n1050, mult_21_C241_n1049, 
      mult_21_C241_n1048, mult_21_C241_n1047, mult_21_C241_n1046, 
      mult_21_C241_n1045, mult_21_C241_n1044, mult_21_C241_n1043, 
      mult_21_C241_n1042, mult_21_C241_n1041, mult_21_C241_n1040, 
      mult_21_C241_n1039, mult_21_C241_n1038, mult_21_C241_n1037, 
      mult_21_C241_n1036, mult_21_C241_n1035, mult_21_C241_n1034, 
      mult_21_C241_n1033, mult_21_C241_n1032, mult_21_C241_n1031, 
      mult_21_C241_n1030, mult_21_C241_n1029, mult_21_C241_n1028, 
      mult_21_C241_n1027, mult_21_C241_n1026, mult_21_C241_n1025, 
      mult_21_C241_n1024, mult_21_C241_n1023, mult_21_C241_n1022, 
      mult_21_C241_n1021, mult_21_C241_n1020, mult_21_C241_n1019, 
      mult_21_C241_n1018, mult_21_C241_n1017, mult_21_C241_n1016, 
      mult_21_C241_n1015, mult_21_C241_n1014, mult_21_C241_n1013, 
      mult_21_C241_n1012, mult_21_C241_n1011, mult_21_C241_n1010, 
      mult_21_C241_n1009, mult_21_C241_n1008, mult_21_C241_n1007, 
      mult_21_C241_n1006, mult_21_C241_n1005, mult_21_C241_n1004, 
      mult_21_C241_n1003, mult_21_C241_n1002, mult_21_C241_n1001, 
      mult_21_C241_n1000, mult_21_C241_n999, mult_21_C241_n998, 
      mult_21_C241_n997, mult_21_C241_n996, mult_21_C241_n995, 
      mult_21_C241_n994, mult_21_C241_n993, mult_21_C241_n992, 
      mult_21_C241_n991, mult_21_C241_n990, mult_21_C241_n989, 
      mult_21_C241_n988, mult_21_C241_n987, mult_21_C241_n986, 
      mult_21_C241_n985, mult_21_C241_n984, mult_21_C241_n983, 
      mult_21_C241_n982, mult_21_C241_n981, mult_21_C241_n980, 
      mult_21_C241_n979, mult_21_C241_n978, mult_21_C241_n977, 
      mult_21_C241_n976, mult_21_C241_n975, mult_21_C241_n974, 
      mult_21_C241_n973, mult_21_C241_n972, mult_21_C241_n971, 
      mult_21_C241_n970, mult_21_C241_n969, mult_21_C241_n968, 
      mult_21_C241_n967, mult_21_C241_n966, mult_21_C241_n965, 
      mult_21_C241_n964, mult_21_C241_n963, mult_21_C241_n962, 
      mult_21_C241_n961, mult_21_C241_n960, mult_21_C241_n959, 
      mult_21_C241_n958, mult_21_C241_n957, mult_21_C241_n956, 
      mult_21_C241_n955, mult_21_C241_n953, mult_21_C241_n952, 
      mult_21_C241_n951, mult_21_C241_n950, mult_21_C241_n949, 
      mult_21_C241_n948, mult_21_C241_n947, mult_21_C241_n946, 
      mult_21_C241_n945, mult_21_C241_n944, mult_21_C241_n943, 
      mult_21_C241_n942, mult_21_C241_n941, mult_21_C241_n940, 
      mult_21_C241_n939, mult_21_C241_n923, mult_21_C241_n922, 
      mult_21_C241_n921, mult_21_C241_n920, mult_21_C241_n919, 
      mult_21_C241_n918, mult_21_C241_n917, mult_21_C241_n916, 
      mult_21_C241_n915, mult_21_C241_n914, mult_21_C241_n913, 
      mult_21_C241_n912, mult_21_C241_n911, mult_21_C241_n910, 
      mult_21_C241_n909, mult_21_C241_n908, mult_21_C241_n907, 
      mult_21_C241_n906, mult_21_C241_n905, mult_21_C241_n904, 
      mult_21_C241_n903, mult_21_C241_n902, mult_21_C241_n901, 
      mult_21_C241_n900, mult_21_C241_n899, mult_21_C241_n898, 
      mult_21_C241_n897, mult_21_C241_n896, mult_21_C241_n895, 
      mult_21_C241_n894, mult_21_C241_n893, mult_21_C241_n892, 
      mult_21_C241_n891, mult_21_C241_n890, mult_21_C241_n889, 
      mult_21_C241_n888, mult_21_C241_n887, mult_21_C241_n886, 
      mult_21_C241_n885, mult_21_C241_n884, mult_21_C241_n883, 
      mult_21_C241_n882, mult_21_C241_n881, mult_21_C241_n880, 
      mult_21_C241_n879, mult_21_C241_n878, mult_21_C241_n877, 
      mult_21_C241_n876, mult_21_C241_n875, mult_21_C241_n874, 
      mult_21_C241_n873, mult_21_C241_n872, mult_21_C241_n871, 
      mult_21_C241_n870, mult_21_C241_n869, mult_21_C241_n868, 
      mult_21_C241_n867, mult_21_C241_n866, mult_21_C241_n865, 
      mult_21_C241_n864, mult_21_C241_n863, mult_21_C241_n862, 
      mult_21_C241_n861, mult_21_C241_n860, mult_21_C241_n859, 
      mult_21_C241_n858, mult_21_C241_n857, mult_21_C241_n856, 
      mult_21_C241_n855, mult_21_C241_n854, mult_21_C241_n853, 
      mult_21_C241_n852, mult_21_C241_n851, mult_21_C241_n850, 
      mult_21_C241_n849, mult_21_C241_n848, mult_21_C241_n847, 
      mult_21_C241_n846, mult_21_C241_n845, mult_21_C241_n844, 
      mult_21_C241_n843, mult_21_C241_n842, mult_21_C241_n841, 
      mult_21_C241_n840, mult_21_C241_n839, mult_21_C241_n838, 
      mult_21_C241_n837, mult_21_C241_n836, mult_21_C241_n835, 
      mult_21_C241_n834, mult_21_C241_n833, mult_21_C241_n832, 
      mult_21_C241_n831, mult_21_C241_n830, mult_21_C241_n829, 
      mult_21_C241_n828, mult_21_C241_n827, mult_21_C241_n826, 
      mult_21_C241_n825, mult_21_C241_n824, mult_21_C241_n823, 
      mult_21_C241_n822, mult_21_C241_n821, mult_21_C241_n820, 
      mult_21_C241_n819, mult_21_C241_n818, mult_21_C241_n817, 
      mult_21_C241_n816, mult_21_C241_n815, mult_21_C241_n814, 
      mult_21_C241_n813, mult_21_C241_n812, mult_21_C241_n811, 
      mult_21_C241_n810, mult_21_C241_n809, mult_21_C241_n808, 
      mult_21_C241_n807, mult_21_C241_n806, mult_21_C241_n805, 
      mult_21_C241_n804, mult_21_C241_n803, mult_21_C241_n802, 
      mult_21_C241_n801, mult_21_C241_n800, mult_21_C241_n799, 
      mult_21_C241_n798, mult_21_C241_n797, mult_21_C241_n796, 
      mult_21_C241_n795, mult_21_C241_n794, mult_21_C241_n793, 
      mult_21_C241_n792, mult_21_C241_n791, mult_21_C241_n790, 
      mult_21_C241_n789, mult_21_C241_n788, mult_21_C241_n787, 
      mult_21_C241_n786, mult_21_C241_n785, mult_21_C241_n784, 
      mult_21_C241_n783, mult_21_C241_n782, mult_21_C241_n781, 
      mult_21_C241_n780, mult_21_C241_n779, mult_21_C241_n778, 
      mult_21_C241_n777, mult_21_C241_n776, mult_21_C241_n775, 
      mult_21_C241_n774, mult_21_C241_n773, mult_21_C241_n772, 
      mult_21_C241_n771, mult_21_C241_n770, mult_21_C241_n769, 
      mult_21_C241_n768, mult_21_C241_n767, mult_21_C241_n766, 
      mult_21_C241_n765, mult_21_C241_n764, mult_21_C241_n763, 
      mult_21_C241_n762, mult_21_C241_n761, mult_21_C241_n760, 
      mult_21_C241_n759, mult_21_C241_n758, mult_21_C241_n757, 
      mult_21_C241_n756, mult_21_C241_n755, mult_21_C241_n754, 
      mult_21_C241_n753, mult_21_C241_n752, mult_21_C241_n751, 
      mult_21_C241_n750, mult_21_C241_n749, mult_21_C241_n748, 
      mult_21_C241_n747, mult_21_C241_n746, mult_21_C241_n745, 
      mult_21_C241_n744, mult_21_C241_n743, mult_21_C241_n742, 
      mult_21_C241_n741, mult_21_C241_n740, mult_21_C241_n739, 
      mult_21_C241_n738, mult_21_C241_n737, mult_21_C241_n736, 
      mult_21_C241_n735, mult_21_C241_n734, mult_21_C241_n733, 
      mult_21_C241_n732, mult_21_C241_n731, mult_21_C241_n730, 
      mult_21_C241_n729, mult_21_C241_n728, mult_21_C241_n727, 
      mult_21_C241_n726, mult_21_C241_n725, mult_21_C241_n724, 
      mult_21_C241_n723, mult_21_C241_n722, mult_21_C241_n721, 
      mult_21_C241_n720, mult_21_C241_n719, mult_21_C241_n718, 
      mult_21_C241_n717, mult_21_C241_n716, mult_21_C241_n715, 
      mult_21_C241_n714, mult_21_C241_n713, mult_21_C241_n712, 
      mult_21_C241_n711, mult_21_C241_n710, mult_21_C241_n709, 
      mult_21_C241_n708, mult_21_C241_n707, mult_21_C241_n706, 
      mult_21_C241_n705, mult_21_C241_n704, mult_21_C241_n703, 
      mult_21_C241_n702, mult_21_C241_n701, mult_21_C241_n700, 
      mult_21_C241_n699, mult_21_C241_n698, mult_21_C241_n697, 
      mult_21_C241_n696, mult_21_C241_n695, mult_21_C241_n694, 
      mult_21_C241_n693, mult_21_C241_n692, mult_21_C241_n691, 
      mult_21_C241_n690, mult_21_C241_n689, mult_21_C241_n688, 
      mult_21_C241_n687, mult_21_C241_n686, mult_21_C241_n685, 
      mult_21_C241_n684, mult_21_C241_n683, mult_21_C241_n682, 
      mult_21_C241_n681, mult_21_C241_n680, mult_21_C241_n679, 
      mult_21_C241_n678, mult_21_C241_n677, mult_21_C241_n676, 
      mult_21_C241_n675, mult_21_C241_n674, mult_21_C241_n673, 
      mult_21_C241_n672, mult_21_C241_n671, mult_21_C241_n670, 
      mult_21_C241_n669, mult_21_C241_n668, mult_21_C241_n667, 
      mult_21_C241_n666, mult_21_C241_n665, mult_21_C241_n664, 
      mult_21_C241_n663, mult_21_C241_n662, mult_21_C241_n661, 
      mult_21_C241_n660, mult_21_C241_n659, mult_21_C241_n658, 
      mult_21_C241_n657, mult_21_C241_n656, mult_21_C241_n655, 
      mult_21_C241_n654, mult_21_C241_n653, mult_21_C241_n652, 
      mult_21_C241_n651, mult_21_C241_n650, mult_21_C241_n649, 
      mult_21_C241_n648, mult_21_C241_n647, mult_21_C241_n646, 
      mult_21_C241_n645, mult_21_C241_n644, mult_21_C241_n643, 
      mult_21_C241_n642, mult_21_C241_n641, mult_21_C241_n640, 
      mult_21_C241_n639, mult_21_C241_n638, mult_21_C241_n637, 
      mult_21_C241_n636, mult_21_C241_n635, mult_21_C241_n634, 
      mult_21_C241_n633, mult_21_C241_n632, mult_21_C241_n631, 
      mult_21_C241_n630, mult_21_C241_n629, mult_21_C241_n628, 
      mult_21_C241_n627, mult_21_C241_n626, mult_21_C241_n625, 
      mult_21_C241_n624, mult_21_C241_n623, mult_21_C241_n622, 
      mult_21_C241_n621, mult_21_C241_n620, mult_21_C241_n619, 
      mult_21_C241_n618, mult_21_C241_n617, mult_21_C241_n616, 
      mult_21_C241_n615, mult_21_C241_n614, mult_21_C241_n613, 
      mult_21_C241_n612, mult_21_C241_n611, mult_21_C241_n610, 
      mult_21_C241_n609, mult_21_C241_n608, mult_21_C241_n607, 
      mult_21_C241_n606, mult_21_C241_n605, mult_21_C241_n604, 
      mult_21_C241_n603, mult_21_C241_n602, mult_21_C241_n601, 
      mult_21_C241_n600, mult_21_C241_n599, mult_21_C241_n598, 
      mult_21_C241_n597, mult_21_C241_n596, mult_21_C241_n595, 
      mult_21_C241_n594, mult_21_C241_n593, mult_21_C241_n592, 
      mult_21_C241_n591, mult_21_C241_n590, mult_21_C241_n589, 
      mult_21_C241_n588, mult_21_C241_n587, mult_21_C241_n586, 
      mult_21_C241_n585, mult_21_C241_n584, mult_21_C241_n583, 
      mult_21_C241_n582, mult_21_C241_n581, mult_21_C241_n580, 
      mult_21_C241_n579, mult_21_C241_n578, mult_21_C241_n577, 
      mult_21_C241_n576, mult_21_C241_n575, mult_21_C241_n574, 
      mult_21_C241_n573, mult_21_C241_n572, mult_21_C241_n571, 
      mult_21_C241_n570, mult_21_C241_n569, mult_21_C241_n568, 
      mult_21_C241_n567, mult_21_C241_n566, mult_21_C241_n565, 
      mult_21_C241_n564, mult_21_C241_n563, mult_21_C241_n562, 
      mult_21_C241_n561, mult_21_C241_n560, mult_21_C241_n559, 
      mult_21_C241_n558, mult_21_C241_n557, mult_21_C241_n556, 
      mult_21_C241_n555, mult_21_C241_n554, mult_21_C241_n553, 
      mult_21_C241_n552, mult_21_C241_n551, mult_21_C241_n550, 
      mult_21_C241_n549, mult_21_C241_n548, mult_21_C241_n547, 
      mult_21_C241_n546, mult_21_C241_n545, mult_21_C241_n544, 
      mult_21_C241_n543, mult_21_C241_n542, mult_21_C241_n541, 
      mult_21_C241_n540, mult_21_C241_n539, mult_21_C241_n538, 
      mult_21_C241_n537, mult_21_C241_n536, mult_21_C241_n535, 
      mult_21_C241_n534, mult_21_C241_n533, mult_21_C241_n532, 
      mult_21_C241_n531, mult_21_C241_n530, mult_21_C241_n529, 
      mult_21_C241_n528, mult_21_C241_n527, mult_21_C241_n526, 
      mult_21_C241_n525, mult_21_C241_n524, mult_21_C241_n523, 
      mult_21_C241_n522, mult_21_C241_n521, mult_21_C241_n520, 
      mult_21_C241_n519, mult_21_C241_n518, mult_21_C241_n517, 
      mult_21_C241_n516, mult_21_C241_n515, mult_21_C241_n514, 
      mult_21_C241_n513, mult_21_C241_n512, mult_21_C241_n511, 
      mult_21_C241_n510, mult_21_C241_n509, mult_21_C241_n508, 
      mult_21_C241_n507, mult_21_C241_n506, mult_21_C241_n505, 
      mult_21_C241_n504, mult_21_C241_n503, mult_21_C241_n502, 
      mult_21_C241_n501, mult_21_C241_n500, mult_21_C241_n499, 
      mult_21_C241_n498, mult_21_C241_n497, mult_21_C241_n496, 
      mult_21_C241_n495, mult_21_C241_n494, mult_21_C241_n493, 
      mult_21_C241_n492, mult_21_C241_n491, mult_21_C241_n490, 
      mult_21_C241_n489, mult_21_C241_n488, mult_21_C241_n487, 
      mult_21_C241_n486, mult_21_C241_n485, mult_21_C241_n484, 
      mult_21_C241_n483, mult_21_C241_n482, mult_21_C241_n481, 
      mult_21_C241_n480, mult_21_C241_n479, mult_21_C241_n478, 
      mult_21_C241_n477, mult_21_C241_n476, mult_21_C241_n475, 
      mult_21_C241_n474, mult_21_C241_n473, mult_21_C241_n472, 
      mult_21_C241_n471, mult_21_C241_n470, mult_21_C241_n469, 
      mult_21_C241_n468, mult_21_C241_n467, mult_21_C241_n466, 
      mult_21_C241_n465, mult_21_C241_n464, mult_21_C241_n463, 
      mult_21_C241_n462, mult_21_C241_n461, mult_21_C241_n460, 
      mult_21_C241_n459, mult_21_C241_n458, mult_21_C241_n457, 
      mult_21_C241_n456, mult_21_C241_n455, mult_21_C241_n454, 
      mult_21_C241_n453, mult_21_C241_n452, mult_21_C241_n451, 
      mult_21_C241_n450, mult_21_C241_n449, mult_21_C241_n448, 
      mult_21_C241_n447, mult_21_C241_n446, mult_21_C241_n445, 
      mult_21_C241_n444, mult_21_C241_n443, mult_21_C241_n442, 
      mult_21_C241_n441, mult_21_C241_n440, mult_21_C241_n439, 
      mult_21_C241_n438, mult_21_C241_n437, mult_21_C241_n436, 
      mult_21_C241_n435, mult_21_C241_n434, mult_21_C241_n433, 
      mult_21_C241_n432, mult_21_C241_n431, mult_21_C241_n430, 
      mult_21_C241_n429, mult_21_C241_n428, mult_21_C241_n427, 
      mult_21_C241_n426, mult_21_C241_n425, mult_21_C241_n424, 
      mult_21_C241_n423, mult_21_C241_n422, mult_21_C241_n421, 
      mult_21_C241_n420, mult_21_C241_n419, mult_21_C241_n418, 
      mult_21_C241_n417, mult_21_C241_n416, mult_21_C241_n415, 
      mult_21_C241_n414, mult_21_C241_n413, mult_21_C241_n412, 
      mult_21_C241_n411, mult_21_C241_n410, mult_21_C241_n409, 
      mult_21_C241_n408, mult_21_C241_n407, mult_21_C241_n406, 
      mult_21_C241_n405, mult_21_C241_n404, mult_21_C241_n403, 
      mult_21_C241_n402, mult_21_C241_n401, mult_21_C241_n400, 
      mult_21_C241_n399, mult_21_C241_n398, mult_21_C241_n397, 
      mult_21_C241_n396, mult_21_C241_n395, mult_21_C241_n394, 
      mult_21_C241_n393, mult_21_C241_n392, mult_21_C241_n391, 
      mult_21_C241_n390, mult_21_C241_n389, mult_21_C241_n388, 
      mult_21_C241_n387, mult_21_C241_n386, mult_21_C241_n385, 
      mult_21_C241_n384, mult_21_C241_n383, mult_21_C241_n382, 
      mult_21_C241_n381, mult_21_C241_n380, mult_21_C241_n379, 
      mult_21_C241_n378, mult_21_C241_n377, mult_21_C241_n376, 
      mult_21_C241_n375, mult_21_C241_n374, mult_21_C241_n373, 
      mult_21_C241_n372, mult_21_C241_n371, mult_21_C241_n370, 
      mult_21_C241_n369, mult_21_C241_n368, mult_21_C241_n367, 
      mult_21_C241_n366, mult_21_C241_n365, mult_21_C241_n364, 
      mult_21_C241_n363, mult_21_C241_n362, mult_21_C241_n361, 
      mult_21_C241_n360, mult_21_C241_n359, mult_21_C241_n358, 
      mult_21_C241_n357, mult_21_C241_n356, mult_21_C241_n355, 
      mult_21_C241_n354, mult_21_C241_n353, mult_21_C241_n352, 
      mult_21_C241_n351, mult_21_C241_n350, mult_21_C241_n349, 
      mult_21_C241_n348, mult_21_C241_n347, mult_21_C241_n346, 
      mult_21_C241_n345, mult_21_C241_n344, mult_21_C241_n343, 
      mult_21_C241_n342, mult_21_C241_n341, mult_21_C241_n340, 
      mult_21_C241_n339, mult_21_C241_n338, mult_21_C241_n337, 
      mult_21_C241_n336, mult_21_C241_n335, mult_21_C241_n334, 
      mult_21_C241_n333, mult_21_C241_n332, mult_21_C241_n331, 
      mult_21_C241_n330, mult_21_C241_n329, mult_21_C241_n328, 
      mult_21_C241_n327, mult_21_C241_n326, mult_21_C241_n325, 
      mult_21_C241_n324, mult_21_C241_n323, mult_21_C241_n322, 
      mult_21_C241_n321, mult_21_C241_n320, mult_21_C241_n319, 
      mult_21_C241_n318, mult_21_C241_n317, mult_21_C241_n316, 
      mult_21_C241_n315, mult_21_C241_n314, mult_21_C241_n313, 
      mult_21_C241_n312, mult_21_C241_n311, mult_21_C241_n310, 
      mult_21_C241_n309, mult_21_C241_n308, mult_21_C241_n307, 
      mult_21_C241_n306, mult_21_C241_n305, mult_21_C241_n304, 
      mult_21_C241_n303, mult_21_C241_n302, mult_21_C241_n301, 
      mult_21_C241_n300, mult_21_C241_n299, mult_21_C241_n298, 
      mult_21_C241_n297, mult_21_C241_n296, mult_21_C241_n295, 
      mult_21_C241_n294, mult_21_C241_n293, mult_21_C241_n292, 
      mult_21_C241_n291, mult_21_C241_n290, mult_21_C241_n289, 
      mult_21_C241_n288, mult_21_C241_n287, mult_21_C241_n286, 
      mult_21_C241_n285, mult_21_C241_n284, mult_21_C241_n283, 
      mult_21_C241_n282, mult_21_C241_n281, mult_21_C241_n280, 
      mult_21_C241_n279, mult_21_C241_n278, mult_21_C241_n277, 
      mult_21_C241_n276, mult_21_C241_n275, mult_21_C241_n274, 
      mult_21_C241_n273, mult_21_C241_n272, mult_21_C241_n271, 
      mult_21_C241_n270, mult_21_C241_n269, mult_21_C241_n268, 
      mult_21_C241_n267, mult_21_C241_n266, mult_21_C241_n265, 
      mult_21_C241_n264, mult_21_C241_n263, mult_21_C241_n262, 
      mult_21_C241_n261, mult_21_C241_n260, mult_21_C241_n259, 
      mult_21_C241_n258, mult_21_C241_n257, mult_21_C241_n256, 
      mult_21_C241_n255, mult_21_C241_n254, mult_21_C241_n253, 
      mult_21_C241_n252, mult_21_C241_n251, mult_21_C241_n250, 
      mult_21_C241_n249, mult_21_C241_n248, mult_21_C241_n247, 
      mult_21_C241_n246, mult_21_C241_n245, mult_21_C241_n244, 
      mult_21_C241_n243, mult_21_C241_n242, mult_21_C241_n241, 
      mult_21_C241_n240, mult_21_C241_n239, mult_21_C241_n238, 
      mult_21_C241_n237, mult_21_C241_n236, mult_21_C241_n235, 
      mult_21_C241_n234, mult_21_C241_n233, mult_21_C241_n232, 
      mult_21_C241_n231, mult_21_C241_n230, mult_21_C241_n229, 
      mult_21_C241_n228, mult_21_C241_n227, mult_21_C241_n226, 
      mult_21_C241_n225, mult_21_C241_n224, mult_21_C241_n223, 
      mult_21_C241_n222, mult_21_C241_n221, mult_21_C241_n220, 
      mult_21_C241_n219, mult_21_C241_n218, mult_21_C241_n217, 
      mult_21_C241_n216, mult_21_C241_n215, mult_21_C241_n214, 
      mult_21_C241_n213, mult_21_C241_n212, mult_21_C241_n211, 
      mult_21_C241_n210, mult_21_C241_n209, mult_21_C241_n208, 
      mult_21_C241_n207, mult_21_C241_n206, mult_21_C241_n205, 
      mult_21_C241_n204, mult_21_C241_n203, mult_21_C241_n202, 
      mult_21_C241_n186, mult_21_C241_n185, mult_21_C241_n184, 
      mult_21_C241_n183, mult_21_C241_n182, mult_21_C241_n181, 
      mult_21_C241_n180, mult_21_C241_n179, mult_21_C241_n178, 
      mult_21_C241_n177, mult_21_C241_n176, mult_21_C241_n175, 
      mult_21_C241_n174, mult_21_C241_n173, mult_21_C241_n172, 
      mult_21_C241_n171, mult_21_C241_n170, mult_21_C241_n169, 
      mult_21_C241_n168, mult_21_C241_n167, mult_21_C241_n166, 
      mult_21_C241_n165, mult_21_C241_n164, mult_21_C241_n163, 
      mult_21_C241_n162, mult_21_C241_n161, mult_21_C241_n160, 
      mult_21_C241_n159, mult_21_C241_n158, mult_21_C241_n157, 
      mult_21_C241_n156, mult_21_C241_n104, mult_21_C241_n99, mult_21_C241_n94,
      mult_21_C241_n89, mult_21_C241_n84, mult_21_C241_n80, mult_21_C241_n73, 
      mult_21_C241_n66, mult_21_C241_n58, mult_21_C241_n50, mult_21_C241_n42, 
      mult_21_C243_n1451, mult_21_C243_n1450, mult_21_C243_n1449, 
      mult_21_C243_n1448, mult_21_C243_n1447, mult_21_C243_n1446, 
      mult_21_C243_n1445, mult_21_C243_n1444, mult_21_C243_n1443, 
      mult_21_C243_n1442, mult_21_C243_n1441, mult_21_C243_n1440, 
      mult_21_C243_n1439, mult_21_C243_n1438, mult_21_C243_n1437, 
      mult_21_C243_n1436, mult_21_C243_n1435, mult_21_C243_n1434, 
      mult_21_C243_n1433, mult_21_C243_n1432, mult_21_C243_n1431, 
      mult_21_C243_n1430, mult_21_C243_n1429, mult_21_C243_n1428, 
      mult_21_C243_n1427, mult_21_C243_n1426, mult_21_C243_n1425, 
      mult_21_C243_n1424, mult_21_C243_n1423, mult_21_C243_n1422, 
      mult_21_C243_n1421, mult_21_C243_n1420, mult_21_C243_n1419, 
      mult_21_C243_n1418, mult_21_C243_n1417, mult_21_C243_n1416, 
      mult_21_C243_n1415, mult_21_C243_n1414, mult_21_C243_n1413, 
      mult_21_C243_n1412, mult_21_C243_n1411, mult_21_C243_n1410, 
      mult_21_C243_n1409, mult_21_C243_n1408, mult_21_C243_n1407, 
      mult_21_C243_n1406, mult_21_C243_n1405, mult_21_C243_n1404, 
      mult_21_C243_n1403, mult_21_C243_n1402, mult_21_C243_n1401, 
      mult_21_C243_n1400, mult_21_C243_n1399, mult_21_C243_n1398, 
      mult_21_C243_n1397, mult_21_C243_n1396, mult_21_C243_n1395, 
      mult_21_C243_n1394, mult_21_C243_n1393, mult_21_C243_n1392, 
      mult_21_C243_n1391, mult_21_C243_n1390, mult_21_C243_n1389, 
      mult_21_C243_n1388, mult_21_C243_n1387, mult_21_C243_n1386, 
      mult_21_C243_n1385, mult_21_C243_n1384, mult_21_C243_n1383, 
      mult_21_C243_n1382, mult_21_C243_n1381, mult_21_C243_n1380, 
      mult_21_C243_n1379, mult_21_C243_n1378, mult_21_C243_n1377, 
      mult_21_C243_n1376, mult_21_C243_n1375, mult_21_C243_n1226, 
      mult_21_C243_n1225, mult_21_C243_n1224, mult_21_C243_n1223, 
      mult_21_C243_n1222, mult_21_C243_n1221, mult_21_C243_n1220, 
      mult_21_C243_n1219, mult_21_C243_n1218, mult_21_C243_n1217, 
      mult_21_C243_n1216, mult_21_C243_n1215, mult_21_C243_n1214, 
      mult_21_C243_n1213, mult_21_C243_n1212, mult_21_C243_n1211, 
      mult_21_C243_n1210, mult_21_C243_n1209, mult_21_C243_n1208, 
      mult_21_C243_n1207, mult_21_C243_n1206, mult_21_C243_n1205, 
      mult_21_C243_n1204, mult_21_C243_n1203, mult_21_C243_n1202, 
      mult_21_C243_n1201, mult_21_C243_n1200, mult_21_C243_n1199, 
      mult_21_C243_n1198, mult_21_C243_n1197, mult_21_C243_n1196, 
      mult_21_C243_n1195, mult_21_C243_n1194, mult_21_C243_n1193, 
      mult_21_C243_n1192, mult_21_C243_n1191, mult_21_C243_n1190, 
      mult_21_C243_n1189, mult_21_C243_n1188, mult_21_C243_n1187, 
      mult_21_C243_n1186, mult_21_C243_n1185, mult_21_C243_n1184, 
      mult_21_C243_n1183, mult_21_C243_n1182, mult_21_C243_n1181, 
      mult_21_C243_n1180, mult_21_C243_n1179, mult_21_C243_n1178, 
      mult_21_C243_n1177, mult_21_C243_n1176, mult_21_C243_n1175, 
      mult_21_C243_n1174, mult_21_C243_n1173, mult_21_C243_n1172, 
      mult_21_C243_n1171, mult_21_C243_n1170, mult_21_C243_n1169, 
      mult_21_C243_n1168, mult_21_C243_n1167, mult_21_C243_n1166, 
      mult_21_C243_n1165, mult_21_C243_n1164, mult_21_C243_n1163, 
      mult_21_C243_n1162, mult_21_C243_n1161, mult_21_C243_n1160, 
      mult_21_C243_n1159, mult_21_C243_n1158, mult_21_C243_n1157, 
      mult_21_C243_n1156, mult_21_C243_n1155, mult_21_C243_n1154, 
      mult_21_C243_n1153, mult_21_C243_n1152, mult_21_C243_n1151, 
      mult_21_C243_n1150, mult_21_C243_n1149, mult_21_C243_n1148, 
      mult_21_C243_n1147, mult_21_C243_n1146, mult_21_C243_n1145, 
      mult_21_C243_n1144, mult_21_C243_n1143, mult_21_C243_n1142, 
      mult_21_C243_n1141, mult_21_C243_n1140, mult_21_C243_n1139, 
      mult_21_C243_n1138, mult_21_C243_n1137, mult_21_C243_n1136, 
      mult_21_C243_n1135, mult_21_C243_n1134, mult_21_C243_n1133, 
      mult_21_C243_n1132, mult_21_C243_n1131, mult_21_C243_n1130, 
      mult_21_C243_n1129, mult_21_C243_n1128, mult_21_C243_n1127, 
      mult_21_C243_n1126, mult_21_C243_n1125, mult_21_C243_n1124, 
      mult_21_C243_n1123, mult_21_C243_n1122, mult_21_C243_n1121, 
      mult_21_C243_n1120, mult_21_C243_n1119, mult_21_C243_n1118, 
      mult_21_C243_n1117, mult_21_C243_n1116, mult_21_C243_n1115, 
      mult_21_C243_n1114, mult_21_C243_n1113, mult_21_C243_n1112, 
      mult_21_C243_n1111, mult_21_C243_n1110, mult_21_C243_n1109, 
      mult_21_C243_n1108, mult_21_C243_n1107, mult_21_C243_n1106, 
      mult_21_C243_n1105, mult_21_C243_n1104, mult_21_C243_n1103, 
      mult_21_C243_n1102, mult_21_C243_n1101, mult_21_C243_n1100, 
      mult_21_C243_n1099, mult_21_C243_n1098, mult_21_C243_n1097, 
      mult_21_C243_n1096, mult_21_C243_n1095, mult_21_C243_n1094, 
      mult_21_C243_n1093, mult_21_C243_n1092, mult_21_C243_n1091, 
      mult_21_C243_n1090, mult_21_C243_n1089, mult_21_C243_n1088, 
      mult_21_C243_n1087, mult_21_C243_n1086, mult_21_C243_n1085, 
      mult_21_C243_n1084, mult_21_C243_n1083, mult_21_C243_n1082, 
      mult_21_C243_n1081, mult_21_C243_n1080, mult_21_C243_n1079, 
      mult_21_C243_n1078, mult_21_C243_n1077, mult_21_C243_n1076, 
      mult_21_C243_n1075, mult_21_C243_n1074, mult_21_C243_n1073, 
      mult_21_C243_n1072, mult_21_C243_n1071, mult_21_C243_n1070, 
      mult_21_C243_n1069, mult_21_C243_n1068, mult_21_C243_n1067, 
      mult_21_C243_n1066, mult_21_C243_n1065, mult_21_C243_n1064, 
      mult_21_C243_n1063, mult_21_C243_n1062, mult_21_C243_n1061, 
      mult_21_C243_n1060, mult_21_C243_n1059, mult_21_C243_n1058, 
      mult_21_C243_n1057, mult_21_C243_n1056, mult_21_C243_n1055, 
      mult_21_C243_n1054, mult_21_C243_n1053, mult_21_C243_n1052, 
      mult_21_C243_n1051, mult_21_C243_n1050, mult_21_C243_n1049, 
      mult_21_C243_n1048, mult_21_C243_n1047, mult_21_C243_n1046, 
      mult_21_C243_n1045, mult_21_C243_n1044, mult_21_C243_n1043, 
      mult_21_C243_n1042, mult_21_C243_n1041, mult_21_C243_n1040, 
      mult_21_C243_n1039, mult_21_C243_n1038, mult_21_C243_n1037, 
      mult_21_C243_n1036, mult_21_C243_n1035, mult_21_C243_n1034, 
      mult_21_C243_n1033, mult_21_C243_n1032, mult_21_C243_n1031, 
      mult_21_C243_n1030, mult_21_C243_n1029, mult_21_C243_n1028, 
      mult_21_C243_n1027, mult_21_C243_n1026, mult_21_C243_n1025, 
      mult_21_C243_n1024, mult_21_C243_n1023, mult_21_C243_n1022, 
      mult_21_C243_n1021, mult_21_C243_n1020, mult_21_C243_n1019, 
      mult_21_C243_n1018, mult_21_C243_n1017, mult_21_C243_n1016, 
      mult_21_C243_n1015, mult_21_C243_n1014, mult_21_C243_n1013, 
      mult_21_C243_n1012, mult_21_C243_n1011, mult_21_C243_n1010, 
      mult_21_C243_n1009, mult_21_C243_n1008, mult_21_C243_n1007, 
      mult_21_C243_n1006, mult_21_C243_n1005, mult_21_C243_n1004, 
      mult_21_C243_n1003, mult_21_C243_n1002, mult_21_C243_n1001, 
      mult_21_C243_n1000, mult_21_C243_n999, mult_21_C243_n998, 
      mult_21_C243_n997, mult_21_C243_n996, mult_21_C243_n995, 
      mult_21_C243_n994, mult_21_C243_n993, mult_21_C243_n992, 
      mult_21_C243_n991, mult_21_C243_n990, mult_21_C243_n989, 
      mult_21_C243_n988, mult_21_C243_n987, mult_21_C243_n986, 
      mult_21_C243_n985, mult_21_C243_n984, mult_21_C243_n983, 
      mult_21_C243_n982, mult_21_C243_n981, mult_21_C243_n980, 
      mult_21_C243_n979, mult_21_C243_n978, mult_21_C243_n977, 
      mult_21_C243_n976, mult_21_C243_n975, mult_21_C243_n974, 
      mult_21_C243_n973, mult_21_C243_n972, mult_21_C243_n971, 
      mult_21_C243_n970, mult_21_C243_n969, mult_21_C243_n968, 
      mult_21_C243_n967, mult_21_C243_n966, mult_21_C243_n965, 
      mult_21_C243_n964, mult_21_C243_n963, mult_21_C243_n962, 
      mult_21_C243_n961, mult_21_C243_n960, mult_21_C243_n959, 
      mult_21_C243_n958, mult_21_C243_n957, mult_21_C243_n956, 
      mult_21_C243_n955, mult_21_C243_n953, mult_21_C243_n952, 
      mult_21_C243_n951, mult_21_C243_n950, mult_21_C243_n949, 
      mult_21_C243_n948, mult_21_C243_n947, mult_21_C243_n946, 
      mult_21_C243_n945, mult_21_C243_n944, mult_21_C243_n943, 
      mult_21_C243_n942, mult_21_C243_n941, mult_21_C243_n940, 
      mult_21_C243_n939, mult_21_C243_n923, mult_21_C243_n922, 
      mult_21_C243_n921, mult_21_C243_n920, mult_21_C243_n919, 
      mult_21_C243_n918, mult_21_C243_n917, mult_21_C243_n916, 
      mult_21_C243_n915, mult_21_C243_n914, mult_21_C243_n913, 
      mult_21_C243_n912, mult_21_C243_n911, mult_21_C243_n910, 
      mult_21_C243_n909, mult_21_C243_n908, mult_21_C243_n907, 
      mult_21_C243_n906, mult_21_C243_n905, mult_21_C243_n904, 
      mult_21_C243_n903, mult_21_C243_n902, mult_21_C243_n901, 
      mult_21_C243_n900, mult_21_C243_n899, mult_21_C243_n898, 
      mult_21_C243_n897, mult_21_C243_n896, mult_21_C243_n895, 
      mult_21_C243_n894, mult_21_C243_n893, mult_21_C243_n892, 
      mult_21_C243_n891, mult_21_C243_n890, mult_21_C243_n889, 
      mult_21_C243_n888, mult_21_C243_n887, mult_21_C243_n886, 
      mult_21_C243_n885, mult_21_C243_n884, mult_21_C243_n883, 
      mult_21_C243_n882, mult_21_C243_n881, mult_21_C243_n880, 
      mult_21_C243_n879, mult_21_C243_n878, mult_21_C243_n877, 
      mult_21_C243_n876, mult_21_C243_n875, mult_21_C243_n874, 
      mult_21_C243_n873, mult_21_C243_n872, mult_21_C243_n871, 
      mult_21_C243_n870, mult_21_C243_n869, mult_21_C243_n868, 
      mult_21_C243_n867, mult_21_C243_n866, mult_21_C243_n865, 
      mult_21_C243_n864, mult_21_C243_n863, mult_21_C243_n862, 
      mult_21_C243_n861, mult_21_C243_n860, mult_21_C243_n859, 
      mult_21_C243_n858, mult_21_C243_n857, mult_21_C243_n856, 
      mult_21_C243_n855, mult_21_C243_n854, mult_21_C243_n853, 
      mult_21_C243_n852, mult_21_C243_n851, mult_21_C243_n850, 
      mult_21_C243_n849, mult_21_C243_n848, mult_21_C243_n847, 
      mult_21_C243_n846, mult_21_C243_n845, mult_21_C243_n844, 
      mult_21_C243_n843, mult_21_C243_n842, mult_21_C243_n841, 
      mult_21_C243_n840, mult_21_C243_n839, mult_21_C243_n838, 
      mult_21_C243_n837, mult_21_C243_n836, mult_21_C243_n835, 
      mult_21_C243_n834, mult_21_C243_n833, mult_21_C243_n832, 
      mult_21_C243_n831, mult_21_C243_n830, mult_21_C243_n829, 
      mult_21_C243_n828, mult_21_C243_n827, mult_21_C243_n826, 
      mult_21_C243_n825, mult_21_C243_n824, mult_21_C243_n823, 
      mult_21_C243_n822, mult_21_C243_n821, mult_21_C243_n820, 
      mult_21_C243_n819, mult_21_C243_n818, mult_21_C243_n817, 
      mult_21_C243_n816, mult_21_C243_n815, mult_21_C243_n814, 
      mult_21_C243_n813, mult_21_C243_n812, mult_21_C243_n811, 
      mult_21_C243_n810, mult_21_C243_n809, mult_21_C243_n808, 
      mult_21_C243_n807, mult_21_C243_n806, mult_21_C243_n805, 
      mult_21_C243_n804, mult_21_C243_n803, mult_21_C243_n802, 
      mult_21_C243_n801, mult_21_C243_n800, mult_21_C243_n799, 
      mult_21_C243_n798, mult_21_C243_n797, mult_21_C243_n796, 
      mult_21_C243_n795, mult_21_C243_n794, mult_21_C243_n793, 
      mult_21_C243_n792, mult_21_C243_n791, mult_21_C243_n790, 
      mult_21_C243_n789, mult_21_C243_n788, mult_21_C243_n787, 
      mult_21_C243_n786, mult_21_C243_n785, mult_21_C243_n784, 
      mult_21_C243_n783, mult_21_C243_n782, mult_21_C243_n781, 
      mult_21_C243_n780, mult_21_C243_n779, mult_21_C243_n778, 
      mult_21_C243_n777, mult_21_C243_n776, mult_21_C243_n775, 
      mult_21_C243_n774, mult_21_C243_n773, mult_21_C243_n772, 
      mult_21_C243_n771, mult_21_C243_n770, mult_21_C243_n769, 
      mult_21_C243_n768, mult_21_C243_n767, mult_21_C243_n766, 
      mult_21_C243_n765, mult_21_C243_n764, mult_21_C243_n763, 
      mult_21_C243_n762, mult_21_C243_n761, mult_21_C243_n760, 
      mult_21_C243_n759, mult_21_C243_n758, mult_21_C243_n757, 
      mult_21_C243_n756, mult_21_C243_n755, mult_21_C243_n754, 
      mult_21_C243_n753, mult_21_C243_n752, mult_21_C243_n751, 
      mult_21_C243_n750, mult_21_C243_n749, mult_21_C243_n748, 
      mult_21_C243_n747, mult_21_C243_n746, mult_21_C243_n745, 
      mult_21_C243_n744, mult_21_C243_n743, mult_21_C243_n742, 
      mult_21_C243_n741, mult_21_C243_n740, mult_21_C243_n739, 
      mult_21_C243_n738, mult_21_C243_n737, mult_21_C243_n736, 
      mult_21_C243_n735, mult_21_C243_n734, mult_21_C243_n733, 
      mult_21_C243_n732, mult_21_C243_n731, mult_21_C243_n730, 
      mult_21_C243_n729, mult_21_C243_n728, mult_21_C243_n727, 
      mult_21_C243_n726, mult_21_C243_n725, mult_21_C243_n724, 
      mult_21_C243_n723, mult_21_C243_n722, mult_21_C243_n721, 
      mult_21_C243_n720, mult_21_C243_n719, mult_21_C243_n718, 
      mult_21_C243_n717, mult_21_C243_n716, mult_21_C243_n715, 
      mult_21_C243_n714, mult_21_C243_n713, mult_21_C243_n712, 
      mult_21_C243_n711, mult_21_C243_n710, mult_21_C243_n709, 
      mult_21_C243_n708, mult_21_C243_n707, mult_21_C243_n706, 
      mult_21_C243_n705, mult_21_C243_n704, mult_21_C243_n703, 
      mult_21_C243_n702, mult_21_C243_n701, mult_21_C243_n700, 
      mult_21_C243_n699, mult_21_C243_n698, mult_21_C243_n697, 
      mult_21_C243_n696, mult_21_C243_n695, mult_21_C243_n694, 
      mult_21_C243_n693, mult_21_C243_n692, mult_21_C243_n691, 
      mult_21_C243_n690, mult_21_C243_n689, mult_21_C243_n688, 
      mult_21_C243_n687, mult_21_C243_n686, mult_21_C243_n685, 
      mult_21_C243_n684, mult_21_C243_n683, mult_21_C243_n682, 
      mult_21_C243_n681, mult_21_C243_n680, mult_21_C243_n679, 
      mult_21_C243_n678, mult_21_C243_n677, mult_21_C243_n676, 
      mult_21_C243_n675, mult_21_C243_n674, mult_21_C243_n673, 
      mult_21_C243_n672, mult_21_C243_n671, mult_21_C243_n670, 
      mult_21_C243_n669, mult_21_C243_n668, mult_21_C243_n667, 
      mult_21_C243_n666, mult_21_C243_n665, mult_21_C243_n664, 
      mult_21_C243_n663, mult_21_C243_n662, mult_21_C243_n661, 
      mult_21_C243_n660, mult_21_C243_n659, mult_21_C243_n658, 
      mult_21_C243_n657, mult_21_C243_n656, mult_21_C243_n655, 
      mult_21_C243_n654, mult_21_C243_n653, mult_21_C243_n652, 
      mult_21_C243_n651, mult_21_C243_n650, mult_21_C243_n649, 
      mult_21_C243_n648, mult_21_C243_n647, mult_21_C243_n646, 
      mult_21_C243_n645, mult_21_C243_n644, mult_21_C243_n643, 
      mult_21_C243_n642, mult_21_C243_n641, mult_21_C243_n640, 
      mult_21_C243_n639, mult_21_C243_n638, mult_21_C243_n637, 
      mult_21_C243_n636, mult_21_C243_n635, mult_21_C243_n634, 
      mult_21_C243_n633, mult_21_C243_n632, mult_21_C243_n631, 
      mult_21_C243_n630, mult_21_C243_n629, mult_21_C243_n628, 
      mult_21_C243_n627, mult_21_C243_n626, mult_21_C243_n625, 
      mult_21_C243_n624, mult_21_C243_n623, mult_21_C243_n622, 
      mult_21_C243_n621, mult_21_C243_n620, mult_21_C243_n619, 
      mult_21_C243_n618, mult_21_C243_n617, mult_21_C243_n616, 
      mult_21_C243_n615, mult_21_C243_n614, mult_21_C243_n613, 
      mult_21_C243_n612, mult_21_C243_n611, mult_21_C243_n610, 
      mult_21_C243_n609, mult_21_C243_n608, mult_21_C243_n607, 
      mult_21_C243_n606, mult_21_C243_n605, mult_21_C243_n604, 
      mult_21_C243_n603, mult_21_C243_n602, mult_21_C243_n601, 
      mult_21_C243_n600, mult_21_C243_n599, mult_21_C243_n598, 
      mult_21_C243_n597, mult_21_C243_n596, mult_21_C243_n595, 
      mult_21_C243_n594, mult_21_C243_n593, mult_21_C243_n592, 
      mult_21_C243_n591, mult_21_C243_n590, mult_21_C243_n589, 
      mult_21_C243_n588, mult_21_C243_n587, mult_21_C243_n586, 
      mult_21_C243_n585, mult_21_C243_n584, mult_21_C243_n583, 
      mult_21_C243_n582, mult_21_C243_n581, mult_21_C243_n580, 
      mult_21_C243_n579, mult_21_C243_n578, mult_21_C243_n577, 
      mult_21_C243_n576, mult_21_C243_n575, mult_21_C243_n574, 
      mult_21_C243_n573, mult_21_C243_n572, mult_21_C243_n571, 
      mult_21_C243_n570, mult_21_C243_n569, mult_21_C243_n568, 
      mult_21_C243_n567, mult_21_C243_n566, mult_21_C243_n565, 
      mult_21_C243_n564, mult_21_C243_n563, mult_21_C243_n562, 
      mult_21_C243_n561, mult_21_C243_n560, mult_21_C243_n559, 
      mult_21_C243_n558, mult_21_C243_n557, mult_21_C243_n556, 
      mult_21_C243_n555, mult_21_C243_n554, mult_21_C243_n553, 
      mult_21_C243_n552, mult_21_C243_n551, mult_21_C243_n550, 
      mult_21_C243_n549, mult_21_C243_n548, mult_21_C243_n547, 
      mult_21_C243_n546, mult_21_C243_n545, mult_21_C243_n544, 
      mult_21_C243_n543, mult_21_C243_n542, mult_21_C243_n541, 
      mult_21_C243_n540, mult_21_C243_n539, mult_21_C243_n538, 
      mult_21_C243_n537, mult_21_C243_n536, mult_21_C243_n535, 
      mult_21_C243_n534, mult_21_C243_n533, mult_21_C243_n532, 
      mult_21_C243_n531, mult_21_C243_n530, mult_21_C243_n529, 
      mult_21_C243_n528, mult_21_C243_n527, mult_21_C243_n526, 
      mult_21_C243_n525, mult_21_C243_n524, mult_21_C243_n523, 
      mult_21_C243_n522, mult_21_C243_n521, mult_21_C243_n520, 
      mult_21_C243_n519, mult_21_C243_n518, mult_21_C243_n517, 
      mult_21_C243_n516, mult_21_C243_n515, mult_21_C243_n514, 
      mult_21_C243_n513, mult_21_C243_n512, mult_21_C243_n511, 
      mult_21_C243_n510, mult_21_C243_n509, mult_21_C243_n508, 
      mult_21_C243_n507, mult_21_C243_n506, mult_21_C243_n505, 
      mult_21_C243_n504, mult_21_C243_n503, mult_21_C243_n502, 
      mult_21_C243_n501, mult_21_C243_n500, mult_21_C243_n499, 
      mult_21_C243_n498, mult_21_C243_n497, mult_21_C243_n496, 
      mult_21_C243_n495, mult_21_C243_n494, mult_21_C243_n493, 
      mult_21_C243_n492, mult_21_C243_n491, mult_21_C243_n490, 
      mult_21_C243_n489, mult_21_C243_n488, mult_21_C243_n487, 
      mult_21_C243_n486, mult_21_C243_n485, mult_21_C243_n484, 
      mult_21_C243_n483, mult_21_C243_n482, mult_21_C243_n481, 
      mult_21_C243_n480, mult_21_C243_n479, mult_21_C243_n478, 
      mult_21_C243_n477, mult_21_C243_n476, mult_21_C243_n475, 
      mult_21_C243_n474, mult_21_C243_n473, mult_21_C243_n472, 
      mult_21_C243_n471, mult_21_C243_n470, mult_21_C243_n469, 
      mult_21_C243_n468, mult_21_C243_n467, mult_21_C243_n466, 
      mult_21_C243_n465, mult_21_C243_n464, mult_21_C243_n463, 
      mult_21_C243_n462, mult_21_C243_n461, mult_21_C243_n460, 
      mult_21_C243_n459, mult_21_C243_n458, mult_21_C243_n457, 
      mult_21_C243_n456, mult_21_C243_n455, mult_21_C243_n454, 
      mult_21_C243_n453, mult_21_C243_n452, mult_21_C243_n451, 
      mult_21_C243_n450, mult_21_C243_n449, mult_21_C243_n448, 
      mult_21_C243_n447, mult_21_C243_n446, mult_21_C243_n445, 
      mult_21_C243_n444, mult_21_C243_n443, mult_21_C243_n442, 
      mult_21_C243_n441, mult_21_C243_n440, mult_21_C243_n439, 
      mult_21_C243_n438, mult_21_C243_n437, mult_21_C243_n436, 
      mult_21_C243_n435, mult_21_C243_n434, mult_21_C243_n433, 
      mult_21_C243_n432, mult_21_C243_n431, mult_21_C243_n430, 
      mult_21_C243_n429, mult_21_C243_n428, mult_21_C243_n427, 
      mult_21_C243_n426, mult_21_C243_n425, mult_21_C243_n424, 
      mult_21_C243_n423, mult_21_C243_n422, mult_21_C243_n421, 
      mult_21_C243_n420, mult_21_C243_n419, mult_21_C243_n418, 
      mult_21_C243_n417, mult_21_C243_n416, mult_21_C243_n415, 
      mult_21_C243_n414, mult_21_C243_n413, mult_21_C243_n412, 
      mult_21_C243_n411, mult_21_C243_n410, mult_21_C243_n409, 
      mult_21_C243_n408, mult_21_C243_n407, mult_21_C243_n406, 
      mult_21_C243_n405, mult_21_C243_n404, mult_21_C243_n403, 
      mult_21_C243_n402, mult_21_C243_n401, mult_21_C243_n400, 
      mult_21_C243_n399, mult_21_C243_n398, mult_21_C243_n397, 
      mult_21_C243_n396, mult_21_C243_n395, mult_21_C243_n394, 
      mult_21_C243_n393, mult_21_C243_n392, mult_21_C243_n391, 
      mult_21_C243_n390, mult_21_C243_n389, mult_21_C243_n388, 
      mult_21_C243_n387, mult_21_C243_n386, mult_21_C243_n385, 
      mult_21_C243_n384, mult_21_C243_n383, mult_21_C243_n382, 
      mult_21_C243_n381, mult_21_C243_n380, mult_21_C243_n379, 
      mult_21_C243_n378, mult_21_C243_n377, mult_21_C243_n376, 
      mult_21_C243_n375, mult_21_C243_n374, mult_21_C243_n373, 
      mult_21_C243_n372, mult_21_C243_n371, mult_21_C243_n370, 
      mult_21_C243_n369, mult_21_C243_n368, mult_21_C243_n367, 
      mult_21_C243_n366, mult_21_C243_n365, mult_21_C243_n364, 
      mult_21_C243_n363, mult_21_C243_n362, mult_21_C243_n361, 
      mult_21_C243_n360, mult_21_C243_n359, mult_21_C243_n358, 
      mult_21_C243_n357, mult_21_C243_n356, mult_21_C243_n355, 
      mult_21_C243_n354, mult_21_C243_n353, mult_21_C243_n352, 
      mult_21_C243_n351, mult_21_C243_n350, mult_21_C243_n349, 
      mult_21_C243_n348, mult_21_C243_n347, mult_21_C243_n346, 
      mult_21_C243_n345, mult_21_C243_n344, mult_21_C243_n343, 
      mult_21_C243_n342, mult_21_C243_n341, mult_21_C243_n340, 
      mult_21_C243_n339, mult_21_C243_n338, mult_21_C243_n337, 
      mult_21_C243_n336, mult_21_C243_n335, mult_21_C243_n334, 
      mult_21_C243_n333, mult_21_C243_n332, mult_21_C243_n331, 
      mult_21_C243_n330, mult_21_C243_n329, mult_21_C243_n328, 
      mult_21_C243_n327, mult_21_C243_n326, mult_21_C243_n325, 
      mult_21_C243_n324, mult_21_C243_n323, mult_21_C243_n322, 
      mult_21_C243_n321, mult_21_C243_n320, mult_21_C243_n319, 
      mult_21_C243_n318, mult_21_C243_n317, mult_21_C243_n316, 
      mult_21_C243_n315, mult_21_C243_n314, mult_21_C243_n313, 
      mult_21_C243_n312, mult_21_C243_n311, mult_21_C243_n310, 
      mult_21_C243_n309, mult_21_C243_n308, mult_21_C243_n307, 
      mult_21_C243_n306, mult_21_C243_n305, mult_21_C243_n304, 
      mult_21_C243_n303, mult_21_C243_n302, mult_21_C243_n301, 
      mult_21_C243_n300, mult_21_C243_n299, mult_21_C243_n298, 
      mult_21_C243_n297, mult_21_C243_n296, mult_21_C243_n295, 
      mult_21_C243_n294, mult_21_C243_n293, mult_21_C243_n292, 
      mult_21_C243_n291, mult_21_C243_n290, mult_21_C243_n289, 
      mult_21_C243_n288, mult_21_C243_n287, mult_21_C243_n286, 
      mult_21_C243_n285, mult_21_C243_n284, mult_21_C243_n283, 
      mult_21_C243_n282, mult_21_C243_n281, mult_21_C243_n280, 
      mult_21_C243_n279, mult_21_C243_n278, mult_21_C243_n277, 
      mult_21_C243_n276, mult_21_C243_n275, mult_21_C243_n274, 
      mult_21_C243_n273, mult_21_C243_n272, mult_21_C243_n271, 
      mult_21_C243_n270, mult_21_C243_n269, mult_21_C243_n268, 
      mult_21_C243_n267, mult_21_C243_n266, mult_21_C243_n265, 
      mult_21_C243_n264, mult_21_C243_n263, mult_21_C243_n262, 
      mult_21_C243_n261, mult_21_C243_n260, mult_21_C243_n259, 
      mult_21_C243_n258, mult_21_C243_n257, mult_21_C243_n256, 
      mult_21_C243_n255, mult_21_C243_n254, mult_21_C243_n253, 
      mult_21_C243_n252, mult_21_C243_n251, mult_21_C243_n250, 
      mult_21_C243_n249, mult_21_C243_n248, mult_21_C243_n247, 
      mult_21_C243_n246, mult_21_C243_n245, mult_21_C243_n244, 
      mult_21_C243_n243, mult_21_C243_n242, mult_21_C243_n241, 
      mult_21_C243_n240, mult_21_C243_n239, mult_21_C243_n238, 
      mult_21_C243_n237, mult_21_C243_n236, mult_21_C243_n235, 
      mult_21_C243_n234, mult_21_C243_n233, mult_21_C243_n232, 
      mult_21_C243_n231, mult_21_C243_n230, mult_21_C243_n229, 
      mult_21_C243_n228, mult_21_C243_n227, mult_21_C243_n226, 
      mult_21_C243_n225, mult_21_C243_n224, mult_21_C243_n223, 
      mult_21_C243_n222, mult_21_C243_n221, mult_21_C243_n220, 
      mult_21_C243_n219, mult_21_C243_n218, mult_21_C243_n217, 
      mult_21_C243_n216, mult_21_C243_n215, mult_21_C243_n214, 
      mult_21_C243_n213, mult_21_C243_n212, mult_21_C243_n211, 
      mult_21_C243_n210, mult_21_C243_n209, mult_21_C243_n208, 
      mult_21_C243_n207, mult_21_C243_n206, mult_21_C243_n205, 
      mult_21_C243_n204, mult_21_C243_n203, mult_21_C243_n202, 
      mult_21_C243_n186, mult_21_C243_n185, mult_21_C243_n184, 
      mult_21_C243_n183, mult_21_C243_n182, mult_21_C243_n181, 
      mult_21_C243_n180, mult_21_C243_n179, mult_21_C243_n178, 
      mult_21_C243_n177, mult_21_C243_n176, mult_21_C243_n175, 
      mult_21_C243_n174, mult_21_C243_n173, mult_21_C243_n172, 
      mult_21_C243_n171, mult_21_C243_n170, mult_21_C243_n169, 
      mult_21_C243_n168, mult_21_C243_n167, mult_21_C243_n166, 
      mult_21_C243_n165, mult_21_C243_n164, mult_21_C243_n163, 
      mult_21_C243_n162, mult_21_C243_n161, mult_21_C243_n160, 
      mult_21_C243_n159, mult_21_C243_n158, mult_21_C243_n157, 
      mult_21_C243_n156, mult_21_C243_n104, mult_21_C243_n99, mult_21_C243_n94,
      mult_21_C243_n89, mult_21_C243_n84, mult_21_C243_n80, mult_21_C243_n73, 
      mult_21_C243_n66, mult_21_C243_n58, mult_21_C243_n50, mult_21_C243_n42, 
      mult_21_C245_n1448, mult_21_C245_n1447, mult_21_C245_n1446, 
      mult_21_C245_n1445, mult_21_C245_n1444, mult_21_C245_n1443, 
      mult_21_C245_n1442, mult_21_C245_n1441, mult_21_C245_n1440, 
      mult_21_C245_n1439, mult_21_C245_n1438, mult_21_C245_n1437, 
      mult_21_C245_n1436, mult_21_C245_n1435, mult_21_C245_n1434, 
      mult_21_C245_n1433, mult_21_C245_n1432, mult_21_C245_n1431, 
      mult_21_C245_n1430, mult_21_C245_n1429, mult_21_C245_n1428, 
      mult_21_C245_n1427, mult_21_C245_n1426, mult_21_C245_n1425, 
      mult_21_C245_n1424, mult_21_C245_n1423, mult_21_C245_n1422, 
      mult_21_C245_n1421, mult_21_C245_n1420, mult_21_C245_n1419, 
      mult_21_C245_n1418, mult_21_C245_n1417, mult_21_C245_n1416, 
      mult_21_C245_n1415, mult_21_C245_n1414, mult_21_C245_n1413, 
      mult_21_C245_n1412, mult_21_C245_n1411, mult_21_C245_n1410, 
      mult_21_C245_n1409, mult_21_C245_n1408, mult_21_C245_n1407, 
      mult_21_C245_n1406, mult_21_C245_n1405, mult_21_C245_n1404, 
      mult_21_C245_n1403, mult_21_C245_n1402, mult_21_C245_n1401, 
      mult_21_C245_n1400, mult_21_C245_n1399, mult_21_C245_n1398, 
      mult_21_C245_n1397, mult_21_C245_n1396, mult_21_C245_n1395, 
      mult_21_C245_n1394, mult_21_C245_n1393, mult_21_C245_n1392, 
      mult_21_C245_n1391, mult_21_C245_n1390, mult_21_C245_n1389, 
      mult_21_C245_n1388, mult_21_C245_n1387, mult_21_C245_n1386, 
      mult_21_C245_n1385, mult_21_C245_n1384, mult_21_C245_n1383, 
      mult_21_C245_n1382, mult_21_C245_n1381, mult_21_C245_n1380, 
      mult_21_C245_n1379, mult_21_C245_n1378, mult_21_C245_n1377, 
      mult_21_C245_n1376, mult_21_C245_n1375, mult_21_C245_n1226, 
      mult_21_C245_n1225, mult_21_C245_n1224, mult_21_C245_n1223, 
      mult_21_C245_n1222, mult_21_C245_n1221, mult_21_C245_n1220, 
      mult_21_C245_n1219, mult_21_C245_n1218, mult_21_C245_n1217, 
      mult_21_C245_n1216, mult_21_C245_n1215, mult_21_C245_n1214, 
      mult_21_C245_n1213, mult_21_C245_n1212, mult_21_C245_n1211, 
      mult_21_C245_n1210, mult_21_C245_n1209, mult_21_C245_n1208, 
      mult_21_C245_n1207, mult_21_C245_n1206, mult_21_C245_n1205, 
      mult_21_C245_n1204, mult_21_C245_n1203, mult_21_C245_n1202, 
      mult_21_C245_n1201, mult_21_C245_n1200, mult_21_C245_n1199, 
      mult_21_C245_n1198, mult_21_C245_n1197, mult_21_C245_n1196, 
      mult_21_C245_n1195, mult_21_C245_n1194, mult_21_C245_n1193, 
      mult_21_C245_n1192, mult_21_C245_n1191, mult_21_C245_n1190, 
      mult_21_C245_n1189, mult_21_C245_n1188, mult_21_C245_n1187, 
      mult_21_C245_n1186, mult_21_C245_n1185, mult_21_C245_n1184, 
      mult_21_C245_n1183, mult_21_C245_n1182, mult_21_C245_n1181, 
      mult_21_C245_n1180, mult_21_C245_n1179, mult_21_C245_n1178, 
      mult_21_C245_n1177, mult_21_C245_n1176, mult_21_C245_n1175, 
      mult_21_C245_n1174, mult_21_C245_n1173, mult_21_C245_n1172, 
      mult_21_C245_n1171, mult_21_C245_n1170, mult_21_C245_n1169, 
      mult_21_C245_n1168, mult_21_C245_n1167, mult_21_C245_n1166, 
      mult_21_C245_n1165, mult_21_C245_n1164, mult_21_C245_n1163, 
      mult_21_C245_n1162, mult_21_C245_n1161, mult_21_C245_n1160, 
      mult_21_C245_n1159, mult_21_C245_n1158, mult_21_C245_n1157, 
      mult_21_C245_n1156, mult_21_C245_n1155, mult_21_C245_n1154, 
      mult_21_C245_n1153, mult_21_C245_n1152, mult_21_C245_n1151, 
      mult_21_C245_n1150, mult_21_C245_n1149, mult_21_C245_n1148, 
      mult_21_C245_n1147, mult_21_C245_n1146, mult_21_C245_n1145, 
      mult_21_C245_n1144, mult_21_C245_n1143, mult_21_C245_n1142, 
      mult_21_C245_n1141, mult_21_C245_n1140, mult_21_C245_n1139, 
      mult_21_C245_n1138, mult_21_C245_n1137, mult_21_C245_n1136, 
      mult_21_C245_n1135, mult_21_C245_n1134, mult_21_C245_n1133, 
      mult_21_C245_n1132, mult_21_C245_n1131, mult_21_C245_n1130, 
      mult_21_C245_n1129, mult_21_C245_n1128, mult_21_C245_n1127, 
      mult_21_C245_n1126, mult_21_C245_n1125, mult_21_C245_n1124, 
      mult_21_C245_n1123, mult_21_C245_n1122, mult_21_C245_n1121, 
      mult_21_C245_n1120, mult_21_C245_n1119, mult_21_C245_n1118, 
      mult_21_C245_n1117, mult_21_C245_n1116, mult_21_C245_n1115, 
      mult_21_C245_n1114, mult_21_C245_n1113, mult_21_C245_n1112, 
      mult_21_C245_n1111, mult_21_C245_n1110, mult_21_C245_n1109, 
      mult_21_C245_n1108, mult_21_C245_n1107, mult_21_C245_n1106, 
      mult_21_C245_n1105, mult_21_C245_n1104, mult_21_C245_n1103, 
      mult_21_C245_n1102, mult_21_C245_n1101, mult_21_C245_n1100, 
      mult_21_C245_n1099, mult_21_C245_n1098, mult_21_C245_n1097, 
      mult_21_C245_n1096, mult_21_C245_n1095, mult_21_C245_n1094, 
      mult_21_C245_n1093, mult_21_C245_n1092, mult_21_C245_n1091, 
      mult_21_C245_n1090, mult_21_C245_n1089, mult_21_C245_n1088, 
      mult_21_C245_n1087, mult_21_C245_n1086, mult_21_C245_n1085, 
      mult_21_C245_n1084, mult_21_C245_n1083, mult_21_C245_n1082, 
      mult_21_C245_n1081, mult_21_C245_n1080, mult_21_C245_n1079, 
      mult_21_C245_n1078, mult_21_C245_n1077, mult_21_C245_n1076, 
      mult_21_C245_n1075, mult_21_C245_n1074, mult_21_C245_n1073, 
      mult_21_C245_n1072, mult_21_C245_n1071, mult_21_C245_n1070, 
      mult_21_C245_n1069, mult_21_C245_n1068, mult_21_C245_n1067, 
      mult_21_C245_n1066, mult_21_C245_n1065, mult_21_C245_n1064, 
      mult_21_C245_n1063, mult_21_C245_n1062, mult_21_C245_n1061, 
      mult_21_C245_n1060, mult_21_C245_n1059, mult_21_C245_n1058, 
      mult_21_C245_n1057, mult_21_C245_n1056, mult_21_C245_n1055, 
      mult_21_C245_n1054, mult_21_C245_n1053, mult_21_C245_n1052, 
      mult_21_C245_n1051, mult_21_C245_n1050, mult_21_C245_n1049, 
      mult_21_C245_n1048, mult_21_C245_n1047, mult_21_C245_n1046, 
      mult_21_C245_n1045, mult_21_C245_n1044, mult_21_C245_n1043, 
      mult_21_C245_n1042, mult_21_C245_n1041, mult_21_C245_n1040, 
      mult_21_C245_n1039, mult_21_C245_n1038, mult_21_C245_n1037, 
      mult_21_C245_n1036, mult_21_C245_n1035, mult_21_C245_n1034, 
      mult_21_C245_n1033, mult_21_C245_n1032, mult_21_C245_n1031, 
      mult_21_C245_n1030, mult_21_C245_n1029, mult_21_C245_n1028, 
      mult_21_C245_n1027, mult_21_C245_n1026, mult_21_C245_n1025, 
      mult_21_C245_n1024, mult_21_C245_n1023, mult_21_C245_n1022, 
      mult_21_C245_n1021, mult_21_C245_n1020, mult_21_C245_n1019, 
      mult_21_C245_n1018, mult_21_C245_n1017, mult_21_C245_n1016, 
      mult_21_C245_n1015, mult_21_C245_n1014, mult_21_C245_n1013, 
      mult_21_C245_n1012, mult_21_C245_n1011, mult_21_C245_n1010, 
      mult_21_C245_n1009, mult_21_C245_n1008, mult_21_C245_n1007, 
      mult_21_C245_n1006, mult_21_C245_n1005, mult_21_C245_n1004, 
      mult_21_C245_n1003, mult_21_C245_n1002, mult_21_C245_n1001, 
      mult_21_C245_n1000, mult_21_C245_n999, mult_21_C245_n998, 
      mult_21_C245_n997, mult_21_C245_n996, mult_21_C245_n995, 
      mult_21_C245_n994, mult_21_C245_n993, mult_21_C245_n992, 
      mult_21_C245_n991, mult_21_C245_n990, mult_21_C245_n989, 
      mult_21_C245_n988, mult_21_C245_n987, mult_21_C245_n986, 
      mult_21_C245_n985, mult_21_C245_n984, mult_21_C245_n983, 
      mult_21_C245_n982, mult_21_C245_n981, mult_21_C245_n980, 
      mult_21_C245_n979, mult_21_C245_n978, mult_21_C245_n977, 
      mult_21_C245_n976, mult_21_C245_n975, mult_21_C245_n974, 
      mult_21_C245_n973, mult_21_C245_n972, mult_21_C245_n971, 
      mult_21_C245_n970, mult_21_C245_n969, mult_21_C245_n968, 
      mult_21_C245_n967, mult_21_C245_n966, mult_21_C245_n965, 
      mult_21_C245_n964, mult_21_C245_n963, mult_21_C245_n962, 
      mult_21_C245_n961, mult_21_C245_n960, mult_21_C245_n959, 
      mult_21_C245_n958, mult_21_C245_n957, mult_21_C245_n956, 
      mult_21_C245_n955, mult_21_C245_n953, mult_21_C245_n952, 
      mult_21_C245_n951, mult_21_C245_n950, mult_21_C245_n949, 
      mult_21_C245_n948, mult_21_C245_n947, mult_21_C245_n946, 
      mult_21_C245_n945, mult_21_C245_n944, mult_21_C245_n943, 
      mult_21_C245_n942, mult_21_C245_n941, mult_21_C245_n940, 
      mult_21_C245_n939, mult_21_C245_n923, mult_21_C245_n922, 
      mult_21_C245_n921, mult_21_C245_n920, mult_21_C245_n919, 
      mult_21_C245_n918, mult_21_C245_n917, mult_21_C245_n916, 
      mult_21_C245_n915, mult_21_C245_n914, mult_21_C245_n913, 
      mult_21_C245_n912, mult_21_C245_n911, mult_21_C245_n910, 
      mult_21_C245_n909, mult_21_C245_n908, mult_21_C245_n907, 
      mult_21_C245_n906, mult_21_C245_n905, mult_21_C245_n904, 
      mult_21_C245_n903, mult_21_C245_n902, mult_21_C245_n901, 
      mult_21_C245_n900, mult_21_C245_n899, mult_21_C245_n898, 
      mult_21_C245_n897, mult_21_C245_n896, mult_21_C245_n895, 
      mult_21_C245_n894, mult_21_C245_n893, mult_21_C245_n892, 
      mult_21_C245_n891, mult_21_C245_n890, mult_21_C245_n889, 
      mult_21_C245_n888, mult_21_C245_n887, mult_21_C245_n886, 
      mult_21_C245_n885, mult_21_C245_n884, mult_21_C245_n883, 
      mult_21_C245_n882, mult_21_C245_n881, mult_21_C245_n880, 
      mult_21_C245_n879, mult_21_C245_n878, mult_21_C245_n877, 
      mult_21_C245_n876, mult_21_C245_n875, mult_21_C245_n874, 
      mult_21_C245_n873, mult_21_C245_n872, mult_21_C245_n871, 
      mult_21_C245_n870, mult_21_C245_n869, mult_21_C245_n868, 
      mult_21_C245_n867, mult_21_C245_n866, mult_21_C245_n865, 
      mult_21_C245_n864, mult_21_C245_n863, mult_21_C245_n862, 
      mult_21_C245_n861, mult_21_C245_n860, mult_21_C245_n859, 
      mult_21_C245_n858, mult_21_C245_n857, mult_21_C245_n856, 
      mult_21_C245_n855, mult_21_C245_n854, mult_21_C245_n853, 
      mult_21_C245_n852, mult_21_C245_n851, mult_21_C245_n850, 
      mult_21_C245_n849, mult_21_C245_n848, mult_21_C245_n847, 
      mult_21_C245_n846, mult_21_C245_n845, mult_21_C245_n844, 
      mult_21_C245_n843, mult_21_C245_n842, mult_21_C245_n841, 
      mult_21_C245_n840, mult_21_C245_n839, mult_21_C245_n838, 
      mult_21_C245_n837, mult_21_C245_n836, mult_21_C245_n835, 
      mult_21_C245_n834, mult_21_C245_n833, mult_21_C245_n832, 
      mult_21_C245_n831, mult_21_C245_n830, mult_21_C245_n829, 
      mult_21_C245_n828, mult_21_C245_n827, mult_21_C245_n826, 
      mult_21_C245_n825, mult_21_C245_n824, mult_21_C245_n823, 
      mult_21_C245_n822, mult_21_C245_n821, mult_21_C245_n820, 
      mult_21_C245_n819, mult_21_C245_n818, mult_21_C245_n817, 
      mult_21_C245_n816, mult_21_C245_n815, mult_21_C245_n814, 
      mult_21_C245_n813, mult_21_C245_n812, mult_21_C245_n811, 
      mult_21_C245_n810, mult_21_C245_n809, mult_21_C245_n808, 
      mult_21_C245_n807, mult_21_C245_n806, mult_21_C245_n805, 
      mult_21_C245_n804, mult_21_C245_n803, mult_21_C245_n802, 
      mult_21_C245_n801, mult_21_C245_n800, mult_21_C245_n799, 
      mult_21_C245_n798, mult_21_C245_n797, mult_21_C245_n796, 
      mult_21_C245_n795, mult_21_C245_n794, mult_21_C245_n793, 
      mult_21_C245_n792, mult_21_C245_n791, mult_21_C245_n790, 
      mult_21_C245_n789, mult_21_C245_n788, mult_21_C245_n787, 
      mult_21_C245_n786, mult_21_C245_n785, mult_21_C245_n784, 
      mult_21_C245_n783, mult_21_C245_n782, mult_21_C245_n781, 
      mult_21_C245_n780, mult_21_C245_n779, mult_21_C245_n778, 
      mult_21_C245_n777, mult_21_C245_n776, mult_21_C245_n775, 
      mult_21_C245_n774, mult_21_C245_n773, mult_21_C245_n772, 
      mult_21_C245_n771, mult_21_C245_n770, mult_21_C245_n769, 
      mult_21_C245_n768, mult_21_C245_n767, mult_21_C245_n766, 
      mult_21_C245_n765, mult_21_C245_n764, mult_21_C245_n763, 
      mult_21_C245_n762, mult_21_C245_n761, mult_21_C245_n760, 
      mult_21_C245_n759, mult_21_C245_n758, mult_21_C245_n757, 
      mult_21_C245_n756, mult_21_C245_n755, mult_21_C245_n754, 
      mult_21_C245_n753, mult_21_C245_n752, mult_21_C245_n751, 
      mult_21_C245_n750, mult_21_C245_n749, mult_21_C245_n748, 
      mult_21_C245_n747, mult_21_C245_n746, mult_21_C245_n745, 
      mult_21_C245_n744, mult_21_C245_n743, mult_21_C245_n742, 
      mult_21_C245_n741, mult_21_C245_n740, mult_21_C245_n739, 
      mult_21_C245_n738, mult_21_C245_n737, mult_21_C245_n736, 
      mult_21_C245_n735, mult_21_C245_n734, mult_21_C245_n733, 
      mult_21_C245_n732, mult_21_C245_n731, mult_21_C245_n730, 
      mult_21_C245_n729, mult_21_C245_n728, mult_21_C245_n727, 
      mult_21_C245_n726, mult_21_C245_n725, mult_21_C245_n724, 
      mult_21_C245_n723, mult_21_C245_n722, mult_21_C245_n721, 
      mult_21_C245_n720, mult_21_C245_n719, mult_21_C245_n718, 
      mult_21_C245_n717, mult_21_C245_n716, mult_21_C245_n715, 
      mult_21_C245_n714, mult_21_C245_n713, mult_21_C245_n712, 
      mult_21_C245_n711, mult_21_C245_n710, mult_21_C245_n709, 
      mult_21_C245_n708, mult_21_C245_n707, mult_21_C245_n706, 
      mult_21_C245_n705, mult_21_C245_n704, mult_21_C245_n703, 
      mult_21_C245_n702, mult_21_C245_n701, mult_21_C245_n700, 
      mult_21_C245_n699, mult_21_C245_n698, mult_21_C245_n697, 
      mult_21_C245_n696, mult_21_C245_n695, mult_21_C245_n694, 
      mult_21_C245_n693, mult_21_C245_n692, mult_21_C245_n691, 
      mult_21_C245_n690, mult_21_C245_n689, mult_21_C245_n688, 
      mult_21_C245_n687, mult_21_C245_n686, mult_21_C245_n685, 
      mult_21_C245_n684, mult_21_C245_n683, mult_21_C245_n682, 
      mult_21_C245_n681, mult_21_C245_n680, mult_21_C245_n679, 
      mult_21_C245_n678, mult_21_C245_n677, mult_21_C245_n676, 
      mult_21_C245_n675, mult_21_C245_n674, mult_21_C245_n673, 
      mult_21_C245_n672, mult_21_C245_n671, mult_21_C245_n670, 
      mult_21_C245_n669, mult_21_C245_n668, mult_21_C245_n667, 
      mult_21_C245_n666, mult_21_C245_n665, mult_21_C245_n664, 
      mult_21_C245_n663, mult_21_C245_n662, mult_21_C245_n661, 
      mult_21_C245_n660, mult_21_C245_n659, mult_21_C245_n658, 
      mult_21_C245_n657, mult_21_C245_n656, mult_21_C245_n655, 
      mult_21_C245_n654, mult_21_C245_n653, mult_21_C245_n652, 
      mult_21_C245_n651, mult_21_C245_n650, mult_21_C245_n649, 
      mult_21_C245_n648, mult_21_C245_n647, mult_21_C245_n646, 
      mult_21_C245_n645, mult_21_C245_n644, mult_21_C245_n643, 
      mult_21_C245_n642, mult_21_C245_n641, mult_21_C245_n640, 
      mult_21_C245_n639, mult_21_C245_n638, mult_21_C245_n637, 
      mult_21_C245_n636, mult_21_C245_n635, mult_21_C245_n634, 
      mult_21_C245_n633, mult_21_C245_n632, mult_21_C245_n631, 
      mult_21_C245_n630, mult_21_C245_n629, mult_21_C245_n628, 
      mult_21_C245_n627, mult_21_C245_n626, mult_21_C245_n625, 
      mult_21_C245_n624, mult_21_C245_n623, mult_21_C245_n622, 
      mult_21_C245_n621, mult_21_C245_n620, mult_21_C245_n619, 
      mult_21_C245_n618, mult_21_C245_n617, mult_21_C245_n616, 
      mult_21_C245_n615, mult_21_C245_n614, mult_21_C245_n613, 
      mult_21_C245_n612, mult_21_C245_n611, mult_21_C245_n610, 
      mult_21_C245_n609, mult_21_C245_n608, mult_21_C245_n607, 
      mult_21_C245_n606, mult_21_C245_n605, mult_21_C245_n604, 
      mult_21_C245_n603, mult_21_C245_n602, mult_21_C245_n601, 
      mult_21_C245_n600, mult_21_C245_n599, mult_21_C245_n598, 
      mult_21_C245_n597, mult_21_C245_n596, mult_21_C245_n595, 
      mult_21_C245_n594, mult_21_C245_n593, mult_21_C245_n592, 
      mult_21_C245_n591, mult_21_C245_n590, mult_21_C245_n589, 
      mult_21_C245_n588, mult_21_C245_n587, mult_21_C245_n586, 
      mult_21_C245_n585, mult_21_C245_n584, mult_21_C245_n583, 
      mult_21_C245_n582, mult_21_C245_n581, mult_21_C245_n580, 
      mult_21_C245_n579, mult_21_C245_n578, mult_21_C245_n577, 
      mult_21_C245_n576, mult_21_C245_n575, mult_21_C245_n574, 
      mult_21_C245_n573, mult_21_C245_n572, mult_21_C245_n571, 
      mult_21_C245_n570, mult_21_C245_n569, mult_21_C245_n568, 
      mult_21_C245_n567, mult_21_C245_n566, mult_21_C245_n565, 
      mult_21_C245_n564, mult_21_C245_n563, mult_21_C245_n562, 
      mult_21_C245_n561, mult_21_C245_n560, mult_21_C245_n559, 
      mult_21_C245_n558, mult_21_C245_n557, mult_21_C245_n556, 
      mult_21_C245_n555, mult_21_C245_n554, mult_21_C245_n553, 
      mult_21_C245_n552, mult_21_C245_n551, mult_21_C245_n550, 
      mult_21_C245_n549, mult_21_C245_n548, mult_21_C245_n547, 
      mult_21_C245_n546, mult_21_C245_n545, mult_21_C245_n544, 
      mult_21_C245_n543, mult_21_C245_n542, mult_21_C245_n541, 
      mult_21_C245_n540, mult_21_C245_n539, mult_21_C245_n538, 
      mult_21_C245_n537, mult_21_C245_n536, mult_21_C245_n535, 
      mult_21_C245_n534, mult_21_C245_n533, mult_21_C245_n532, 
      mult_21_C245_n531, mult_21_C245_n530, mult_21_C245_n529, 
      mult_21_C245_n528, mult_21_C245_n527, mult_21_C245_n526, 
      mult_21_C245_n525, mult_21_C245_n524, mult_21_C245_n523, 
      mult_21_C245_n522, mult_21_C245_n521, mult_21_C245_n520, 
      mult_21_C245_n519, mult_21_C245_n518, mult_21_C245_n517, 
      mult_21_C245_n516, mult_21_C245_n515, mult_21_C245_n514, 
      mult_21_C245_n513, mult_21_C245_n512, mult_21_C245_n511, 
      mult_21_C245_n510, mult_21_C245_n509, mult_21_C245_n508, 
      mult_21_C245_n507, mult_21_C245_n506, mult_21_C245_n505, 
      mult_21_C245_n504, mult_21_C245_n503, mult_21_C245_n502, 
      mult_21_C245_n501, mult_21_C245_n500, mult_21_C245_n499, 
      mult_21_C245_n498, mult_21_C245_n497, mult_21_C245_n496, 
      mult_21_C245_n495, mult_21_C245_n494, mult_21_C245_n493, 
      mult_21_C245_n492, mult_21_C245_n491, mult_21_C245_n490, 
      mult_21_C245_n489, mult_21_C245_n488, mult_21_C245_n487, 
      mult_21_C245_n486, mult_21_C245_n485, mult_21_C245_n484, 
      mult_21_C245_n483, mult_21_C245_n482, mult_21_C245_n481, 
      mult_21_C245_n480, mult_21_C245_n479, mult_21_C245_n478, 
      mult_21_C245_n477, mult_21_C245_n476, mult_21_C245_n475, 
      mult_21_C245_n474, mult_21_C245_n473, mult_21_C245_n472, 
      mult_21_C245_n471, mult_21_C245_n470, mult_21_C245_n469, 
      mult_21_C245_n468, mult_21_C245_n467, mult_21_C245_n466, 
      mult_21_C245_n465, mult_21_C245_n464, mult_21_C245_n463, 
      mult_21_C245_n462, mult_21_C245_n461, mult_21_C245_n460, 
      mult_21_C245_n459, mult_21_C245_n458, mult_21_C245_n457, 
      mult_21_C245_n456, mult_21_C245_n455, mult_21_C245_n454, 
      mult_21_C245_n453, mult_21_C245_n452, mult_21_C245_n451, 
      mult_21_C245_n450, mult_21_C245_n449, mult_21_C245_n448, 
      mult_21_C245_n447, mult_21_C245_n446, mult_21_C245_n445, 
      mult_21_C245_n444, mult_21_C245_n443, mult_21_C245_n442, 
      mult_21_C245_n441, mult_21_C245_n440, mult_21_C245_n439, 
      mult_21_C245_n438, mult_21_C245_n437, mult_21_C245_n436, 
      mult_21_C245_n435, mult_21_C245_n434, mult_21_C245_n433, 
      mult_21_C245_n432, mult_21_C245_n431, mult_21_C245_n430, 
      mult_21_C245_n429, mult_21_C245_n428, mult_21_C245_n427, 
      mult_21_C245_n426, mult_21_C245_n425, mult_21_C245_n424, 
      mult_21_C245_n423, mult_21_C245_n422, mult_21_C245_n421, 
      mult_21_C245_n420, mult_21_C245_n419, mult_21_C245_n418, 
      mult_21_C245_n417, mult_21_C245_n416, mult_21_C245_n415, 
      mult_21_C245_n414, mult_21_C245_n413, mult_21_C245_n412, 
      mult_21_C245_n411, mult_21_C245_n410, mult_21_C245_n409, 
      mult_21_C245_n408, mult_21_C245_n407, mult_21_C245_n406, 
      mult_21_C245_n405, mult_21_C245_n404, mult_21_C245_n403, 
      mult_21_C245_n402, mult_21_C245_n401, mult_21_C245_n400, 
      mult_21_C245_n399, mult_21_C245_n398, mult_21_C245_n397, 
      mult_21_C245_n396, mult_21_C245_n395, mult_21_C245_n394, 
      mult_21_C245_n393, mult_21_C245_n392, mult_21_C245_n391, 
      mult_21_C245_n390, mult_21_C245_n389, mult_21_C245_n388, 
      mult_21_C245_n387, mult_21_C245_n386, mult_21_C245_n385, 
      mult_21_C245_n384, mult_21_C245_n383, mult_21_C245_n382, 
      mult_21_C245_n381, mult_21_C245_n380, mult_21_C245_n379, 
      mult_21_C245_n378, mult_21_C245_n377, mult_21_C245_n376, 
      mult_21_C245_n375, mult_21_C245_n374, mult_21_C245_n373, 
      mult_21_C245_n372, mult_21_C245_n371, mult_21_C245_n370, 
      mult_21_C245_n369, mult_21_C245_n368, mult_21_C245_n367, 
      mult_21_C245_n366, mult_21_C245_n365, mult_21_C245_n364, 
      mult_21_C245_n363, mult_21_C245_n362, mult_21_C245_n361, 
      mult_21_C245_n360, mult_21_C245_n359, mult_21_C245_n358, 
      mult_21_C245_n357, mult_21_C245_n356, mult_21_C245_n355, 
      mult_21_C245_n354, mult_21_C245_n353, mult_21_C245_n352, 
      mult_21_C245_n351, mult_21_C245_n350, mult_21_C245_n349, 
      mult_21_C245_n348, mult_21_C245_n347, mult_21_C245_n346, 
      mult_21_C245_n345, mult_21_C245_n344, mult_21_C245_n343, 
      mult_21_C245_n342, mult_21_C245_n341, mult_21_C245_n340, 
      mult_21_C245_n339, mult_21_C245_n338, mult_21_C245_n337, 
      mult_21_C245_n336, mult_21_C245_n335, mult_21_C245_n334, 
      mult_21_C245_n333, mult_21_C245_n332, mult_21_C245_n331, 
      mult_21_C245_n330, mult_21_C245_n329, mult_21_C245_n328, 
      mult_21_C245_n327, mult_21_C245_n326, mult_21_C245_n325, 
      mult_21_C245_n324, mult_21_C245_n323, mult_21_C245_n322, 
      mult_21_C245_n321, mult_21_C245_n320, mult_21_C245_n319, 
      mult_21_C245_n318, mult_21_C245_n317, mult_21_C245_n316, 
      mult_21_C245_n315, mult_21_C245_n314, mult_21_C245_n313, 
      mult_21_C245_n312, mult_21_C245_n311, mult_21_C245_n310, 
      mult_21_C245_n309, mult_21_C245_n308, mult_21_C245_n307, 
      mult_21_C245_n306, mult_21_C245_n305, mult_21_C245_n304, 
      mult_21_C245_n303, mult_21_C245_n302, mult_21_C245_n301, 
      mult_21_C245_n300, mult_21_C245_n299, mult_21_C245_n298, 
      mult_21_C245_n297, mult_21_C245_n296, mult_21_C245_n295, 
      mult_21_C245_n294, mult_21_C245_n293, mult_21_C245_n292, 
      mult_21_C245_n291, mult_21_C245_n290, mult_21_C245_n289, 
      mult_21_C245_n288, mult_21_C245_n287, mult_21_C245_n286, 
      mult_21_C245_n285, mult_21_C245_n284, mult_21_C245_n283, 
      mult_21_C245_n282, mult_21_C245_n281, mult_21_C245_n280, 
      mult_21_C245_n279, mult_21_C245_n278, mult_21_C245_n277, 
      mult_21_C245_n276, mult_21_C245_n275, mult_21_C245_n274, 
      mult_21_C245_n273, mult_21_C245_n272, mult_21_C245_n271, 
      mult_21_C245_n270, mult_21_C245_n269, mult_21_C245_n268, 
      mult_21_C245_n267, mult_21_C245_n266, mult_21_C245_n265, 
      mult_21_C245_n264, mult_21_C245_n263, mult_21_C245_n262, 
      mult_21_C245_n261, mult_21_C245_n260, mult_21_C245_n259, 
      mult_21_C245_n258, mult_21_C245_n257, mult_21_C245_n256, 
      mult_21_C245_n255, mult_21_C245_n254, mult_21_C245_n253, 
      mult_21_C245_n252, mult_21_C245_n251, mult_21_C245_n250, 
      mult_21_C245_n249, mult_21_C245_n248, mult_21_C245_n247, 
      mult_21_C245_n246, mult_21_C245_n245, mult_21_C245_n244, 
      mult_21_C245_n243, mult_21_C245_n242, mult_21_C245_n241, 
      mult_21_C245_n240, mult_21_C245_n239, mult_21_C245_n238, 
      mult_21_C245_n237, mult_21_C245_n236, mult_21_C245_n235, 
      mult_21_C245_n234, mult_21_C245_n233, mult_21_C245_n232, 
      mult_21_C245_n231, mult_21_C245_n230, mult_21_C245_n229, 
      mult_21_C245_n228, mult_21_C245_n227, mult_21_C245_n226, 
      mult_21_C245_n225, mult_21_C245_n224, mult_21_C245_n223, 
      mult_21_C245_n222, mult_21_C245_n221, mult_21_C245_n220, 
      mult_21_C245_n219, mult_21_C245_n218, mult_21_C245_n217, 
      mult_21_C245_n216, mult_21_C245_n215, mult_21_C245_n214, 
      mult_21_C245_n213, mult_21_C245_n212, mult_21_C245_n211, 
      mult_21_C245_n210, mult_21_C245_n209, mult_21_C245_n208, 
      mult_21_C245_n207, mult_21_C245_n206, mult_21_C245_n205, 
      mult_21_C245_n204, mult_21_C245_n203, mult_21_C245_n202, 
      mult_21_C245_n186, mult_21_C245_n185, mult_21_C245_n184, 
      mult_21_C245_n183, mult_21_C245_n182, mult_21_C245_n181, 
      mult_21_C245_n180, mult_21_C245_n179, mult_21_C245_n178, 
      mult_21_C245_n177, mult_21_C245_n176, mult_21_C245_n175, 
      mult_21_C245_n174, mult_21_C245_n173, mult_21_C245_n172, 
      mult_21_C245_n171, mult_21_C245_n170, mult_21_C245_n169, 
      mult_21_C245_n168, mult_21_C245_n167, mult_21_C245_n166, 
      mult_21_C245_n165, mult_21_C245_n164, mult_21_C245_n163, 
      mult_21_C245_n162, mult_21_C245_n161, mult_21_C245_n160, 
      mult_21_C245_n159, mult_21_C245_n158, mult_21_C245_n157, 
      mult_21_C245_n156, mult_21_C245_n104, mult_21_C245_n99, mult_21_C245_n94,
      mult_21_C245_n89, mult_21_C245_n84, mult_21_C245_n80, mult_21_C245_n73, 
      mult_21_C245_n66, mult_21_C245_n58, mult_21_C245_n50, mult_21_C245_n42, 
      mult_21_C247_n1457, mult_21_C247_n1456, mult_21_C247_n1455, 
      mult_21_C247_n1454, mult_21_C247_n1453, mult_21_C247_n1452, 
      mult_21_C247_n1451, mult_21_C247_n1450, mult_21_C247_n1449, 
      mult_21_C247_n1448, mult_21_C247_n1447, mult_21_C247_n1446, 
      mult_21_C247_n1445, mult_21_C247_n1444, mult_21_C247_n1443, 
      mult_21_C247_n1442, mult_21_C247_n1441, mult_21_C247_n1440, 
      mult_21_C247_n1439, mult_21_C247_n1438, mult_21_C247_n1437, 
      mult_21_C247_n1436, mult_21_C247_n1435, mult_21_C247_n1434, 
      mult_21_C247_n1433, mult_21_C247_n1432, mult_21_C247_n1431, 
      mult_21_C247_n1430, mult_21_C247_n1429, mult_21_C247_n1428, 
      mult_21_C247_n1427, mult_21_C247_n1426, mult_21_C247_n1425, 
      mult_21_C247_n1424, mult_21_C247_n1423, mult_21_C247_n1422, 
      mult_21_C247_n1421, mult_21_C247_n1420, mult_21_C247_n1419, 
      mult_21_C247_n1418, mult_21_C247_n1417, mult_21_C247_n1416, 
      mult_21_C247_n1415, mult_21_C247_n1414, mult_21_C247_n1413, 
      mult_21_C247_n1412, mult_21_C247_n1411, mult_21_C247_n1410, 
      mult_21_C247_n1409, mult_21_C247_n1408, mult_21_C247_n1407, 
      mult_21_C247_n1406, mult_21_C247_n1405, mult_21_C247_n1404, 
      mult_21_C247_n1403, mult_21_C247_n1402, mult_21_C247_n1401, 
      mult_21_C247_n1400, mult_21_C247_n1399, mult_21_C247_n1398, 
      mult_21_C247_n1397, mult_21_C247_n1396, mult_21_C247_n1395, 
      mult_21_C247_n1394, mult_21_C247_n1393, mult_21_C247_n1392, 
      mult_21_C247_n1391, mult_21_C247_n1390, mult_21_C247_n1389, 
      mult_21_C247_n1388, mult_21_C247_n1387, mult_21_C247_n1386, 
      mult_21_C247_n1385, mult_21_C247_n1384, mult_21_C247_n1383, 
      mult_21_C247_n1382, mult_21_C247_n1381, mult_21_C247_n1380, 
      mult_21_C247_n1379, mult_21_C247_n1378, mult_21_C247_n1377, 
      mult_21_C247_n1376, mult_21_C247_n1375, mult_21_C247_n1226, 
      mult_21_C247_n1225, mult_21_C247_n1224, mult_21_C247_n1223, 
      mult_21_C247_n1222, mult_21_C247_n1221, mult_21_C247_n1220, 
      mult_21_C247_n1219, mult_21_C247_n1218, mult_21_C247_n1217, 
      mult_21_C247_n1216, mult_21_C247_n1215, mult_21_C247_n1214, 
      mult_21_C247_n1213, mult_21_C247_n1212, mult_21_C247_n1211, 
      mult_21_C247_n1210, mult_21_C247_n1209, mult_21_C247_n1208, 
      mult_21_C247_n1207, mult_21_C247_n1206, mult_21_C247_n1205, 
      mult_21_C247_n1204, mult_21_C247_n1203, mult_21_C247_n1202, 
      mult_21_C247_n1201, mult_21_C247_n1200, mult_21_C247_n1199, 
      mult_21_C247_n1198, mult_21_C247_n1197, mult_21_C247_n1196, 
      mult_21_C247_n1195, mult_21_C247_n1194, mult_21_C247_n1193, 
      mult_21_C247_n1192, mult_21_C247_n1191, mult_21_C247_n1190, 
      mult_21_C247_n1189, mult_21_C247_n1188, mult_21_C247_n1187, 
      mult_21_C247_n1186, mult_21_C247_n1185, mult_21_C247_n1184, 
      mult_21_C247_n1183, mult_21_C247_n1182, mult_21_C247_n1181, 
      mult_21_C247_n1180, mult_21_C247_n1179, mult_21_C247_n1178, 
      mult_21_C247_n1177, mult_21_C247_n1176, mult_21_C247_n1175, 
      mult_21_C247_n1174, mult_21_C247_n1173, mult_21_C247_n1172, 
      mult_21_C247_n1171, mult_21_C247_n1170, mult_21_C247_n1169, 
      mult_21_C247_n1168, mult_21_C247_n1167, mult_21_C247_n1166, 
      mult_21_C247_n1165, mult_21_C247_n1164, mult_21_C247_n1163, 
      mult_21_C247_n1162, mult_21_C247_n1161, mult_21_C247_n1160, 
      mult_21_C247_n1159, mult_21_C247_n1158, mult_21_C247_n1157, 
      mult_21_C247_n1156, mult_21_C247_n1155, mult_21_C247_n1154, 
      mult_21_C247_n1153, mult_21_C247_n1152, mult_21_C247_n1151, 
      mult_21_C247_n1150, mult_21_C247_n1149, mult_21_C247_n1148, 
      mult_21_C247_n1147, mult_21_C247_n1146, mult_21_C247_n1145, 
      mult_21_C247_n1144, mult_21_C247_n1143, mult_21_C247_n1142, 
      mult_21_C247_n1141, mult_21_C247_n1140, mult_21_C247_n1139, 
      mult_21_C247_n1138, mult_21_C247_n1137, mult_21_C247_n1136, 
      mult_21_C247_n1135, mult_21_C247_n1134, mult_21_C247_n1133, 
      mult_21_C247_n1132, mult_21_C247_n1131, mult_21_C247_n1130, 
      mult_21_C247_n1129, mult_21_C247_n1128, mult_21_C247_n1127, 
      mult_21_C247_n1126, mult_21_C247_n1125, mult_21_C247_n1124, 
      mult_21_C247_n1123, mult_21_C247_n1122, mult_21_C247_n1121, 
      mult_21_C247_n1120, mult_21_C247_n1119, mult_21_C247_n1118, 
      mult_21_C247_n1117, mult_21_C247_n1116, mult_21_C247_n1115, 
      mult_21_C247_n1114, mult_21_C247_n1113, mult_21_C247_n1112, 
      mult_21_C247_n1111, mult_21_C247_n1110, mult_21_C247_n1109, 
      mult_21_C247_n1108, mult_21_C247_n1107, mult_21_C247_n1106, 
      mult_21_C247_n1105, mult_21_C247_n1104, mult_21_C247_n1103, 
      mult_21_C247_n1102, mult_21_C247_n1101, mult_21_C247_n1100, 
      mult_21_C247_n1099, mult_21_C247_n1098, mult_21_C247_n1097, 
      mult_21_C247_n1096, mult_21_C247_n1095, mult_21_C247_n1094, 
      mult_21_C247_n1093, mult_21_C247_n1092, mult_21_C247_n1091, 
      mult_21_C247_n1090, mult_21_C247_n1089, mult_21_C247_n1088, 
      mult_21_C247_n1087, mult_21_C247_n1086, mult_21_C247_n1085, 
      mult_21_C247_n1084, mult_21_C247_n1083, mult_21_C247_n1082, 
      mult_21_C247_n1081, mult_21_C247_n1080, mult_21_C247_n1079, 
      mult_21_C247_n1078, mult_21_C247_n1077, mult_21_C247_n1076, 
      mult_21_C247_n1075, mult_21_C247_n1074, mult_21_C247_n1073, 
      mult_21_C247_n1072, mult_21_C247_n1071, mult_21_C247_n1070, 
      mult_21_C247_n1069, mult_21_C247_n1068, mult_21_C247_n1067, 
      mult_21_C247_n1066, mult_21_C247_n1065, mult_21_C247_n1064, 
      mult_21_C247_n1063, mult_21_C247_n1062, mult_21_C247_n1061, 
      mult_21_C247_n1060, mult_21_C247_n1059, mult_21_C247_n1058, 
      mult_21_C247_n1057, mult_21_C247_n1056, mult_21_C247_n1055, 
      mult_21_C247_n1054, mult_21_C247_n1053, mult_21_C247_n1052, 
      mult_21_C247_n1051, mult_21_C247_n1050, mult_21_C247_n1049, 
      mult_21_C247_n1048, mult_21_C247_n1047, mult_21_C247_n1046, 
      mult_21_C247_n1045, mult_21_C247_n1044, mult_21_C247_n1043, 
      mult_21_C247_n1042, mult_21_C247_n1041, mult_21_C247_n1040, 
      mult_21_C247_n1039, mult_21_C247_n1038, mult_21_C247_n1037, 
      mult_21_C247_n1036, mult_21_C247_n1035, mult_21_C247_n1034, 
      mult_21_C247_n1033, mult_21_C247_n1032, mult_21_C247_n1031, 
      mult_21_C247_n1030, mult_21_C247_n1029, mult_21_C247_n1028, 
      mult_21_C247_n1027, mult_21_C247_n1026, mult_21_C247_n1025, 
      mult_21_C247_n1024, mult_21_C247_n1023, mult_21_C247_n1022, 
      mult_21_C247_n1021, mult_21_C247_n1020, mult_21_C247_n1019, 
      mult_21_C247_n1018, mult_21_C247_n1017, mult_21_C247_n1016, 
      mult_21_C247_n1015, mult_21_C247_n1014, mult_21_C247_n1013, 
      mult_21_C247_n1012, mult_21_C247_n1011, mult_21_C247_n1010, 
      mult_21_C247_n1009, mult_21_C247_n1008, mult_21_C247_n1007, 
      mult_21_C247_n1006, mult_21_C247_n1005, mult_21_C247_n1004, 
      mult_21_C247_n1003, mult_21_C247_n1002, mult_21_C247_n1001, 
      mult_21_C247_n1000, mult_21_C247_n999, mult_21_C247_n998, 
      mult_21_C247_n997, mult_21_C247_n996, mult_21_C247_n995, 
      mult_21_C247_n994, mult_21_C247_n993, mult_21_C247_n992, 
      mult_21_C247_n991, mult_21_C247_n990, mult_21_C247_n989, 
      mult_21_C247_n988, mult_21_C247_n987, mult_21_C247_n986, 
      mult_21_C247_n985, mult_21_C247_n984, mult_21_C247_n983, 
      mult_21_C247_n982, mult_21_C247_n981, mult_21_C247_n980, 
      mult_21_C247_n979, mult_21_C247_n978, mult_21_C247_n977, 
      mult_21_C247_n976, mult_21_C247_n975, mult_21_C247_n974, 
      mult_21_C247_n973, mult_21_C247_n972, mult_21_C247_n971, 
      mult_21_C247_n970, mult_21_C247_n969, mult_21_C247_n968, 
      mult_21_C247_n967, mult_21_C247_n966, mult_21_C247_n965, 
      mult_21_C247_n964, mult_21_C247_n963, mult_21_C247_n962, 
      mult_21_C247_n961, mult_21_C247_n960, mult_21_C247_n959, 
      mult_21_C247_n958, mult_21_C247_n957, mult_21_C247_n956, 
      mult_21_C247_n955, mult_21_C247_n953, mult_21_C247_n952, 
      mult_21_C247_n951, mult_21_C247_n950, mult_21_C247_n949, 
      mult_21_C247_n948, mult_21_C247_n947, mult_21_C247_n946, 
      mult_21_C247_n945, mult_21_C247_n944, mult_21_C247_n943, 
      mult_21_C247_n942, mult_21_C247_n941, mult_21_C247_n940, 
      mult_21_C247_n939, mult_21_C247_n923, mult_21_C247_n922, 
      mult_21_C247_n921, mult_21_C247_n920, mult_21_C247_n919, 
      mult_21_C247_n918, mult_21_C247_n917, mult_21_C247_n916, 
      mult_21_C247_n915, mult_21_C247_n914, mult_21_C247_n913, 
      mult_21_C247_n912, mult_21_C247_n911, mult_21_C247_n910, 
      mult_21_C247_n909, mult_21_C247_n908, mult_21_C247_n907, 
      mult_21_C247_n906, mult_21_C247_n905, mult_21_C247_n904, 
      mult_21_C247_n903, mult_21_C247_n902, mult_21_C247_n901, 
      mult_21_C247_n900, mult_21_C247_n899, mult_21_C247_n898, 
      mult_21_C247_n897, mult_21_C247_n896, mult_21_C247_n895, 
      mult_21_C247_n894, mult_21_C247_n893, mult_21_C247_n892, 
      mult_21_C247_n891, mult_21_C247_n890, mult_21_C247_n889, 
      mult_21_C247_n888, mult_21_C247_n887, mult_21_C247_n886, 
      mult_21_C247_n885, mult_21_C247_n884, mult_21_C247_n883, 
      mult_21_C247_n882, mult_21_C247_n881, mult_21_C247_n880, 
      mult_21_C247_n879, mult_21_C247_n878, mult_21_C247_n877, 
      mult_21_C247_n876, mult_21_C247_n875, mult_21_C247_n874, 
      mult_21_C247_n873, mult_21_C247_n872, mult_21_C247_n871, 
      mult_21_C247_n870, mult_21_C247_n869, mult_21_C247_n868, 
      mult_21_C247_n867, mult_21_C247_n866, mult_21_C247_n865, 
      mult_21_C247_n864, mult_21_C247_n863, mult_21_C247_n862, 
      mult_21_C247_n861, mult_21_C247_n860, mult_21_C247_n859, 
      mult_21_C247_n858, mult_21_C247_n857, mult_21_C247_n856, 
      mult_21_C247_n855, mult_21_C247_n854, mult_21_C247_n853, 
      mult_21_C247_n852, mult_21_C247_n851, mult_21_C247_n850, 
      mult_21_C247_n849, mult_21_C247_n848, mult_21_C247_n847, 
      mult_21_C247_n846, mult_21_C247_n845, mult_21_C247_n844, 
      mult_21_C247_n843, mult_21_C247_n842, mult_21_C247_n841, 
      mult_21_C247_n840, mult_21_C247_n839, mult_21_C247_n838, 
      mult_21_C247_n837, mult_21_C247_n836, mult_21_C247_n835, 
      mult_21_C247_n834, mult_21_C247_n833, mult_21_C247_n832, 
      mult_21_C247_n831, mult_21_C247_n830, mult_21_C247_n829, 
      mult_21_C247_n828, mult_21_C247_n827, mult_21_C247_n826, 
      mult_21_C247_n825, mult_21_C247_n824, mult_21_C247_n823, 
      mult_21_C247_n822, mult_21_C247_n821, mult_21_C247_n820, 
      mult_21_C247_n819, mult_21_C247_n818, mult_21_C247_n817, 
      mult_21_C247_n816, mult_21_C247_n815, mult_21_C247_n814, 
      mult_21_C247_n813, mult_21_C247_n812, mult_21_C247_n811, 
      mult_21_C247_n810, mult_21_C247_n809, mult_21_C247_n808, 
      mult_21_C247_n807, mult_21_C247_n806, mult_21_C247_n805, 
      mult_21_C247_n804, mult_21_C247_n803, mult_21_C247_n802, 
      mult_21_C247_n801, mult_21_C247_n800, mult_21_C247_n799, 
      mult_21_C247_n798, mult_21_C247_n797, mult_21_C247_n796, 
      mult_21_C247_n795, mult_21_C247_n794, mult_21_C247_n793, 
      mult_21_C247_n792, mult_21_C247_n791, mult_21_C247_n790, 
      mult_21_C247_n789, mult_21_C247_n788, mult_21_C247_n787, 
      mult_21_C247_n786, mult_21_C247_n785, mult_21_C247_n784, 
      mult_21_C247_n783, mult_21_C247_n782, mult_21_C247_n781, 
      mult_21_C247_n780, mult_21_C247_n779, mult_21_C247_n778, 
      mult_21_C247_n777, mult_21_C247_n776, mult_21_C247_n775, 
      mult_21_C247_n774, mult_21_C247_n773, mult_21_C247_n772, 
      mult_21_C247_n771, mult_21_C247_n770, mult_21_C247_n769, 
      mult_21_C247_n768, mult_21_C247_n767, mult_21_C247_n766, 
      mult_21_C247_n765, mult_21_C247_n764, mult_21_C247_n763, 
      mult_21_C247_n762, mult_21_C247_n761, mult_21_C247_n760, 
      mult_21_C247_n759, mult_21_C247_n758, mult_21_C247_n757, 
      mult_21_C247_n756, mult_21_C247_n755, mult_21_C247_n754, 
      mult_21_C247_n753, mult_21_C247_n752, mult_21_C247_n751, 
      mult_21_C247_n750, mult_21_C247_n749, mult_21_C247_n748, 
      mult_21_C247_n747, mult_21_C247_n746, mult_21_C247_n745, 
      mult_21_C247_n744, mult_21_C247_n743, mult_21_C247_n742, 
      mult_21_C247_n741, mult_21_C247_n740, mult_21_C247_n739, 
      mult_21_C247_n738, mult_21_C247_n737, mult_21_C247_n736, 
      mult_21_C247_n735, mult_21_C247_n734, mult_21_C247_n733, 
      mult_21_C247_n732, mult_21_C247_n731, mult_21_C247_n730, 
      mult_21_C247_n729, mult_21_C247_n728, mult_21_C247_n727, 
      mult_21_C247_n726, mult_21_C247_n725, mult_21_C247_n724, 
      mult_21_C247_n723, mult_21_C247_n722, mult_21_C247_n721, 
      mult_21_C247_n720, mult_21_C247_n719, mult_21_C247_n718, 
      mult_21_C247_n717, mult_21_C247_n716, mult_21_C247_n715, 
      mult_21_C247_n714, mult_21_C247_n713, mult_21_C247_n712, 
      mult_21_C247_n711, mult_21_C247_n710, mult_21_C247_n709, 
      mult_21_C247_n708, mult_21_C247_n707, mult_21_C247_n706, 
      mult_21_C247_n705, mult_21_C247_n704, mult_21_C247_n703, 
      mult_21_C247_n702, mult_21_C247_n701, mult_21_C247_n700, 
      mult_21_C247_n699, mult_21_C247_n698, mult_21_C247_n697, 
      mult_21_C247_n696, mult_21_C247_n695, mult_21_C247_n694, 
      mult_21_C247_n693, mult_21_C247_n692, mult_21_C247_n691, 
      mult_21_C247_n690, mult_21_C247_n689, mult_21_C247_n688, 
      mult_21_C247_n687, mult_21_C247_n686, mult_21_C247_n685, 
      mult_21_C247_n684, mult_21_C247_n683, mult_21_C247_n682, 
      mult_21_C247_n681, mult_21_C247_n680, mult_21_C247_n679, 
      mult_21_C247_n678, mult_21_C247_n677, mult_21_C247_n676, 
      mult_21_C247_n675, mult_21_C247_n674, mult_21_C247_n673, 
      mult_21_C247_n672, mult_21_C247_n671, mult_21_C247_n670, 
      mult_21_C247_n669, mult_21_C247_n668, mult_21_C247_n667, 
      mult_21_C247_n666, mult_21_C247_n665, mult_21_C247_n664, 
      mult_21_C247_n663, mult_21_C247_n662, mult_21_C247_n661, 
      mult_21_C247_n660, mult_21_C247_n659, mult_21_C247_n658, 
      mult_21_C247_n657, mult_21_C247_n656, mult_21_C247_n655, 
      mult_21_C247_n654, mult_21_C247_n653, mult_21_C247_n652, 
      mult_21_C247_n651, mult_21_C247_n650, mult_21_C247_n649, 
      mult_21_C247_n648, mult_21_C247_n647, mult_21_C247_n646, 
      mult_21_C247_n645, mult_21_C247_n644, mult_21_C247_n643, 
      mult_21_C247_n642, mult_21_C247_n641, mult_21_C247_n640, 
      mult_21_C247_n639, mult_21_C247_n638, mult_21_C247_n637, 
      mult_21_C247_n636, mult_21_C247_n635, mult_21_C247_n634, 
      mult_21_C247_n633, mult_21_C247_n632, mult_21_C247_n631, 
      mult_21_C247_n630, mult_21_C247_n629, mult_21_C247_n628, 
      mult_21_C247_n627, mult_21_C247_n626, mult_21_C247_n625, 
      mult_21_C247_n624, mult_21_C247_n623, mult_21_C247_n622, 
      mult_21_C247_n621, mult_21_C247_n620, mult_21_C247_n619, 
      mult_21_C247_n618, mult_21_C247_n617, mult_21_C247_n616, 
      mult_21_C247_n615, mult_21_C247_n614, mult_21_C247_n613, 
      mult_21_C247_n612, mult_21_C247_n611, mult_21_C247_n610, 
      mult_21_C247_n609, mult_21_C247_n608, mult_21_C247_n607, 
      mult_21_C247_n606, mult_21_C247_n605, mult_21_C247_n604, 
      mult_21_C247_n603, mult_21_C247_n602, mult_21_C247_n601, 
      mult_21_C247_n600, mult_21_C247_n599, mult_21_C247_n598, 
      mult_21_C247_n597, mult_21_C247_n596, mult_21_C247_n595, 
      mult_21_C247_n594, mult_21_C247_n593, mult_21_C247_n592, 
      mult_21_C247_n591, mult_21_C247_n590, mult_21_C247_n589, 
      mult_21_C247_n588, mult_21_C247_n587, mult_21_C247_n586, 
      mult_21_C247_n585, mult_21_C247_n584, mult_21_C247_n583, 
      mult_21_C247_n582, mult_21_C247_n581, mult_21_C247_n580, 
      mult_21_C247_n579, mult_21_C247_n578, mult_21_C247_n577, 
      mult_21_C247_n576, mult_21_C247_n575, mult_21_C247_n574, 
      mult_21_C247_n573, mult_21_C247_n572, mult_21_C247_n571, 
      mult_21_C247_n570, mult_21_C247_n569, mult_21_C247_n568, 
      mult_21_C247_n567, mult_21_C247_n566, mult_21_C247_n565, 
      mult_21_C247_n564, mult_21_C247_n563, mult_21_C247_n562, 
      mult_21_C247_n561, mult_21_C247_n560, mult_21_C247_n559, 
      mult_21_C247_n558, mult_21_C247_n557, mult_21_C247_n556, 
      mult_21_C247_n555, mult_21_C247_n554, mult_21_C247_n553, 
      mult_21_C247_n552, mult_21_C247_n551, mult_21_C247_n550, 
      mult_21_C247_n549, mult_21_C247_n548, mult_21_C247_n547, 
      mult_21_C247_n546, mult_21_C247_n545, mult_21_C247_n544, 
      mult_21_C247_n543, mult_21_C247_n542, mult_21_C247_n541, 
      mult_21_C247_n540, mult_21_C247_n539, mult_21_C247_n538, 
      mult_21_C247_n537, mult_21_C247_n536, mult_21_C247_n535, 
      mult_21_C247_n534, mult_21_C247_n533, mult_21_C247_n532, 
      mult_21_C247_n531, mult_21_C247_n530, mult_21_C247_n529, 
      mult_21_C247_n528, mult_21_C247_n527, mult_21_C247_n526, 
      mult_21_C247_n525, mult_21_C247_n524, mult_21_C247_n523, 
      mult_21_C247_n522, mult_21_C247_n521, mult_21_C247_n520, 
      mult_21_C247_n519, mult_21_C247_n518, mult_21_C247_n517, 
      mult_21_C247_n516, mult_21_C247_n515, mult_21_C247_n514, 
      mult_21_C247_n513, mult_21_C247_n512, mult_21_C247_n511, 
      mult_21_C247_n510, mult_21_C247_n509, mult_21_C247_n508, 
      mult_21_C247_n507, mult_21_C247_n506, mult_21_C247_n505, 
      mult_21_C247_n504, mult_21_C247_n503, mult_21_C247_n502, 
      mult_21_C247_n501, mult_21_C247_n500, mult_21_C247_n499, 
      mult_21_C247_n498, mult_21_C247_n497, mult_21_C247_n496, 
      mult_21_C247_n495, mult_21_C247_n494, mult_21_C247_n493, 
      mult_21_C247_n492, mult_21_C247_n491, mult_21_C247_n490, 
      mult_21_C247_n489, mult_21_C247_n488, mult_21_C247_n487, 
      mult_21_C247_n486, mult_21_C247_n485, mult_21_C247_n484, 
      mult_21_C247_n483, mult_21_C247_n482, mult_21_C247_n481, 
      mult_21_C247_n480, mult_21_C247_n479, mult_21_C247_n478, 
      mult_21_C247_n477, mult_21_C247_n476, mult_21_C247_n475, 
      mult_21_C247_n474, mult_21_C247_n473, mult_21_C247_n472, 
      mult_21_C247_n471, mult_21_C247_n470, mult_21_C247_n469, 
      mult_21_C247_n468, mult_21_C247_n467, mult_21_C247_n466, 
      mult_21_C247_n465, mult_21_C247_n464, mult_21_C247_n463, 
      mult_21_C247_n462, mult_21_C247_n461, mult_21_C247_n460, 
      mult_21_C247_n459, mult_21_C247_n458, mult_21_C247_n457, 
      mult_21_C247_n456, mult_21_C247_n455, mult_21_C247_n454, 
      mult_21_C247_n453, mult_21_C247_n452, mult_21_C247_n451, 
      mult_21_C247_n450, mult_21_C247_n449, mult_21_C247_n448, 
      mult_21_C247_n447, mult_21_C247_n446, mult_21_C247_n445, 
      mult_21_C247_n444, mult_21_C247_n443, mult_21_C247_n442, 
      mult_21_C247_n441, mult_21_C247_n440, mult_21_C247_n439, 
      mult_21_C247_n438, mult_21_C247_n437, mult_21_C247_n436, 
      mult_21_C247_n435, mult_21_C247_n434, mult_21_C247_n433, 
      mult_21_C247_n432, mult_21_C247_n431, mult_21_C247_n430, 
      mult_21_C247_n429, mult_21_C247_n428, mult_21_C247_n427, 
      mult_21_C247_n426, mult_21_C247_n425, mult_21_C247_n424, 
      mult_21_C247_n423, mult_21_C247_n422, mult_21_C247_n421, 
      mult_21_C247_n420, mult_21_C247_n419, mult_21_C247_n418, 
      mult_21_C247_n417, mult_21_C247_n416, mult_21_C247_n415, 
      mult_21_C247_n414, mult_21_C247_n413, mult_21_C247_n412, 
      mult_21_C247_n411, mult_21_C247_n410, mult_21_C247_n409, 
      mult_21_C247_n408, mult_21_C247_n407, mult_21_C247_n406, 
      mult_21_C247_n405, mult_21_C247_n404, mult_21_C247_n403, 
      mult_21_C247_n402, mult_21_C247_n401, mult_21_C247_n400, 
      mult_21_C247_n399, mult_21_C247_n398, mult_21_C247_n397, 
      mult_21_C247_n396, mult_21_C247_n395, mult_21_C247_n394, 
      mult_21_C247_n393, mult_21_C247_n392, mult_21_C247_n391, 
      mult_21_C247_n390, mult_21_C247_n389, mult_21_C247_n388, 
      mult_21_C247_n387, mult_21_C247_n386, mult_21_C247_n385, 
      mult_21_C247_n384, mult_21_C247_n383, mult_21_C247_n382, 
      mult_21_C247_n381, mult_21_C247_n380, mult_21_C247_n379, 
      mult_21_C247_n378, mult_21_C247_n377, mult_21_C247_n376, 
      mult_21_C247_n375, mult_21_C247_n374, mult_21_C247_n373, 
      mult_21_C247_n372, mult_21_C247_n371, mult_21_C247_n370, 
      mult_21_C247_n369, mult_21_C247_n368, mult_21_C247_n367, 
      mult_21_C247_n366, mult_21_C247_n365, mult_21_C247_n364, 
      mult_21_C247_n363, mult_21_C247_n362, mult_21_C247_n361, 
      mult_21_C247_n360, mult_21_C247_n359, mult_21_C247_n358, 
      mult_21_C247_n357, mult_21_C247_n356, mult_21_C247_n355, 
      mult_21_C247_n354, mult_21_C247_n353, mult_21_C247_n352, 
      mult_21_C247_n351, mult_21_C247_n350, mult_21_C247_n349, 
      mult_21_C247_n348, mult_21_C247_n347, mult_21_C247_n346, 
      mult_21_C247_n345, mult_21_C247_n344, mult_21_C247_n343, 
      mult_21_C247_n342, mult_21_C247_n341, mult_21_C247_n340, 
      mult_21_C247_n339, mult_21_C247_n338, mult_21_C247_n337, 
      mult_21_C247_n336, mult_21_C247_n335, mult_21_C247_n334, 
      mult_21_C247_n333, mult_21_C247_n332, mult_21_C247_n331, 
      mult_21_C247_n330, mult_21_C247_n329, mult_21_C247_n328, 
      mult_21_C247_n327, mult_21_C247_n326, mult_21_C247_n325, 
      mult_21_C247_n324, mult_21_C247_n323, mult_21_C247_n322, 
      mult_21_C247_n321, mult_21_C247_n320, mult_21_C247_n319, 
      mult_21_C247_n318, mult_21_C247_n317, mult_21_C247_n316, 
      mult_21_C247_n315, mult_21_C247_n314, mult_21_C247_n313, 
      mult_21_C247_n312, mult_21_C247_n311, mult_21_C247_n310, 
      mult_21_C247_n309, mult_21_C247_n308, mult_21_C247_n307, 
      mult_21_C247_n306, mult_21_C247_n305, mult_21_C247_n304, 
      mult_21_C247_n303, mult_21_C247_n302, mult_21_C247_n301, 
      mult_21_C247_n300, mult_21_C247_n299, mult_21_C247_n298, 
      mult_21_C247_n297, mult_21_C247_n296, mult_21_C247_n295, 
      mult_21_C247_n294, mult_21_C247_n293, mult_21_C247_n292, 
      mult_21_C247_n291, mult_21_C247_n290, mult_21_C247_n289, 
      mult_21_C247_n288, mult_21_C247_n287, mult_21_C247_n286, 
      mult_21_C247_n285, mult_21_C247_n284, mult_21_C247_n283, 
      mult_21_C247_n282, mult_21_C247_n281, mult_21_C247_n280, 
      mult_21_C247_n279, mult_21_C247_n278, mult_21_C247_n277, 
      mult_21_C247_n276, mult_21_C247_n275, mult_21_C247_n274, 
      mult_21_C247_n273, mult_21_C247_n272, mult_21_C247_n271, 
      mult_21_C247_n270, mult_21_C247_n269, mult_21_C247_n268, 
      mult_21_C247_n267, mult_21_C247_n266, mult_21_C247_n265, 
      mult_21_C247_n264, mult_21_C247_n263, mult_21_C247_n262, 
      mult_21_C247_n261, mult_21_C247_n260, mult_21_C247_n259, 
      mult_21_C247_n258, mult_21_C247_n257, mult_21_C247_n256, 
      mult_21_C247_n255, mult_21_C247_n254, mult_21_C247_n253, 
      mult_21_C247_n252, mult_21_C247_n251, mult_21_C247_n250, 
      mult_21_C247_n249, mult_21_C247_n248, mult_21_C247_n247, 
      mult_21_C247_n246, mult_21_C247_n245, mult_21_C247_n244, 
      mult_21_C247_n243, mult_21_C247_n242, mult_21_C247_n241, 
      mult_21_C247_n240, mult_21_C247_n239, mult_21_C247_n238, 
      mult_21_C247_n237, mult_21_C247_n236, mult_21_C247_n235, 
      mult_21_C247_n234, mult_21_C247_n233, mult_21_C247_n232, 
      mult_21_C247_n231, mult_21_C247_n230, mult_21_C247_n229, 
      mult_21_C247_n228, mult_21_C247_n227, mult_21_C247_n226, 
      mult_21_C247_n225, mult_21_C247_n224, mult_21_C247_n223, 
      mult_21_C247_n222, mult_21_C247_n221, mult_21_C247_n220, 
      mult_21_C247_n219, mult_21_C247_n218, mult_21_C247_n217, 
      mult_21_C247_n216, mult_21_C247_n215, mult_21_C247_n214, 
      mult_21_C247_n213, mult_21_C247_n212, mult_21_C247_n211, 
      mult_21_C247_n210, mult_21_C247_n209, mult_21_C247_n208, 
      mult_21_C247_n207, mult_21_C247_n206, mult_21_C247_n205, 
      mult_21_C247_n204, mult_21_C247_n203, mult_21_C247_n202, 
      mult_21_C247_n186, mult_21_C247_n185, mult_21_C247_n184, 
      mult_21_C247_n183, mult_21_C247_n182, mult_21_C247_n181, 
      mult_21_C247_n180, mult_21_C247_n179, mult_21_C247_n178, 
      mult_21_C247_n177, mult_21_C247_n176, mult_21_C247_n175, 
      mult_21_C247_n174, mult_21_C247_n173, mult_21_C247_n172, 
      mult_21_C247_n171, mult_21_C247_n170, mult_21_C247_n169, 
      mult_21_C247_n168, mult_21_C247_n167, mult_21_C247_n166, 
      mult_21_C247_n165, mult_21_C247_n164, mult_21_C247_n163, 
      mult_21_C247_n162, mult_21_C247_n161, mult_21_C247_n160, 
      mult_21_C247_n159, mult_21_C247_n158, mult_21_C247_n157, 
      mult_21_C247_n156, mult_21_C247_n104, mult_21_C247_n99, mult_21_C247_n94,
      mult_21_C247_n89, mult_21_C247_n84, mult_21_C247_n80, mult_21_C247_n73, 
      mult_21_C247_n66, mult_21_C247_n58, mult_21_C247_n50, mult_21_C247_n42, 
      mult_21_C249_n1454, mult_21_C249_n1453, mult_21_C249_n1452, 
      mult_21_C249_n1451, mult_21_C249_n1450, mult_21_C249_n1449, 
      mult_21_C249_n1448, mult_21_C249_n1447, mult_21_C249_n1446, 
      mult_21_C249_n1445, mult_21_C249_n1444, mult_21_C249_n1443, 
      mult_21_C249_n1442, mult_21_C249_n1441, mult_21_C249_n1440, 
      mult_21_C249_n1439, mult_21_C249_n1438, mult_21_C249_n1437, 
      mult_21_C249_n1436, mult_21_C249_n1435, mult_21_C249_n1434, 
      mult_21_C249_n1433, mult_21_C249_n1432, mult_21_C249_n1431, 
      mult_21_C249_n1430, mult_21_C249_n1429, mult_21_C249_n1428, 
      mult_21_C249_n1427, mult_21_C249_n1426, mult_21_C249_n1425, 
      mult_21_C249_n1424, mult_21_C249_n1423, mult_21_C249_n1422, 
      mult_21_C249_n1421, mult_21_C249_n1420, mult_21_C249_n1419, 
      mult_21_C249_n1418, mult_21_C249_n1417, mult_21_C249_n1416, 
      mult_21_C249_n1415, mult_21_C249_n1414, mult_21_C249_n1413, 
      mult_21_C249_n1412, mult_21_C249_n1411, mult_21_C249_n1410, 
      mult_21_C249_n1409, mult_21_C249_n1408, mult_21_C249_n1407, 
      mult_21_C249_n1406, mult_21_C249_n1405, mult_21_C249_n1404, 
      mult_21_C249_n1403, mult_21_C249_n1402, mult_21_C249_n1401, 
      mult_21_C249_n1400, mult_21_C249_n1399, mult_21_C249_n1398, 
      mult_21_C249_n1397, mult_21_C249_n1396, mult_21_C249_n1395, 
      mult_21_C249_n1394, mult_21_C249_n1393, mult_21_C249_n1392, 
      mult_21_C249_n1391, mult_21_C249_n1390, mult_21_C249_n1389, 
      mult_21_C249_n1388, mult_21_C249_n1387, mult_21_C249_n1386, 
      mult_21_C249_n1385, mult_21_C249_n1384, mult_21_C249_n1383, 
      mult_21_C249_n1382, mult_21_C249_n1381, mult_21_C249_n1380, 
      mult_21_C249_n1379, mult_21_C249_n1378, mult_21_C249_n1377, 
      mult_21_C249_n1376, mult_21_C249_n1375, mult_21_C249_n1226, 
      mult_21_C249_n1225, mult_21_C249_n1224, mult_21_C249_n1223, 
      mult_21_C249_n1222, mult_21_C249_n1221, mult_21_C249_n1220, 
      mult_21_C249_n1219, mult_21_C249_n1218, mult_21_C249_n1217, 
      mult_21_C249_n1216, mult_21_C249_n1215, mult_21_C249_n1214, 
      mult_21_C249_n1213, mult_21_C249_n1212, mult_21_C249_n1211, 
      mult_21_C249_n1210, mult_21_C249_n1209, mult_21_C249_n1208, 
      mult_21_C249_n1207, mult_21_C249_n1206, mult_21_C249_n1205, 
      mult_21_C249_n1204, mult_21_C249_n1203, mult_21_C249_n1202, 
      mult_21_C249_n1201, mult_21_C249_n1200, mult_21_C249_n1199, 
      mult_21_C249_n1198, mult_21_C249_n1197, mult_21_C249_n1196, 
      mult_21_C249_n1195, mult_21_C249_n1194, mult_21_C249_n1193, 
      mult_21_C249_n1192, mult_21_C249_n1191, mult_21_C249_n1190, 
      mult_21_C249_n1189, mult_21_C249_n1188, mult_21_C249_n1187, 
      mult_21_C249_n1186, mult_21_C249_n1185, mult_21_C249_n1184, 
      mult_21_C249_n1183, mult_21_C249_n1182, mult_21_C249_n1181, 
      mult_21_C249_n1180, mult_21_C249_n1179, mult_21_C249_n1178, 
      mult_21_C249_n1177, mult_21_C249_n1176, mult_21_C249_n1175, 
      mult_21_C249_n1174, mult_21_C249_n1173, mult_21_C249_n1172, 
      mult_21_C249_n1171, mult_21_C249_n1170, mult_21_C249_n1169, 
      mult_21_C249_n1168, mult_21_C249_n1167, mult_21_C249_n1166, 
      mult_21_C249_n1165, mult_21_C249_n1164, mult_21_C249_n1163, 
      mult_21_C249_n1162, mult_21_C249_n1161, mult_21_C249_n1160, 
      mult_21_C249_n1159, mult_21_C249_n1158, mult_21_C249_n1157, 
      mult_21_C249_n1156, mult_21_C249_n1155, mult_21_C249_n1154, 
      mult_21_C249_n1153, mult_21_C249_n1152, mult_21_C249_n1151, 
      mult_21_C249_n1150, mult_21_C249_n1149, mult_21_C249_n1148, 
      mult_21_C249_n1147, mult_21_C249_n1146, mult_21_C249_n1145, 
      mult_21_C249_n1144, mult_21_C249_n1143, mult_21_C249_n1142, 
      mult_21_C249_n1141, mult_21_C249_n1140, mult_21_C249_n1139, 
      mult_21_C249_n1138, mult_21_C249_n1137, mult_21_C249_n1136, 
      mult_21_C249_n1135, mult_21_C249_n1134, mult_21_C249_n1133, 
      mult_21_C249_n1132, mult_21_C249_n1131, mult_21_C249_n1130, 
      mult_21_C249_n1129, mult_21_C249_n1128, mult_21_C249_n1127, 
      mult_21_C249_n1126, mult_21_C249_n1125, mult_21_C249_n1124, 
      mult_21_C249_n1123, mult_21_C249_n1122, mult_21_C249_n1121, 
      mult_21_C249_n1120, mult_21_C249_n1119, mult_21_C249_n1118, 
      mult_21_C249_n1117, mult_21_C249_n1116, mult_21_C249_n1115, 
      mult_21_C249_n1114, mult_21_C249_n1113, mult_21_C249_n1112, 
      mult_21_C249_n1111, mult_21_C249_n1110, mult_21_C249_n1109, 
      mult_21_C249_n1108, mult_21_C249_n1107, mult_21_C249_n1106, 
      mult_21_C249_n1105, mult_21_C249_n1104, mult_21_C249_n1103, 
      mult_21_C249_n1102, mult_21_C249_n1101, mult_21_C249_n1100, 
      mult_21_C249_n1099, mult_21_C249_n1098, mult_21_C249_n1097, 
      mult_21_C249_n1096, mult_21_C249_n1095, mult_21_C249_n1094, 
      mult_21_C249_n1093, mult_21_C249_n1092, mult_21_C249_n1091, 
      mult_21_C249_n1090, mult_21_C249_n1089, mult_21_C249_n1088, 
      mult_21_C249_n1087, mult_21_C249_n1086, mult_21_C249_n1085, 
      mult_21_C249_n1084, mult_21_C249_n1083, mult_21_C249_n1082, 
      mult_21_C249_n1081, mult_21_C249_n1080, mult_21_C249_n1079, 
      mult_21_C249_n1078, mult_21_C249_n1077, mult_21_C249_n1076, 
      mult_21_C249_n1075, mult_21_C249_n1074, mult_21_C249_n1073, 
      mult_21_C249_n1072, mult_21_C249_n1071, mult_21_C249_n1070, 
      mult_21_C249_n1069, mult_21_C249_n1068, mult_21_C249_n1067, 
      mult_21_C249_n1066, mult_21_C249_n1065, mult_21_C249_n1064, 
      mult_21_C249_n1063, mult_21_C249_n1062, mult_21_C249_n1061, 
      mult_21_C249_n1060, mult_21_C249_n1059, mult_21_C249_n1058, 
      mult_21_C249_n1057, mult_21_C249_n1056, mult_21_C249_n1055, 
      mult_21_C249_n1054, mult_21_C249_n1053, mult_21_C249_n1052, 
      mult_21_C249_n1051, mult_21_C249_n1050, mult_21_C249_n1049, 
      mult_21_C249_n1048, mult_21_C249_n1047, mult_21_C249_n1046, 
      mult_21_C249_n1045, mult_21_C249_n1044, mult_21_C249_n1043, 
      mult_21_C249_n1042, mult_21_C249_n1041, mult_21_C249_n1040, 
      mult_21_C249_n1039, mult_21_C249_n1038, mult_21_C249_n1037, 
      mult_21_C249_n1036, mult_21_C249_n1035, mult_21_C249_n1034, 
      mult_21_C249_n1033, mult_21_C249_n1032, mult_21_C249_n1031, 
      mult_21_C249_n1030, mult_21_C249_n1029, mult_21_C249_n1028, 
      mult_21_C249_n1027, mult_21_C249_n1026, mult_21_C249_n1025, 
      mult_21_C249_n1024, mult_21_C249_n1023, mult_21_C249_n1022, 
      mult_21_C249_n1021, mult_21_C249_n1020, mult_21_C249_n1019, 
      mult_21_C249_n1018, mult_21_C249_n1017, mult_21_C249_n1016, 
      mult_21_C249_n1015, mult_21_C249_n1014, mult_21_C249_n1013, 
      mult_21_C249_n1012, mult_21_C249_n1011, mult_21_C249_n1010, 
      mult_21_C249_n1009, mult_21_C249_n1008, mult_21_C249_n1007, 
      mult_21_C249_n1006, mult_21_C249_n1005, mult_21_C249_n1004, 
      mult_21_C249_n1003, mult_21_C249_n1002, mult_21_C249_n1001, 
      mult_21_C249_n1000, mult_21_C249_n999, mult_21_C249_n998, 
      mult_21_C249_n997, mult_21_C249_n996, mult_21_C249_n995, 
      mult_21_C249_n994, mult_21_C249_n993, mult_21_C249_n992, 
      mult_21_C249_n991, mult_21_C249_n990, mult_21_C249_n989, 
      mult_21_C249_n988, mult_21_C249_n987, mult_21_C249_n986, 
      mult_21_C249_n985, mult_21_C249_n984, mult_21_C249_n983, 
      mult_21_C249_n982, mult_21_C249_n981, mult_21_C249_n980, 
      mult_21_C249_n979, mult_21_C249_n978, mult_21_C249_n977, 
      mult_21_C249_n976, mult_21_C249_n975, mult_21_C249_n974, 
      mult_21_C249_n973, mult_21_C249_n972, mult_21_C249_n971, 
      mult_21_C249_n970, mult_21_C249_n969, mult_21_C249_n968, 
      mult_21_C249_n967, mult_21_C249_n966, mult_21_C249_n965, 
      mult_21_C249_n964, mult_21_C249_n963, mult_21_C249_n962, 
      mult_21_C249_n961, mult_21_C249_n960, mult_21_C249_n959, 
      mult_21_C249_n958, mult_21_C249_n957, mult_21_C249_n956, 
      mult_21_C249_n955, mult_21_C249_n953, mult_21_C249_n952, 
      mult_21_C249_n951, mult_21_C249_n950, mult_21_C249_n949, 
      mult_21_C249_n948, mult_21_C249_n947, mult_21_C249_n946, 
      mult_21_C249_n945, mult_21_C249_n944, mult_21_C249_n943, 
      mult_21_C249_n942, mult_21_C249_n941, mult_21_C249_n940, 
      mult_21_C249_n939, mult_21_C249_n923, mult_21_C249_n922, 
      mult_21_C249_n921, mult_21_C249_n920, mult_21_C249_n919, 
      mult_21_C249_n918, mult_21_C249_n917, mult_21_C249_n916, 
      mult_21_C249_n915, mult_21_C249_n914, mult_21_C249_n913, 
      mult_21_C249_n912, mult_21_C249_n911, mult_21_C249_n910, 
      mult_21_C249_n909, mult_21_C249_n908, mult_21_C249_n907, 
      mult_21_C249_n906, mult_21_C249_n905, mult_21_C249_n904, 
      mult_21_C249_n903, mult_21_C249_n902, mult_21_C249_n901, 
      mult_21_C249_n900, mult_21_C249_n899, mult_21_C249_n898, 
      mult_21_C249_n897, mult_21_C249_n896, mult_21_C249_n895, 
      mult_21_C249_n894, mult_21_C249_n893, mult_21_C249_n892, 
      mult_21_C249_n891, mult_21_C249_n890, mult_21_C249_n889, 
      mult_21_C249_n888, mult_21_C249_n887, mult_21_C249_n886, 
      mult_21_C249_n885, mult_21_C249_n884, mult_21_C249_n883, 
      mult_21_C249_n882, mult_21_C249_n881, mult_21_C249_n880, 
      mult_21_C249_n879, mult_21_C249_n878, mult_21_C249_n877, 
      mult_21_C249_n876, mult_21_C249_n875, mult_21_C249_n874, 
      mult_21_C249_n873, mult_21_C249_n872, mult_21_C249_n871, 
      mult_21_C249_n870, mult_21_C249_n869, mult_21_C249_n868, 
      mult_21_C249_n867, mult_21_C249_n866, mult_21_C249_n865, 
      mult_21_C249_n864, mult_21_C249_n863, mult_21_C249_n862, 
      mult_21_C249_n861, mult_21_C249_n860, mult_21_C249_n859, 
      mult_21_C249_n858, mult_21_C249_n857, mult_21_C249_n856, 
      mult_21_C249_n855, mult_21_C249_n854, mult_21_C249_n853, 
      mult_21_C249_n852, mult_21_C249_n851, mult_21_C249_n850, 
      mult_21_C249_n849, mult_21_C249_n848, mult_21_C249_n847, 
      mult_21_C249_n846, mult_21_C249_n845, mult_21_C249_n844, 
      mult_21_C249_n843, mult_21_C249_n842, mult_21_C249_n841, 
      mult_21_C249_n840, mult_21_C249_n839, mult_21_C249_n838, 
      mult_21_C249_n837, mult_21_C249_n836, mult_21_C249_n835, 
      mult_21_C249_n834, mult_21_C249_n833, mult_21_C249_n832, 
      mult_21_C249_n831, mult_21_C249_n830, mult_21_C249_n829, 
      mult_21_C249_n828, mult_21_C249_n827, mult_21_C249_n826, 
      mult_21_C249_n825, mult_21_C249_n824, mult_21_C249_n823, 
      mult_21_C249_n822, mult_21_C249_n821, mult_21_C249_n820, 
      mult_21_C249_n819, mult_21_C249_n818, mult_21_C249_n817, 
      mult_21_C249_n816, mult_21_C249_n815, mult_21_C249_n814, 
      mult_21_C249_n813, mult_21_C249_n812, mult_21_C249_n811, 
      mult_21_C249_n810, mult_21_C249_n809, mult_21_C249_n808, 
      mult_21_C249_n807, mult_21_C249_n806, mult_21_C249_n805, 
      mult_21_C249_n804, mult_21_C249_n803, mult_21_C249_n802, 
      mult_21_C249_n801, mult_21_C249_n800, mult_21_C249_n799, 
      mult_21_C249_n798, mult_21_C249_n797, mult_21_C249_n796, 
      mult_21_C249_n795, mult_21_C249_n794, mult_21_C249_n793, 
      mult_21_C249_n792, mult_21_C249_n791, mult_21_C249_n790, 
      mult_21_C249_n789, mult_21_C249_n788, mult_21_C249_n787, 
      mult_21_C249_n786, mult_21_C249_n785, mult_21_C249_n784, 
      mult_21_C249_n783, mult_21_C249_n782, mult_21_C249_n781, 
      mult_21_C249_n780, mult_21_C249_n779, mult_21_C249_n778, 
      mult_21_C249_n777, mult_21_C249_n776, mult_21_C249_n775, 
      mult_21_C249_n774, mult_21_C249_n773, mult_21_C249_n772, 
      mult_21_C249_n771, mult_21_C249_n770, mult_21_C249_n769, 
      mult_21_C249_n768, mult_21_C249_n767, mult_21_C249_n766, 
      mult_21_C249_n765, mult_21_C249_n764, mult_21_C249_n763, 
      mult_21_C249_n762, mult_21_C249_n761, mult_21_C249_n760, 
      mult_21_C249_n759, mult_21_C249_n758, mult_21_C249_n757, 
      mult_21_C249_n756, mult_21_C249_n755, mult_21_C249_n754, 
      mult_21_C249_n753, mult_21_C249_n752, mult_21_C249_n751, 
      mult_21_C249_n750, mult_21_C249_n749, mult_21_C249_n748, 
      mult_21_C249_n747, mult_21_C249_n746, mult_21_C249_n745, 
      mult_21_C249_n744, mult_21_C249_n743, mult_21_C249_n742, 
      mult_21_C249_n741, mult_21_C249_n740, mult_21_C249_n739, 
      mult_21_C249_n738, mult_21_C249_n737, mult_21_C249_n736, 
      mult_21_C249_n735, mult_21_C249_n734, mult_21_C249_n733, 
      mult_21_C249_n732, mult_21_C249_n731, mult_21_C249_n730, 
      mult_21_C249_n729, mult_21_C249_n728, mult_21_C249_n727, 
      mult_21_C249_n726, mult_21_C249_n725, mult_21_C249_n724, 
      mult_21_C249_n723, mult_21_C249_n722, mult_21_C249_n721, 
      mult_21_C249_n720, mult_21_C249_n719, mult_21_C249_n718, 
      mult_21_C249_n717, mult_21_C249_n716, mult_21_C249_n715, 
      mult_21_C249_n714, mult_21_C249_n713, mult_21_C249_n712, 
      mult_21_C249_n711, mult_21_C249_n710, mult_21_C249_n709, 
      mult_21_C249_n708, mult_21_C249_n707, mult_21_C249_n706, 
      mult_21_C249_n705, mult_21_C249_n704, mult_21_C249_n703, 
      mult_21_C249_n702, mult_21_C249_n701, mult_21_C249_n700, 
      mult_21_C249_n699, mult_21_C249_n698, mult_21_C249_n697, 
      mult_21_C249_n696, mult_21_C249_n695, mult_21_C249_n694, 
      mult_21_C249_n693, mult_21_C249_n692, mult_21_C249_n691, 
      mult_21_C249_n690, mult_21_C249_n689, mult_21_C249_n688, 
      mult_21_C249_n687, mult_21_C249_n686, mult_21_C249_n685, 
      mult_21_C249_n684, mult_21_C249_n683, mult_21_C249_n682, 
      mult_21_C249_n681, mult_21_C249_n680, mult_21_C249_n679, 
      mult_21_C249_n678, mult_21_C249_n677, mult_21_C249_n676, 
      mult_21_C249_n675, mult_21_C249_n674, mult_21_C249_n673, 
      mult_21_C249_n672, mult_21_C249_n671, mult_21_C249_n670, 
      mult_21_C249_n669, mult_21_C249_n668, mult_21_C249_n667, 
      mult_21_C249_n666, mult_21_C249_n665, mult_21_C249_n664, 
      mult_21_C249_n663, mult_21_C249_n662, mult_21_C249_n661, 
      mult_21_C249_n660, mult_21_C249_n659, mult_21_C249_n658, 
      mult_21_C249_n657, mult_21_C249_n656, mult_21_C249_n655, 
      mult_21_C249_n654, mult_21_C249_n653, mult_21_C249_n652, 
      mult_21_C249_n651, mult_21_C249_n650, mult_21_C249_n649, 
      mult_21_C249_n648, mult_21_C249_n647, mult_21_C249_n646, 
      mult_21_C249_n645, mult_21_C249_n644, mult_21_C249_n643, 
      mult_21_C249_n642, mult_21_C249_n641, mult_21_C249_n640, 
      mult_21_C249_n639, mult_21_C249_n638, mult_21_C249_n637, 
      mult_21_C249_n636, mult_21_C249_n635, mult_21_C249_n634, 
      mult_21_C249_n633, mult_21_C249_n632, mult_21_C249_n631, 
      mult_21_C249_n630, mult_21_C249_n629, mult_21_C249_n628, 
      mult_21_C249_n627, mult_21_C249_n626, mult_21_C249_n625, 
      mult_21_C249_n624, mult_21_C249_n623, mult_21_C249_n622, 
      mult_21_C249_n621, mult_21_C249_n620, mult_21_C249_n619, 
      mult_21_C249_n618, mult_21_C249_n617, mult_21_C249_n616, 
      mult_21_C249_n615, mult_21_C249_n614, mult_21_C249_n613, 
      mult_21_C249_n612, mult_21_C249_n611, mult_21_C249_n610, 
      mult_21_C249_n609, mult_21_C249_n608, mult_21_C249_n607, 
      mult_21_C249_n606, mult_21_C249_n605, mult_21_C249_n604, 
      mult_21_C249_n603, mult_21_C249_n602, mult_21_C249_n601, 
      mult_21_C249_n600, mult_21_C249_n599, mult_21_C249_n598, 
      mult_21_C249_n597, mult_21_C249_n596, mult_21_C249_n595, 
      mult_21_C249_n594, mult_21_C249_n593, mult_21_C249_n592, 
      mult_21_C249_n591, mult_21_C249_n590, mult_21_C249_n589, 
      mult_21_C249_n588, mult_21_C249_n587, mult_21_C249_n586, 
      mult_21_C249_n585, mult_21_C249_n584, mult_21_C249_n583, 
      mult_21_C249_n582, mult_21_C249_n581, mult_21_C249_n580, 
      mult_21_C249_n579, mult_21_C249_n578, mult_21_C249_n577, 
      mult_21_C249_n576, mult_21_C249_n575, mult_21_C249_n574, 
      mult_21_C249_n573, mult_21_C249_n572, mult_21_C249_n571, 
      mult_21_C249_n570, mult_21_C249_n569, mult_21_C249_n568, 
      mult_21_C249_n567, mult_21_C249_n566, mult_21_C249_n565, 
      mult_21_C249_n564, mult_21_C249_n563, mult_21_C249_n562, 
      mult_21_C249_n561, mult_21_C249_n560, mult_21_C249_n559, 
      mult_21_C249_n558, mult_21_C249_n557, mult_21_C249_n556, 
      mult_21_C249_n555, mult_21_C249_n554, mult_21_C249_n553, 
      mult_21_C249_n552, mult_21_C249_n551, mult_21_C249_n550, 
      mult_21_C249_n549, mult_21_C249_n548, mult_21_C249_n547, 
      mult_21_C249_n546, mult_21_C249_n545, mult_21_C249_n544, 
      mult_21_C249_n543, mult_21_C249_n542, mult_21_C249_n541, 
      mult_21_C249_n540, mult_21_C249_n539, mult_21_C249_n538, 
      mult_21_C249_n537, mult_21_C249_n536, mult_21_C249_n535, 
      mult_21_C249_n534, mult_21_C249_n533, mult_21_C249_n532, 
      mult_21_C249_n531, mult_21_C249_n530, mult_21_C249_n529, 
      mult_21_C249_n528, mult_21_C249_n527, mult_21_C249_n526, 
      mult_21_C249_n525, mult_21_C249_n524, mult_21_C249_n523, 
      mult_21_C249_n522, mult_21_C249_n521, mult_21_C249_n520, 
      mult_21_C249_n519, mult_21_C249_n518, mult_21_C249_n517, 
      mult_21_C249_n516, mult_21_C249_n515, mult_21_C249_n514, 
      mult_21_C249_n513, mult_21_C249_n512, mult_21_C249_n511, 
      mult_21_C249_n510, mult_21_C249_n509, mult_21_C249_n508, 
      mult_21_C249_n507, mult_21_C249_n506, mult_21_C249_n505, 
      mult_21_C249_n504, mult_21_C249_n503, mult_21_C249_n502, 
      mult_21_C249_n501, mult_21_C249_n500, mult_21_C249_n499, 
      mult_21_C249_n498, mult_21_C249_n497, mult_21_C249_n496, 
      mult_21_C249_n495, mult_21_C249_n494, mult_21_C249_n493, 
      mult_21_C249_n492, mult_21_C249_n491, mult_21_C249_n490, 
      mult_21_C249_n489, mult_21_C249_n488, mult_21_C249_n487, 
      mult_21_C249_n486, mult_21_C249_n485, mult_21_C249_n484, 
      mult_21_C249_n483, mult_21_C249_n482, mult_21_C249_n481, 
      mult_21_C249_n480, mult_21_C249_n479, mult_21_C249_n478, 
      mult_21_C249_n477, mult_21_C249_n476, mult_21_C249_n475, 
      mult_21_C249_n474, mult_21_C249_n473, mult_21_C249_n472, 
      mult_21_C249_n471, mult_21_C249_n470, mult_21_C249_n469, 
      mult_21_C249_n468, mult_21_C249_n467, mult_21_C249_n466, 
      mult_21_C249_n465, mult_21_C249_n464, mult_21_C249_n463, 
      mult_21_C249_n462, mult_21_C249_n461, mult_21_C249_n460, 
      mult_21_C249_n459, mult_21_C249_n458, mult_21_C249_n457, 
      mult_21_C249_n456, mult_21_C249_n455, mult_21_C249_n454, 
      mult_21_C249_n453, mult_21_C249_n452, mult_21_C249_n451, 
      mult_21_C249_n450, mult_21_C249_n449, mult_21_C249_n448, 
      mult_21_C249_n447, mult_21_C249_n446, mult_21_C249_n445, 
      mult_21_C249_n444, mult_21_C249_n443, mult_21_C249_n442, 
      mult_21_C249_n441, mult_21_C249_n440, mult_21_C249_n439, 
      mult_21_C249_n438, mult_21_C249_n437, mult_21_C249_n436, 
      mult_21_C249_n435, mult_21_C249_n434, mult_21_C249_n433, 
      mult_21_C249_n432, mult_21_C249_n431, mult_21_C249_n430, 
      mult_21_C249_n429, mult_21_C249_n428, mult_21_C249_n427, 
      mult_21_C249_n426, mult_21_C249_n425, mult_21_C249_n424, 
      mult_21_C249_n423, mult_21_C249_n422, mult_21_C249_n421, 
      mult_21_C249_n420, mult_21_C249_n419, mult_21_C249_n418, 
      mult_21_C249_n417, mult_21_C249_n416, mult_21_C249_n415, 
      mult_21_C249_n414, mult_21_C249_n413, mult_21_C249_n412, 
      mult_21_C249_n411, mult_21_C249_n410, mult_21_C249_n409, 
      mult_21_C249_n408, mult_21_C249_n407, mult_21_C249_n406, 
      mult_21_C249_n405, mult_21_C249_n404, mult_21_C249_n403, 
      mult_21_C249_n402, mult_21_C249_n401, mult_21_C249_n400, 
      mult_21_C249_n399, mult_21_C249_n398, mult_21_C249_n397, 
      mult_21_C249_n396, mult_21_C249_n395, mult_21_C249_n394, 
      mult_21_C249_n393, mult_21_C249_n392, mult_21_C249_n391, 
      mult_21_C249_n390, mult_21_C249_n389, mult_21_C249_n388, 
      mult_21_C249_n387, mult_21_C249_n386, mult_21_C249_n385, 
      mult_21_C249_n384, mult_21_C249_n383, mult_21_C249_n382, 
      mult_21_C249_n381, mult_21_C249_n380, mult_21_C249_n379, 
      mult_21_C249_n378, mult_21_C249_n377, mult_21_C249_n376, 
      mult_21_C249_n375, mult_21_C249_n374, mult_21_C249_n373, 
      mult_21_C249_n372, mult_21_C249_n371, mult_21_C249_n370, 
      mult_21_C249_n369, mult_21_C249_n368, mult_21_C249_n367, 
      mult_21_C249_n366, mult_21_C249_n365, mult_21_C249_n364, 
      mult_21_C249_n363, mult_21_C249_n362, mult_21_C249_n361, 
      mult_21_C249_n360, mult_21_C249_n359, mult_21_C249_n358, 
      mult_21_C249_n357, mult_21_C249_n356, mult_21_C249_n355, 
      mult_21_C249_n354, mult_21_C249_n353, mult_21_C249_n352, 
      mult_21_C249_n351, mult_21_C249_n350, mult_21_C249_n349, 
      mult_21_C249_n348, mult_21_C249_n347, mult_21_C249_n346, 
      mult_21_C249_n345, mult_21_C249_n344, mult_21_C249_n343, 
      mult_21_C249_n342, mult_21_C249_n341, mult_21_C249_n340, 
      mult_21_C249_n339, mult_21_C249_n338, mult_21_C249_n337, 
      mult_21_C249_n336, mult_21_C249_n335, mult_21_C249_n334, 
      mult_21_C249_n333, mult_21_C249_n332, mult_21_C249_n331, 
      mult_21_C249_n330, mult_21_C249_n329, mult_21_C249_n328, 
      mult_21_C249_n327, mult_21_C249_n326, mult_21_C249_n325, 
      mult_21_C249_n324, mult_21_C249_n323, mult_21_C249_n322, 
      mult_21_C249_n321, mult_21_C249_n320, mult_21_C249_n319, 
      mult_21_C249_n318, mult_21_C249_n317, mult_21_C249_n316, 
      mult_21_C249_n315, mult_21_C249_n314, mult_21_C249_n313, 
      mult_21_C249_n312, mult_21_C249_n311, mult_21_C249_n310, 
      mult_21_C249_n309, mult_21_C249_n308, mult_21_C249_n307, 
      mult_21_C249_n306, mult_21_C249_n305, mult_21_C249_n304, 
      mult_21_C249_n303, mult_21_C249_n302, mult_21_C249_n301, 
      mult_21_C249_n300, mult_21_C249_n299, mult_21_C249_n298, 
      mult_21_C249_n297, mult_21_C249_n296, mult_21_C249_n295, 
      mult_21_C249_n294, mult_21_C249_n293, mult_21_C249_n292, 
      mult_21_C249_n291, mult_21_C249_n290, mult_21_C249_n289, 
      mult_21_C249_n288, mult_21_C249_n287, mult_21_C249_n286, 
      mult_21_C249_n285, mult_21_C249_n284, mult_21_C249_n283, 
      mult_21_C249_n282, mult_21_C249_n281, mult_21_C249_n280, 
      mult_21_C249_n279, mult_21_C249_n278, mult_21_C249_n277, 
      mult_21_C249_n276, mult_21_C249_n275, mult_21_C249_n274, 
      mult_21_C249_n273, mult_21_C249_n272, mult_21_C249_n271, 
      mult_21_C249_n270, mult_21_C249_n269, mult_21_C249_n268, 
      mult_21_C249_n267, mult_21_C249_n266, mult_21_C249_n265, 
      mult_21_C249_n264, mult_21_C249_n263, mult_21_C249_n262, 
      mult_21_C249_n261, mult_21_C249_n260, mult_21_C249_n259, 
      mult_21_C249_n258, mult_21_C249_n257, mult_21_C249_n256, 
      mult_21_C249_n255, mult_21_C249_n254, mult_21_C249_n253, 
      mult_21_C249_n252, mult_21_C249_n251, mult_21_C249_n250, 
      mult_21_C249_n249, mult_21_C249_n248, mult_21_C249_n247, 
      mult_21_C249_n246, mult_21_C249_n245, mult_21_C249_n244, 
      mult_21_C249_n243, mult_21_C249_n242, mult_21_C249_n241, 
      mult_21_C249_n240, mult_21_C249_n239, mult_21_C249_n238, 
      mult_21_C249_n237, mult_21_C249_n236, mult_21_C249_n235, 
      mult_21_C249_n234, mult_21_C249_n233, mult_21_C249_n232, 
      mult_21_C249_n231, mult_21_C249_n230, mult_21_C249_n229, 
      mult_21_C249_n228, mult_21_C249_n227, mult_21_C249_n226, 
      mult_21_C249_n225, mult_21_C249_n224, mult_21_C249_n223, 
      mult_21_C249_n222, mult_21_C249_n221, mult_21_C249_n220, 
      mult_21_C249_n219, mult_21_C249_n218, mult_21_C249_n217, 
      mult_21_C249_n216, mult_21_C249_n215, mult_21_C249_n214, 
      mult_21_C249_n213, mult_21_C249_n212, mult_21_C249_n211, 
      mult_21_C249_n210, mult_21_C249_n209, mult_21_C249_n208, 
      mult_21_C249_n207, mult_21_C249_n206, mult_21_C249_n205, 
      mult_21_C249_n204, mult_21_C249_n203, mult_21_C249_n202, 
      mult_21_C249_n186, mult_21_C249_n185, mult_21_C249_n184, 
      mult_21_C249_n183, mult_21_C249_n182, mult_21_C249_n181, 
      mult_21_C249_n180, mult_21_C249_n179, mult_21_C249_n178, 
      mult_21_C249_n177, mult_21_C249_n176, mult_21_C249_n175, 
      mult_21_C249_n174, mult_21_C249_n173, mult_21_C249_n172, 
      mult_21_C249_n171, mult_21_C249_n170, mult_21_C249_n169, 
      mult_21_C249_n168, mult_21_C249_n167, mult_21_C249_n166, 
      mult_21_C249_n165, mult_21_C249_n164, mult_21_C249_n163, 
      mult_21_C249_n162, mult_21_C249_n161, mult_21_C249_n160, 
      mult_21_C249_n159, mult_21_C249_n158, mult_21_C249_n157, 
      mult_21_C249_n156, mult_21_C249_n104, mult_21_C249_n99, mult_21_C249_n94,
      mult_21_C249_n89, mult_21_C249_n84, mult_21_C249_n80, mult_21_C249_n73, 
      mult_21_C249_n66, mult_21_C249_n58, mult_21_C249_n50, mult_21_C249_n42 : 
      std_logic;

begin
   avs_readdata <= ( avs_readdata_31_port, avs_readdata_30_port, 
      avs_readdata_29_port, avs_readdata_28_port, avs_readdata_27_port, 
      avs_readdata_26_port, avs_readdata_25_port, avs_readdata_24_port, 
      avs_readdata_23_port, avs_readdata_22_port, avs_readdata_21_port, 
      avs_readdata_20_port, avs_readdata_19_port, avs_readdata_18_port, 
      avs_readdata_17_port, avs_readdata_16_port, avs_readdata_15_port, 
      avs_readdata_14_port, avs_readdata_13_port, avs_readdata_12_port, 
      avs_readdata_11_port, avs_readdata_10_port, avs_readdata_9_port, 
      avs_readdata_8_port, avs_readdata_7_port, avs_readdata_6_port, 
      avs_readdata_5_port, avs_readdata_4_port, avs_readdata_3_port, 
      avs_readdata_2_port, avs_readdata_1_port, avs_readdata_0_port );
   clk_out <= clk;
   stop_sim <= stop_sim_port;
   
   U3 : OAI22D1 port map( A1 => N63, A2 => n4, B1 => n5, B2 => n697, Z => n201)
                           ;
   U4 : AOI21D1 port map( A1 => out_busy, A2 => n694, B => n684, Z => n5);
   U7 : AOI22D1 port map( A1 => N1978, A2 => n267, B1 => N2010, B2 => n674, Z 
                           => n10);
   U9 : AOI22D1 port map( A1 => N2011, A2 => n12, B1 => avs_readdata_30_port, 
                           B2 => n676, Z => n15);
   U12 : AOI22D1 port map( A1 => N1980, A2 => n267, B1 => N2012, B2 => n674, Z 
                           => n16);
   U14 : AOI22D1 port map( A1 => N2013, A2 => n674, B1 => avs_readdata_28_port,
                           B2 => n676, Z => n18);
   U17 : AOI22D1 port map( A1 => N1982, A2 => n267, B1 => N2014, B2 => n674, Z 
                           => n19);
   U19 : AOI22D1 port map( A1 => N2015, A2 => n674, B1 => avs_readdata_26_port,
                           B2 => n676, Z => n21);
   U22 : AOI22D1 port map( A1 => N1984, A2 => n267, B1 => N2016, B2 => n674, Z 
                           => n22);
   U24 : AOI22D1 port map( A1 => N2017, A2 => n674, B1 => avs_readdata_24_port,
                           B2 => n676, Z => n24);
   U27 : AOI22D1 port map( A1 => N1986, A2 => n267, B1 => N2018, B2 => n674, Z 
                           => n25);
   U29 : AOI22D1 port map( A1 => N2019, A2 => n12, B1 => avs_readdata_22_port, 
                           B2 => n676, Z => n27);
   U32 : AOI22D1 port map( A1 => N1988, A2 => n267, B1 => N2020, B2 => n674, Z 
                           => n28);
   U34 : AOI22D1 port map( A1 => N2021, A2 => n12, B1 => avs_readdata_20_port, 
                           B2 => n676, Z => n30);
   U37 : AOI22D1 port map( A1 => N1990, A2 => n267, B1 => N2022, B2 => n674, Z 
                           => n31);
   U39 : AOI22D1 port map( A1 => N2023, A2 => n12, B1 => avs_readdata_18_port, 
                           B2 => n676, Z => n33);
   U42 : AOI22D1 port map( A1 => N1992, A2 => n267, B1 => N2024, B2 => n674, Z 
                           => n34);
   U44 : AOI22D1 port map( A1 => N2025, A2 => n12, B1 => avs_readdata_16_port, 
                           B2 => n676, Z => n36);
   U47 : AOI22D1 port map( A1 => N1994, A2 => n267, B1 => N2026, B2 => n674, Z 
                           => n37);
   U49 : AOI22D1 port map( A1 => N2027, A2 => n12, B1 => avs_readdata_14_port, 
                           B2 => n676, Z => n39);
   U52 : AOI22D1 port map( A1 => N1996, A2 => n267, B1 => N2028, B2 => n12, Z 
                           => n40);
   U54 : AOI22D1 port map( A1 => N2029, A2 => n12, B1 => avs_readdata_12_port, 
                           B2 => n676, Z => n42);
   U57 : AOI22D1 port map( A1 => N1998, A2 => n267, B1 => N2030, B2 => n12, Z 
                           => n43);
   U59 : AOI22D1 port map( A1 => N2031, A2 => n12, B1 => avs_readdata_10_port, 
                           B2 => n676, Z => n45);
   U62 : AOI22D1 port map( A1 => N2000, A2 => n267, B1 => N2032, B2 => n12, Z 
                           => n46);
   U64 : AOI22D1 port map( A1 => N2033, A2 => n12, B1 => avs_readdata_8_port, 
                           B2 => n676, Z => n48);
   U67 : AOI22D1 port map( A1 => N2002, A2 => n267, B1 => N2034, B2 => n674, Z 
                           => n49);
   U69 : AOI22D1 port map( A1 => N2035, A2 => n12, B1 => avs_readdata_6_port, 
                           B2 => n676, Z => n51);
   U72 : AOI22D1 port map( A1 => N2004, A2 => n267, B1 => N2036, B2 => n674, Z 
                           => n52);
   U74 : AOI22D1 port map( A1 => N2037, A2 => n12, B1 => avs_readdata_4_port, 
                           B2 => n676, Z => n54);
   U77 : AOI22D1 port map( A1 => N2006, A2 => n267, B1 => N2038, B2 => n674, Z 
                           => n55);
   U79 : AOI22D1 port map( A1 => N2039, A2 => n12, B1 => avs_readdata_2_port, 
                           B2 => n676, Z => n57);
   U82 : AOI22D1 port map( A1 => N2008, A2 => n267, B1 => N2040, B2 => n674, Z 
                           => n58);
   U84 : AOI22D1 port map( A1 => N2041, A2 => n674, B1 => avs_readdata_0_port, 
                           B2 => n676, Z => n6100);
   U94 : AOI21D1 port map( A1 => n678, A2 => in_trigger, B => n72, Z => n70);
   U95 : OAI22D1 port map( A1 => n6400, A2 => n73, B1 => n74, B2 => n685, Z => 
                           n72);
   U96 : AOI22D1 port map( A1 => in_busy, A2 => n69, B1 => out_busy, B2 => n68,
                           Z => n73);
   U97 : EXNOR2D1 port map( A1 => n695, A2 => n76, Z => n234);
   U98 : AOI22D1 port map( A1 => n77, A2 => out_busy, B1 => n695, B2 => n685, Z
                           => n76);
   U100 : OAI22D1 port map( A1 => n697, A2 => n4, B1 => n79, B2 => n671, Z => 
                           n235);
   U103 : OAI32D1 port map( A1 => n684, A2 => N62, A3 => n695, B1 => n694, B2 
                           => n81, Z => n236);
   U105 : OAI32D1 port map( A1 => n696, A2 => n695, A3 => n78, B1 => out_busy, 
                           B2 => n685, Z => n81);
   U111 : OAI211D1 port map( A1 => n692, A2 => n84, B => n85, C => n86, Z => 
                           n237);
   U113 : OAI22D1 port map( A1 => n683, A2 => n88, B1 => n89, B2 => n693, Z => 
                           n238);
   U115 : EXNOR2D1 port map( A1 => in_busy, A2 => n161, Z => n239);
   U117 : AOI22D1 port map( A1 => avs_writedata(0), A2 => n677, B1 => 
                           out_trigger, B2 => n74, Z => n92);
   U122 : AOI22D1 port map( A1 => avs_writedata(0), A2 => n678, B1 => 
                           in_trigger, B2 => n96, Z => n95);
   U125 : EXNOR2D1 port map( A1 => n695, A2 => n672, Z => n154);
   U126 : EXNOR2D1 port map( A1 => n687, A2 => in_busy, Z => n156);
   U130 : AOI22D1 port map( A1 => odd, A2 => n91, B1 => n101, B2 => in_busy, Z 
                           => n100);
   U131 : OAI21D1 port map( A1 => in_counter_1_port, A2 => n690, B => n688, Z 
                           => n91);
   U200 : OA21M20D1 port map( A1 => n690, A2 => in_trigger, B => n176, Z => 
                           n161);
   comp_res_reg_4_30 : DFFRPQ1 port map( D => N3391, CK => clk, RB => resetn, Q
                           => comp_res_30_port);
   comp_res_reg_4_28 : DFFRPQ1 port map( D => N3389, CK => clk, RB => resetn, Q
                           => comp_res_28_port);
   comp_res_reg_4_26 : DFFRPQ1 port map( D => N3387, CK => clk, RB => resetn, Q
                           => comp_res_26_port);
   comp_res_reg_4_24 : DFFRPQ1 port map( D => N3385, CK => clk, RB => resetn, Q
                           => comp_res_24_port);
   comp_res_reg_4_22 : DFFRPQ1 port map( D => N3383, CK => clk, RB => resetn, Q
                           => comp_res_22_port);
   comp_res_reg_4_20 : DFFRPQ1 port map( D => N3381, CK => clk, RB => resetn, Q
                           => comp_res_20_port);
   comp_res_reg_4_18 : DFFRPQ1 port map( D => N3379, CK => clk, RB => resetn, Q
                           => comp_res_18_port);
   comp_res_reg_4_16 : DFFRPQ1 port map( D => N3377, CK => clk, RB => resetn, Q
                           => comp_res_16_port);
   comp_res_reg_4_14 : DFFRPQ1 port map( D => N3375, CK => clk, RB => resetn, Q
                           => comp_res_14_port);
   comp_res_reg_4_12 : DFFRPQ1 port map( D => N3373, CK => clk, RB => resetn, Q
                           => comp_res_12_port);
   comp_res_reg_4_10 : DFFRPQ1 port map( D => N3371, CK => clk, RB => resetn, Q
                           => comp_res_10_port);
   comp_res_reg_4_8 : DFFRPQ1 port map( D => N3369, CK => clk, RB => resetn, Q 
                           => comp_res_8_port);
   comp_res_reg_4_6 : DFFRPQ1 port map( D => N3367, CK => clk, RB => resetn, Q 
                           => comp_res_6_port);
   comp_res_reg_4_4 : DFFRPQ1 port map( D => N3365, CK => clk, RB => resetn, Q 
                           => comp_res_4_port);
   comp_res_reg_4_2 : DFFRPQ1 port map( D => N3363, CK => clk, RB => resetn, Q 
                           => comp_res_2_port);
   comp_res_reg_4_0 : DFFRPQ1 port map( D => N3361, CK => clk, RB => resetn, Q 
                           => comp_res_0_port);
   comp_res_reg_4_31 : DFFRPQ1 port map( D => N3392, CK => clk, RB => resetn, Q
                           => comp_res_31_port);
   comp_res_reg_4_29 : DFFRPQ1 port map( D => N3390, CK => clk, RB => resetn, Q
                           => comp_res_29_port);
   comp_res_reg_4_27 : DFFRPQ1 port map( D => N3388, CK => clk, RB => resetn, Q
                           => comp_res_27_port);
   comp_res_reg_4_25 : DFFRPQ1 port map( D => N3386, CK => clk, RB => resetn, Q
                           => comp_res_25_port);
   comp_res_reg_4_23 : DFFRPQ1 port map( D => N3384, CK => clk, RB => resetn, Q
                           => comp_res_23_port);
   comp_res_reg_4_21 : DFFRPQ1 port map( D => N3382, CK => clk, RB => resetn, Q
                           => comp_res_21_port);
   comp_res_reg_4_19 : DFFRPQ1 port map( D => N3380, CK => clk, RB => resetn, Q
                           => comp_res_19_port);
   comp_res_reg_4_17 : DFFRPQ1 port map( D => N3378, CK => clk, RB => resetn, Q
                           => comp_res_17_port);
   comp_res_reg_4_15 : DFFRPQ1 port map( D => N3376, CK => clk, RB => resetn, Q
                           => comp_res_15_port);
   comp_res_reg_4_13 : DFFRPQ1 port map( D => N3374, CK => clk, RB => resetn, Q
                           => comp_res_13_port);
   comp_res_reg_4_11 : DFFRPQ1 port map( D => N3372, CK => clk, RB => resetn, Q
                           => comp_res_11_port);
   comp_res_reg_4_9 : DFFRPQ1 port map( D => N3370, CK => clk, RB => resetn, Q 
                           => comp_res_9_port);
   comp_res_reg_4_7 : DFFRPQ1 port map( D => N3368, CK => clk, RB => resetn, Q 
                           => comp_res_7_port);
   comp_res_reg_4_5 : DFFRPQ1 port map( D => N3366, CK => clk, RB => resetn, Q 
                           => comp_res_5_port);
   comp_res_reg_4_3 : DFFRPQ1 port map( D => N3364, CK => clk, RB => resetn, Q 
                           => comp_res_3_port);
   comp_res_reg_4_1 : DFFRPQ1 port map( D => N3362, CK => clk, RB => resetn, Q 
                           => comp_res_1_port);
   comp_res_reg_3_30 : DFFRPQ1 port map( D => N3359, CK => clk, RB => resetn, Q
                           => comp_res_62_port);
   comp_res_reg_3_28 : DFFRPQ1 port map( D => N3357, CK => clk, RB => resetn, Q
                           => comp_res_60_port);
   comp_res_reg_3_26 : DFFRPQ1 port map( D => N3355, CK => clk, RB => resetn, Q
                           => comp_res_58_port);
   comp_res_reg_3_24 : DFFRPQ1 port map( D => N3353, CK => clk, RB => resetn, Q
                           => comp_res_56_port);
   comp_res_reg_3_22 : DFFRPQ1 port map( D => N3351, CK => clk, RB => resetn, Q
                           => comp_res_54_port);
   comp_res_reg_3_20 : DFFRPQ1 port map( D => N3349, CK => clk, RB => resetn, Q
                           => comp_res_52_port);
   comp_res_reg_3_18 : DFFRPQ1 port map( D => N3347, CK => clk, RB => resetn, Q
                           => comp_res_50_port);
   comp_res_reg_3_16 : DFFRPQ1 port map( D => N3345, CK => clk, RB => resetn, Q
                           => comp_res_48_port);
   comp_res_reg_3_14 : DFFRPQ1 port map( D => N3343, CK => clk, RB => resetn, Q
                           => comp_res_46_port);
   comp_res_reg_3_12 : DFFRPQ1 port map( D => N3341, CK => clk, RB => resetn, Q
                           => comp_res_44_port);
   comp_res_reg_3_10 : DFFRPQ1 port map( D => N3339, CK => clk, RB => resetn, Q
                           => comp_res_42_port);
   comp_res_reg_3_8 : DFFRPQ1 port map( D => N3337, CK => clk, RB => resetn, Q 
                           => comp_res_40_port);
   comp_res_reg_3_6 : DFFRPQ1 port map( D => N3335, CK => clk, RB => resetn, Q 
                           => comp_res_38_port);
   comp_res_reg_3_4 : DFFRPQ1 port map( D => N3333, CK => clk, RB => resetn, Q 
                           => comp_res_36_port);
   comp_res_reg_3_2 : DFFRPQ1 port map( D => N3331, CK => clk, RB => resetn, Q 
                           => comp_res_34_port);
   comp_res_reg_2_30 : DFFRPQ1 port map( D => N3327, CK => clk, RB => resetn, Q
                           => comp_res_94_port);
   comp_res_reg_2_28 : DFFRPQ1 port map( D => N3325, CK => clk, RB => resetn, Q
                           => comp_res_92_port);
   comp_res_reg_2_26 : DFFRPQ1 port map( D => N3323, CK => clk, RB => resetn, Q
                           => comp_res_90_port);
   comp_res_reg_2_24 : DFFRPQ1 port map( D => N3321, CK => clk, RB => resetn, Q
                           => comp_res_88_port);
   comp_res_reg_2_22 : DFFRPQ1 port map( D => N3319, CK => clk, RB => resetn, Q
                           => comp_res_86_port);
   comp_res_reg_2_20 : DFFRPQ1 port map( D => N3317, CK => clk, RB => resetn, Q
                           => comp_res_84_port);
   comp_res_reg_2_18 : DFFRPQ1 port map( D => N3315, CK => clk, RB => resetn, Q
                           => comp_res_82_port);
   comp_res_reg_2_16 : DFFRPQ1 port map( D => N3313, CK => clk, RB => resetn, Q
                           => comp_res_80_port);
   comp_res_reg_2_14 : DFFRPQ1 port map( D => N3311, CK => clk, RB => resetn, Q
                           => comp_res_78_port);
   comp_res_reg_2_12 : DFFRPQ1 port map( D => N3309, CK => clk, RB => resetn, Q
                           => comp_res_76_port);
   comp_res_reg_2_10 : DFFRPQ1 port map( D => N3307, CK => clk, RB => resetn, Q
                           => comp_res_74_port);
   comp_res_reg_2_8 : DFFRPQ1 port map( D => N3305, CK => clk, RB => resetn, Q 
                           => comp_res_72_port);
   comp_res_reg_2_6 : DFFRPQ1 port map( D => N3303, CK => clk, RB => resetn, Q 
                           => comp_res_70_port);
   comp_res_reg_2_4 : DFFRPQ1 port map( D => N3301, CK => clk, RB => resetn, Q 
                           => comp_res_68_port);
   comp_res_reg_2_2 : DFFRPQ1 port map( D => N3299, CK => clk, RB => resetn, Q 
                           => comp_res_66_port);
   comp_res_reg_1_30 : DFFRPQ1 port map( D => N3295, CK => clk, RB => resetn, Q
                           => comp_res_126_port);
   comp_res_reg_1_28 : DFFRPQ1 port map( D => N3293, CK => clk, RB => resetn, Q
                           => comp_res_124_port);
   comp_res_reg_1_26 : DFFRPQ1 port map( D => N3291, CK => clk, RB => resetn, Q
                           => comp_res_122_port);
   comp_res_reg_1_24 : DFFRPQ1 port map( D => N3289, CK => clk, RB => resetn, Q
                           => comp_res_120_port);
   comp_res_reg_1_22 : DFFRPQ1 port map( D => N3287, CK => clk, RB => resetn, Q
                           => comp_res_118_port);
   comp_res_reg_1_20 : DFFRPQ1 port map( D => N3285, CK => clk, RB => resetn, Q
                           => comp_res_116_port);
   comp_res_reg_1_18 : DFFRPQ1 port map( D => N3283, CK => clk, RB => resetn, Q
                           => comp_res_114_port);
   comp_res_reg_1_16 : DFFRPQ1 port map( D => N3281, CK => clk, RB => resetn, Q
                           => comp_res_112_port);
   comp_res_reg_1_14 : DFFRPQ1 port map( D => N3279, CK => clk, RB => resetn, Q
                           => comp_res_110_port);
   comp_res_reg_1_12 : DFFRPQ1 port map( D => N3277, CK => clk, RB => resetn, Q
                           => comp_res_108_port);
   comp_res_reg_1_10 : DFFRPQ1 port map( D => N3275, CK => clk, RB => resetn, Q
                           => comp_res_106_port);
   comp_res_reg_1_8 : DFFRPQ1 port map( D => N3273, CK => clk, RB => resetn, Q 
                           => comp_res_104_port);
   comp_res_reg_1_6 : DFFRPQ1 port map( D => N3271, CK => clk, RB => resetn, Q 
                           => comp_res_102_port);
   comp_res_reg_1_4 : DFFRPQ1 port map( D => N3269, CK => clk, RB => resetn, Q 
                           => comp_res_100_port);
   comp_res_reg_1_2 : DFFRPQ1 port map( D => N3267, CK => clk, RB => resetn, Q 
                           => comp_res_98_port);
   comp_res_reg_0_30 : DFFRPQ1 port map( D => N3263, CK => clk, RB => resetn, Q
                           => comp_res_158_port);
   comp_res_reg_0_28 : DFFRPQ1 port map( D => N3261, CK => clk, RB => resetn, Q
                           => comp_res_156_port);
   comp_res_reg_0_26 : DFFRPQ1 port map( D => N3259, CK => clk, RB => resetn, Q
                           => comp_res_154_port);
   comp_res_reg_0_24 : DFFRPQ1 port map( D => N3257, CK => clk, RB => resetn, Q
                           => comp_res_152_port);
   comp_res_reg_0_22 : DFFRPQ1 port map( D => N3255, CK => clk, RB => resetn, Q
                           => comp_res_150_port);
   comp_res_reg_0_20 : DFFRPQ1 port map( D => N3253, CK => clk, RB => resetn, Q
                           => comp_res_148_port);
   comp_res_reg_0_18 : DFFRPQ1 port map( D => N3251, CK => clk, RB => resetn, Q
                           => comp_res_146_port);
   comp_res_reg_0_16 : DFFRPQ1 port map( D => N3249, CK => clk, RB => resetn, Q
                           => comp_res_144_port);
   comp_res_reg_0_14 : DFFRPQ1 port map( D => N3247, CK => clk, RB => resetn, Q
                           => comp_res_142_port);
   comp_res_reg_0_12 : DFFRPQ1 port map( D => N3245, CK => clk, RB => resetn, Q
                           => comp_res_140_port);
   comp_res_reg_0_10 : DFFRPQ1 port map( D => N3243, CK => clk, RB => resetn, Q
                           => comp_res_138_port);
   comp_res_reg_0_8 : DFFRPQ1 port map( D => N3241, CK => clk, RB => resetn, Q 
                           => comp_res_136_port);
   comp_res_reg_0_6 : DFFRPQ1 port map( D => N3239, CK => clk, RB => resetn, Q 
                           => comp_res_134_port);
   comp_res_reg_0_4 : DFFRPQ1 port map( D => N3237, CK => clk, RB => resetn, Q 
                           => comp_res_132_port);
   comp_res_reg_0_2 : DFFRPQ1 port map( D => N3235, CK => clk, RB => resetn, Q 
                           => comp_res_130_port);
   comp_res_reg_3_0 : DFFRPQ1 port map( D => N3329, CK => clk, RB => resetn, Q 
                           => comp_res_32_port);
   comp_res_reg_2_0 : DFFRPQ1 port map( D => N3297, CK => clk, RB => resetn, Q 
                           => comp_res_64_port);
   comp_res_reg_1_0 : DFFRPQ1 port map( D => N3265, CK => clk, RB => resetn, Q 
                           => comp_res_96_port);
   comp_res_reg_0_0 : DFFRPQ1 port map( D => N3233, CK => clk, RB => resetn, Q 
                           => comp_res_128_port);
   in_buf_reg_7_31 : DFERPQ1 port map( D => siso_data_in(15), CEB => n176, CK 
                           => clk, RB => resetn, Q => in_buf_31_port);
   in_buf_reg_7_29 : DFERPQ1 port map( D => siso_data_in(13), CEB => n176, CK 
                           => clk, RB => resetn, Q => in_buf_29_port);
   in_buf_reg_7_27 : DFERPQ1 port map( D => siso_data_in(11), CEB => n176, CK 
                           => clk, RB => resetn, Q => in_buf_27_port);
   in_buf_reg_7_25 : DFERPQ1 port map( D => siso_data_in(9), CEB => n176, CK =>
                           clk, RB => resetn, Q => in_buf_25_port);
   in_buf_reg_7_23 : DFERPQ1 port map( D => siso_data_in(7), CEB => n176, CK =>
                           clk, RB => resetn, Q => in_buf_23_port);
   in_buf_reg_7_21 : DFERPQ1 port map( D => siso_data_in(5), CEB => n176, CK =>
                           clk, RB => resetn, Q => in_buf_21_port);
   in_buf_reg_7_19 : DFERPQ1 port map( D => siso_data_in(3), CEB => n176, CK =>
                           clk, RB => resetn, Q => in_buf_19_port);
   in_buf_reg_7_17 : DFERPQ1 port map( D => siso_data_in(1), CEB => n176, CK =>
                           clk, RB => resetn, Q => in_buf_17_port);
   in_buf_reg_7_15 : DFERPQ1 port map( D => siso_data_in(15), CEB => n177, CK 
                           => clk, RB => resetn, Q => in_buf_15_port);
   in_buf_reg_7_13 : DFERPQ1 port map( D => siso_data_in(13), CEB => n177, CK 
                           => clk, RB => resetn, Q => in_buf_13_port);
   in_buf_reg_7_11 : DFERPQ1 port map( D => siso_data_in(11), CEB => n177, CK 
                           => clk, RB => resetn, Q => in_buf_11_port);
   in_buf_reg_7_9 : DFERPQ1 port map( D => siso_data_in(9), CEB => n177, CK => 
                           clk, RB => resetn, Q => in_buf_9_port);
   in_buf_reg_7_7 : DFERPQ1 port map( D => siso_data_in(7), CEB => n177, CK => 
                           clk, RB => resetn, Q => in_buf_7_port);
   in_buf_reg_7_5 : DFERPQ1 port map( D => siso_data_in(5), CEB => n177, CK => 
                           clk, RB => resetn, Q => in_buf_5_port);
   in_buf_reg_7_3 : DFERPQ1 port map( D => siso_data_in(3), CEB => n177, CK => 
                           clk, RB => resetn, Q => in_buf_3_port);
   in_buf_reg_7_1 : DFERPQ1 port map( D => siso_data_in(1), CEB => n177, CK => 
                           clk, RB => resetn, Q => in_buf_1_port);
   comp_res_reg_3_31 : DFFRPQ1 port map( D => N3360, CK => clk, RB => resetn, Q
                           => comp_res_63_port);
   comp_res_reg_3_29 : DFFRPQ1 port map( D => N3358, CK => clk, RB => resetn, Q
                           => comp_res_61_port);
   comp_res_reg_3_27 : DFFRPQ1 port map( D => N3356, CK => clk, RB => resetn, Q
                           => comp_res_59_port);
   comp_res_reg_3_25 : DFFRPQ1 port map( D => N3354, CK => clk, RB => resetn, Q
                           => comp_res_57_port);
   comp_res_reg_3_23 : DFFRPQ1 port map( D => N3352, CK => clk, RB => resetn, Q
                           => comp_res_55_port);
   comp_res_reg_3_21 : DFFRPQ1 port map( D => N3350, CK => clk, RB => resetn, Q
                           => comp_res_53_port);
   comp_res_reg_3_19 : DFFRPQ1 port map( D => N3348, CK => clk, RB => resetn, Q
                           => comp_res_51_port);
   comp_res_reg_3_17 : DFFRPQ1 port map( D => N3346, CK => clk, RB => resetn, Q
                           => comp_res_49_port);
   comp_res_reg_3_15 : DFFRPQ1 port map( D => N3344, CK => clk, RB => resetn, Q
                           => comp_res_47_port);
   comp_res_reg_3_13 : DFFRPQ1 port map( D => N3342, CK => clk, RB => resetn, Q
                           => comp_res_45_port);
   comp_res_reg_3_11 : DFFRPQ1 port map( D => N3340, CK => clk, RB => resetn, Q
                           => comp_res_43_port);
   comp_res_reg_3_9 : DFFRPQ1 port map( D => N3338, CK => clk, RB => resetn, Q 
                           => comp_res_41_port);
   comp_res_reg_3_7 : DFFRPQ1 port map( D => N3336, CK => clk, RB => resetn, Q 
                           => comp_res_39_port);
   comp_res_reg_3_5 : DFFRPQ1 port map( D => N3334, CK => clk, RB => resetn, Q 
                           => comp_res_37_port);
   comp_res_reg_3_3 : DFFRPQ1 port map( D => N3332, CK => clk, RB => resetn, Q 
                           => comp_res_35_port);
   comp_res_reg_3_1 : DFFRPQ1 port map( D => N3330, CK => clk, RB => resetn, Q 
                           => comp_res_33_port);
   comp_res_reg_2_31 : DFFRPQ1 port map( D => N3328, CK => clk, RB => resetn, Q
                           => comp_res_95_port);
   comp_res_reg_2_29 : DFFRPQ1 port map( D => N3326, CK => clk, RB => resetn, Q
                           => comp_res_93_port);
   comp_res_reg_2_27 : DFFRPQ1 port map( D => N3324, CK => clk, RB => resetn, Q
                           => comp_res_91_port);
   comp_res_reg_2_25 : DFFRPQ1 port map( D => N3322, CK => clk, RB => resetn, Q
                           => comp_res_89_port);
   comp_res_reg_2_23 : DFFRPQ1 port map( D => N3320, CK => clk, RB => resetn, Q
                           => comp_res_87_port);
   comp_res_reg_2_21 : DFFRPQ1 port map( D => N3318, CK => clk, RB => resetn, Q
                           => comp_res_85_port);
   comp_res_reg_2_19 : DFFRPQ1 port map( D => N3316, CK => clk, RB => resetn, Q
                           => comp_res_83_port);
   comp_res_reg_2_17 : DFFRPQ1 port map( D => N3314, CK => clk, RB => resetn, Q
                           => comp_res_81_port);
   comp_res_reg_2_15 : DFFRPQ1 port map( D => N3312, CK => clk, RB => resetn, Q
                           => comp_res_79_port);
   comp_res_reg_2_13 : DFFRPQ1 port map( D => N3310, CK => clk, RB => resetn, Q
                           => comp_res_77_port);
   comp_res_reg_2_11 : DFFRPQ1 port map( D => N3308, CK => clk, RB => resetn, Q
                           => comp_res_75_port);
   comp_res_reg_2_9 : DFFRPQ1 port map( D => N3306, CK => clk, RB => resetn, Q 
                           => comp_res_73_port);
   comp_res_reg_2_7 : DFFRPQ1 port map( D => N3304, CK => clk, RB => resetn, Q 
                           => comp_res_71_port);
   comp_res_reg_2_5 : DFFRPQ1 port map( D => N3302, CK => clk, RB => resetn, Q 
                           => comp_res_69_port);
   comp_res_reg_2_3 : DFFRPQ1 port map( D => N3300, CK => clk, RB => resetn, Q 
                           => comp_res_67_port);
   comp_res_reg_2_1 : DFFRPQ1 port map( D => N3298, CK => clk, RB => resetn, Q 
                           => comp_res_65_port);
   in_buf_reg_3_31 : DFERPQ1 port map( D => siso_data_in(15), CEB => n168, CK 
                           => clk, RB => resetn, Q => in_buf_159_port);
   in_buf_reg_3_29 : DFERPQ1 port map( D => siso_data_in(13), CEB => n168, CK 
                           => clk, RB => resetn, Q => in_buf_157_port);
   in_buf_reg_3_27 : DFERPQ1 port map( D => siso_data_in(11), CEB => n168, CK 
                           => clk, RB => resetn, Q => in_buf_155_port);
   in_buf_reg_3_25 : DFERPQ1 port map( D => siso_data_in(9), CEB => n168, CK =>
                           clk, RB => resetn, Q => in_buf_153_port);
   in_buf_reg_3_23 : DFERPQ1 port map( D => siso_data_in(7), CEB => n168, CK =>
                           clk, RB => resetn, Q => in_buf_151_port);
   in_buf_reg_3_21 : DFERPQ1 port map( D => siso_data_in(5), CEB => n168, CK =>
                           clk, RB => resetn, Q => in_buf_149_port);
   in_buf_reg_3_19 : DFERPQ1 port map( D => siso_data_in(3), CEB => n168, CK =>
                           clk, RB => resetn, Q => in_buf_147_port);
   in_buf_reg_3_17 : DFERPQ1 port map( D => siso_data_in(1), CEB => n168, CK =>
                           clk, RB => resetn, Q => in_buf_145_port);
   in_buf_reg_3_15 : DFERPQ1 port map( D => siso_data_in(15), CEB => n169, CK 
                           => clk, RB => resetn, Q => in_buf_143_port);
   in_buf_reg_3_13 : DFERPQ1 port map( D => siso_data_in(13), CEB => n169, CK 
                           => clk, RB => resetn, Q => in_buf_141_port);
   in_buf_reg_3_11 : DFERPQ1 port map( D => siso_data_in(11), CEB => n169, CK 
                           => clk, RB => resetn, Q => in_buf_139_port);
   in_buf_reg_3_9 : DFERPQ1 port map( D => siso_data_in(9), CEB => n169, CK => 
                           clk, RB => resetn, Q => in_buf_137_port);
   in_buf_reg_3_7 : DFERPQ1 port map( D => siso_data_in(7), CEB => n169, CK => 
                           clk, RB => resetn, Q => in_buf_135_port);
   in_buf_reg_3_5 : DFERPQ1 port map( D => siso_data_in(5), CEB => n169, CK => 
                           clk, RB => resetn, Q => in_buf_133_port);
   in_buf_reg_3_3 : DFERPQ1 port map( D => siso_data_in(3), CEB => n169, CK => 
                           clk, RB => resetn, Q => in_buf_131_port);
   in_buf_reg_3_1 : DFERPQ1 port map( D => siso_data_in(1), CEB => n169, CK => 
                           clk, RB => resetn, Q => in_buf_129_port);
   in_buf_reg_2_31 : DFERPQ1 port map( D => siso_data_in(15), CEB => n166, CK 
                           => clk, RB => resetn, Q => in_buf_191_port);
   in_buf_reg_2_29 : DFERPQ1 port map( D => siso_data_in(13), CEB => n166, CK 
                           => clk, RB => resetn, Q => in_buf_189_port);
   in_buf_reg_2_27 : DFERPQ1 port map( D => siso_data_in(11), CEB => n166, CK 
                           => clk, RB => resetn, Q => in_buf_187_port);
   in_buf_reg_2_25 : DFERPQ1 port map( D => siso_data_in(9), CEB => n166, CK =>
                           clk, RB => resetn, Q => in_buf_185_port);
   in_buf_reg_2_23 : DFERPQ1 port map( D => siso_data_in(7), CEB => n166, CK =>
                           clk, RB => resetn, Q => in_buf_183_port);
   in_buf_reg_2_21 : DFERPQ1 port map( D => siso_data_in(5), CEB => n166, CK =>
                           clk, RB => resetn, Q => in_buf_181_port);
   in_buf_reg_2_19 : DFERPQ1 port map( D => siso_data_in(3), CEB => n166, CK =>
                           clk, RB => resetn, Q => in_buf_179_port);
   in_buf_reg_2_17 : DFERPQ1 port map( D => siso_data_in(1), CEB => n166, CK =>
                           clk, RB => resetn, Q => in_buf_177_port);
   in_buf_reg_6_31 : DFERPQ1 port map( D => siso_data_in(15), CEB => n174, CK 
                           => clk, RB => resetn, Q => in_buf_63_port);
   in_buf_reg_6_29 : DFERPQ1 port map( D => siso_data_in(13), CEB => n174, CK 
                           => clk, RB => resetn, Q => in_buf_61_port);
   in_buf_reg_6_27 : DFERPQ1 port map( D => siso_data_in(11), CEB => n174, CK 
                           => clk, RB => resetn, Q => in_buf_59_port);
   in_buf_reg_6_25 : DFERPQ1 port map( D => siso_data_in(9), CEB => n174, CK =>
                           clk, RB => resetn, Q => in_buf_57_port);
   in_buf_reg_6_23 : DFERPQ1 port map( D => siso_data_in(7), CEB => n174, CK =>
                           clk, RB => resetn, Q => in_buf_55_port);
   in_buf_reg_6_21 : DFERPQ1 port map( D => siso_data_in(5), CEB => n174, CK =>
                           clk, RB => resetn, Q => in_buf_53_port);
   in_buf_reg_6_19 : DFERPQ1 port map( D => siso_data_in(3), CEB => n174, CK =>
                           clk, RB => resetn, Q => in_buf_51_port);
   in_buf_reg_6_17 : DFERPQ1 port map( D => siso_data_in(1), CEB => n174, CK =>
                           clk, RB => resetn, Q => in_buf_49_port);
   in_buf_reg_2_15 : DFERPQ1 port map( D => siso_data_in(15), CEB => n167, CK 
                           => clk, RB => resetn, Q => in_buf_175_port);
   in_buf_reg_2_13 : DFERPQ1 port map( D => siso_data_in(13), CEB => n167, CK 
                           => clk, RB => resetn, Q => in_buf_173_port);
   in_buf_reg_2_11 : DFERPQ1 port map( D => siso_data_in(11), CEB => n167, CK 
                           => clk, RB => resetn, Q => in_buf_171_port);
   in_buf_reg_2_9 : DFERPQ1 port map( D => siso_data_in(9), CEB => n167, CK => 
                           clk, RB => resetn, Q => in_buf_169_port);
   in_buf_reg_2_7 : DFERPQ1 port map( D => siso_data_in(7), CEB => n167, CK => 
                           clk, RB => resetn, Q => in_buf_167_port);
   in_buf_reg_2_5 : DFERPQ1 port map( D => siso_data_in(5), CEB => n167, CK => 
                           clk, RB => resetn, Q => in_buf_165_port);
   in_buf_reg_2_3 : DFERPQ1 port map( D => siso_data_in(3), CEB => n167, CK => 
                           clk, RB => resetn, Q => in_buf_163_port);
   in_buf_reg_2_1 : DFERPQ1 port map( D => siso_data_in(1), CEB => n167, CK => 
                           clk, RB => resetn, Q => in_buf_161_port);
   in_buf_reg_6_15 : DFERPQ1 port map( D => siso_data_in(15), CEB => n175, CK 
                           => clk, RB => resetn, Q => in_buf_47_port);
   in_buf_reg_6_13 : DFERPQ1 port map( D => siso_data_in(13), CEB => n175, CK 
                           => clk, RB => resetn, Q => in_buf_45_port);
   in_buf_reg_6_11 : DFERPQ1 port map( D => siso_data_in(11), CEB => n175, CK 
                           => clk, RB => resetn, Q => in_buf_43_port);
   in_buf_reg_6_9 : DFERPQ1 port map( D => siso_data_in(9), CEB => n175, CK => 
                           clk, RB => resetn, Q => in_buf_41_port);
   in_buf_reg_6_7 : DFERPQ1 port map( D => siso_data_in(7), CEB => n175, CK => 
                           clk, RB => resetn, Q => in_buf_39_port);
   in_buf_reg_6_5 : DFERPQ1 port map( D => siso_data_in(5), CEB => n175, CK => 
                           clk, RB => resetn, Q => in_buf_37_port);
   in_buf_reg_6_3 : DFERPQ1 port map( D => siso_data_in(3), CEB => n175, CK => 
                           clk, RB => resetn, Q => in_buf_35_port);
   in_buf_reg_6_1 : DFERPQ1 port map( D => siso_data_in(1), CEB => n175, CK => 
                           clk, RB => resetn, Q => in_buf_33_port);
   in_buf_reg_5_31 : DFERPQ1 port map( D => siso_data_in(15), CEB => n172, CK 
                           => clk, RB => resetn, Q => in_buf_95_port);
   in_buf_reg_5_29 : DFERPQ1 port map( D => siso_data_in(13), CEB => n172, CK 
                           => clk, RB => resetn, Q => in_buf_93_port);
   in_buf_reg_5_27 : DFERPQ1 port map( D => siso_data_in(11), CEB => n172, CK 
                           => clk, RB => resetn, Q => in_buf_91_port);
   in_buf_reg_5_25 : DFERPQ1 port map( D => siso_data_in(9), CEB => n172, CK =>
                           clk, RB => resetn, Q => in_buf_89_port);
   in_buf_reg_5_23 : DFERPQ1 port map( D => siso_data_in(7), CEB => n172, CK =>
                           clk, RB => resetn, Q => in_buf_87_port);
   in_buf_reg_5_21 : DFERPQ1 port map( D => siso_data_in(5), CEB => n172, CK =>
                           clk, RB => resetn, Q => in_buf_85_port);
   in_buf_reg_5_19 : DFERPQ1 port map( D => siso_data_in(3), CEB => n172, CK =>
                           clk, RB => resetn, Q => in_buf_83_port);
   in_buf_reg_5_17 : DFERPQ1 port map( D => siso_data_in(1), CEB => n172, CK =>
                           clk, RB => resetn, Q => in_buf_81_port);
   in_buf_reg_5_15 : DFERPQ1 port map( D => siso_data_in(15), CEB => n173, CK 
                           => clk, RB => resetn, Q => in_buf_79_port);
   in_buf_reg_5_13 : DFERPQ1 port map( D => siso_data_in(13), CEB => n173, CK 
                           => clk, RB => resetn, Q => in_buf_77_port);
   in_buf_reg_5_11 : DFERPQ1 port map( D => siso_data_in(11), CEB => n173, CK 
                           => clk, RB => resetn, Q => in_buf_75_port);
   in_buf_reg_5_9 : DFERPQ1 port map( D => siso_data_in(9), CEB => n173, CK => 
                           clk, RB => resetn, Q => in_buf_73_port);
   in_buf_reg_5_7 : DFERPQ1 port map( D => siso_data_in(7), CEB => n173, CK => 
                           clk, RB => resetn, Q => in_buf_71_port);
   in_buf_reg_5_5 : DFERPQ1 port map( D => siso_data_in(5), CEB => n173, CK => 
                           clk, RB => resetn, Q => in_buf_69_port);
   in_buf_reg_5_3 : DFERPQ1 port map( D => siso_data_in(3), CEB => n173, CK => 
                           clk, RB => resetn, Q => in_buf_67_port);
   in_buf_reg_5_1 : DFERPQ1 port map( D => siso_data_in(1), CEB => n173, CK => 
                           clk, RB => resetn, Q => in_buf_65_port);
   comp_res_reg_1_31 : DFFRPQ1 port map( D => N3296, CK => clk, RB => resetn, Q
                           => comp_res_127_port);
   comp_res_reg_1_29 : DFFRPQ1 port map( D => N3294, CK => clk, RB => resetn, Q
                           => comp_res_125_port);
   comp_res_reg_1_27 : DFFRPQ1 port map( D => N3292, CK => clk, RB => resetn, Q
                           => comp_res_123_port);
   comp_res_reg_1_25 : DFFRPQ1 port map( D => N3290, CK => clk, RB => resetn, Q
                           => comp_res_121_port);
   comp_res_reg_1_23 : DFFRPQ1 port map( D => N3288, CK => clk, RB => resetn, Q
                           => comp_res_119_port);
   comp_res_reg_1_21 : DFFRPQ1 port map( D => N3286, CK => clk, RB => resetn, Q
                           => comp_res_117_port);
   comp_res_reg_1_19 : DFFRPQ1 port map( D => N3284, CK => clk, RB => resetn, Q
                           => comp_res_115_port);
   comp_res_reg_1_17 : DFFRPQ1 port map( D => N3282, CK => clk, RB => resetn, Q
                           => comp_res_113_port);
   comp_res_reg_1_15 : DFFRPQ1 port map( D => N3280, CK => clk, RB => resetn, Q
                           => comp_res_111_port);
   comp_res_reg_1_13 : DFFRPQ1 port map( D => N3278, CK => clk, RB => resetn, Q
                           => comp_res_109_port);
   comp_res_reg_1_11 : DFFRPQ1 port map( D => N3276, CK => clk, RB => resetn, Q
                           => comp_res_107_port);
   comp_res_reg_1_9 : DFFRPQ1 port map( D => N3274, CK => clk, RB => resetn, Q 
                           => comp_res_105_port);
   comp_res_reg_1_7 : DFFRPQ1 port map( D => N3272, CK => clk, RB => resetn, Q 
                           => comp_res_103_port);
   comp_res_reg_1_5 : DFFRPQ1 port map( D => N3270, CK => clk, RB => resetn, Q 
                           => comp_res_101_port);
   comp_res_reg_1_3 : DFFRPQ1 port map( D => N3268, CK => clk, RB => resetn, Q 
                           => comp_res_99_port);
   comp_res_reg_1_1 : DFFRPQ1 port map( D => N3266, CK => clk, RB => resetn, Q 
                           => comp_res_97_port);
   comp_res_reg_0_31 : DFFRPQ1 port map( D => N3264, CK => clk, RB => resetn, Q
                           => comp_res_159_port);
   comp_res_reg_0_29 : DFFRPQ1 port map( D => N3262, CK => clk, RB => resetn, Q
                           => comp_res_157_port);
   comp_res_reg_0_27 : DFFRPQ1 port map( D => N3260, CK => clk, RB => resetn, Q
                           => comp_res_155_port);
   comp_res_reg_0_25 : DFFRPQ1 port map( D => N3258, CK => clk, RB => resetn, Q
                           => comp_res_153_port);
   comp_res_reg_0_23 : DFFRPQ1 port map( D => N3256, CK => clk, RB => resetn, Q
                           => comp_res_151_port);
   comp_res_reg_0_21 : DFFRPQ1 port map( D => N3254, CK => clk, RB => resetn, Q
                           => comp_res_149_port);
   comp_res_reg_0_19 : DFFRPQ1 port map( D => N3252, CK => clk, RB => resetn, Q
                           => comp_res_147_port);
   comp_res_reg_0_17 : DFFRPQ1 port map( D => N3250, CK => clk, RB => resetn, Q
                           => comp_res_145_port);
   comp_res_reg_0_15 : DFFRPQ1 port map( D => N3248, CK => clk, RB => resetn, Q
                           => comp_res_143_port);
   comp_res_reg_0_13 : DFFRPQ1 port map( D => N3246, CK => clk, RB => resetn, Q
                           => comp_res_141_port);
   comp_res_reg_0_11 : DFFRPQ1 port map( D => N3244, CK => clk, RB => resetn, Q
                           => comp_res_139_port);
   comp_res_reg_0_9 : DFFRPQ1 port map( D => N3242, CK => clk, RB => resetn, Q 
                           => comp_res_137_port);
   comp_res_reg_0_7 : DFFRPQ1 port map( D => N3240, CK => clk, RB => resetn, Q 
                           => comp_res_135_port);
   comp_res_reg_0_5 : DFFRPQ1 port map( D => N3238, CK => clk, RB => resetn, Q 
                           => comp_res_133_port);
   comp_res_reg_0_3 : DFFRPQ1 port map( D => N3236, CK => clk, RB => resetn, Q 
                           => comp_res_131_port);
   comp_res_reg_0_1 : DFFRPQ1 port map( D => N3234, CK => clk, RB => resetn, Q 
                           => comp_res_129_port);
   in_buf_reg_1_31 : DFERPQ1 port map( D => siso_data_in(15), CEB => n164, CK 
                           => clk, RB => resetn, Q => in_buf_223_port);
   in_buf_reg_1_29 : DFERPQ1 port map( D => siso_data_in(13), CEB => n164, CK 
                           => clk, RB => resetn, Q => in_buf_221_port);
   in_buf_reg_1_27 : DFERPQ1 port map( D => siso_data_in(11), CEB => n164, CK 
                           => clk, RB => resetn, Q => in_buf_219_port);
   in_buf_reg_1_25 : DFERPQ1 port map( D => siso_data_in(9), CEB => n164, CK =>
                           clk, RB => resetn, Q => in_buf_217_port);
   in_buf_reg_1_23 : DFERPQ1 port map( D => siso_data_in(7), CEB => n164, CK =>
                           clk, RB => resetn, Q => in_buf_215_port);
   in_buf_reg_1_21 : DFERPQ1 port map( D => siso_data_in(5), CEB => n164, CK =>
                           clk, RB => resetn, Q => in_buf_213_port);
   in_buf_reg_1_19 : DFERPQ1 port map( D => siso_data_in(3), CEB => n164, CK =>
                           clk, RB => resetn, Q => in_buf_211_port);
   in_buf_reg_1_17 : DFERPQ1 port map( D => siso_data_in(1), CEB => n164, CK =>
                           clk, RB => resetn, Q => in_buf_209_port);
   in_buf_reg_1_15 : DFERPQ1 port map( D => siso_data_in(15), CEB => n165, CK 
                           => clk, RB => resetn, Q => in_buf_207_port);
   in_buf_reg_1_13 : DFERPQ1 port map( D => siso_data_in(13), CEB => n165, CK 
                           => clk, RB => resetn, Q => in_buf_205_port);
   in_buf_reg_1_11 : DFERPQ1 port map( D => siso_data_in(11), CEB => n165, CK 
                           => clk, RB => resetn, Q => in_buf_203_port);
   in_buf_reg_1_9 : DFERPQ1 port map( D => siso_data_in(9), CEB => n165, CK => 
                           clk, RB => resetn, Q => in_buf_201_port);
   in_buf_reg_1_7 : DFERPQ1 port map( D => siso_data_in(7), CEB => n165, CK => 
                           clk, RB => resetn, Q => in_buf_199_port);
   in_buf_reg_1_5 : DFERPQ1 port map( D => siso_data_in(5), CEB => n165, CK => 
                           clk, RB => resetn, Q => in_buf_197_port);
   in_buf_reg_1_3 : DFERPQ1 port map( D => siso_data_in(3), CEB => n165, CK => 
                           clk, RB => resetn, Q => in_buf_195_port);
   in_buf_reg_1_1 : DFERPQ1 port map( D => siso_data_in(1), CEB => n165, CK => 
                           clk, RB => resetn, Q => in_buf_193_port);
   in_buf_reg_4_31 : DFERPQ1 port map( D => siso_data_in(15), CEB => n170, CK 
                           => clk, RB => resetn, Q => in_buf_127_port);
   in_buf_reg_4_29 : DFERPQ1 port map( D => siso_data_in(13), CEB => n170, CK 
                           => clk, RB => resetn, Q => in_buf_125_port);
   in_buf_reg_4_27 : DFERPQ1 port map( D => siso_data_in(11), CEB => n170, CK 
                           => clk, RB => resetn, Q => in_buf_123_port);
   in_buf_reg_4_25 : DFERPQ1 port map( D => siso_data_in(9), CEB => n170, CK =>
                           clk, RB => resetn, Q => in_buf_121_port);
   in_buf_reg_4_23 : DFERPQ1 port map( D => siso_data_in(7), CEB => n170, CK =>
                           clk, RB => resetn, Q => in_buf_119_port);
   in_buf_reg_4_21 : DFERPQ1 port map( D => siso_data_in(5), CEB => n170, CK =>
                           clk, RB => resetn, Q => in_buf_117_port);
   in_buf_reg_4_19 : DFERPQ1 port map( D => siso_data_in(3), CEB => n170, CK =>
                           clk, RB => resetn, Q => in_buf_115_port);
   in_buf_reg_4_17 : DFERPQ1 port map( D => siso_data_in(1), CEB => n170, CK =>
                           clk, RB => resetn, Q => in_buf_113_port);
   in_buf_reg_0_31 : DFERPQ1 port map( D => siso_data_in(15), CEB => n162, CK 
                           => clk, RB => resetn, Q => in_buf_255_port);
   in_buf_reg_0_29 : DFERPQ1 port map( D => siso_data_in(13), CEB => n162, CK 
                           => clk, RB => resetn, Q => in_buf_253_port);
   in_buf_reg_0_27 : DFERPQ1 port map( D => siso_data_in(11), CEB => n162, CK 
                           => clk, RB => resetn, Q => in_buf_251_port);
   in_buf_reg_0_25 : DFERPQ1 port map( D => siso_data_in(9), CEB => n162, CK =>
                           clk, RB => resetn, Q => in_buf_249_port);
   in_buf_reg_0_23 : DFERPQ1 port map( D => siso_data_in(7), CEB => n162, CK =>
                           clk, RB => resetn, Q => in_buf_247_port);
   in_buf_reg_0_21 : DFERPQ1 port map( D => siso_data_in(5), CEB => n162, CK =>
                           clk, RB => resetn, Q => in_buf_245_port);
   in_buf_reg_0_19 : DFERPQ1 port map( D => siso_data_in(3), CEB => n162, CK =>
                           clk, RB => resetn, Q => in_buf_243_port);
   in_buf_reg_0_17 : DFERPQ1 port map( D => siso_data_in(1), CEB => n162, CK =>
                           clk, RB => resetn, Q => in_buf_241_port);
   in_buf_reg_0_15 : DFERPQ1 port map( D => siso_data_in(15), CEB => n163, CK 
                           => clk, RB => resetn, Q => in_buf_239_port);
   in_buf_reg_0_13 : DFERPQ1 port map( D => siso_data_in(13), CEB => n163, CK 
                           => clk, RB => resetn, Q => in_buf_237_port);
   in_buf_reg_0_11 : DFERPQ1 port map( D => siso_data_in(11), CEB => n163, CK 
                           => clk, RB => resetn, Q => in_buf_235_port);
   in_buf_reg_0_9 : DFERPQ1 port map( D => siso_data_in(9), CEB => n163, CK => 
                           clk, RB => resetn, Q => in_buf_233_port);
   in_buf_reg_0_7 : DFERPQ1 port map( D => siso_data_in(7), CEB => n163, CK => 
                           clk, RB => resetn, Q => in_buf_231_port);
   in_buf_reg_0_5 : DFERPQ1 port map( D => siso_data_in(5), CEB => n163, CK => 
                           clk, RB => resetn, Q => in_buf_229_port);
   in_buf_reg_0_3 : DFERPQ1 port map( D => siso_data_in(3), CEB => n163, CK => 
                           clk, RB => resetn, Q => in_buf_227_port);
   in_buf_reg_0_1 : DFERPQ1 port map( D => siso_data_in(1), CEB => n163, CK => 
                           clk, RB => resetn, Q => in_buf_225_port);
   in_buf_reg_4_15 : DFERPQ1 port map( D => siso_data_in(15), CEB => n171, CK 
                           => clk, RB => resetn, Q => in_buf_111_port);
   in_buf_reg_4_13 : DFERPQ1 port map( D => siso_data_in(13), CEB => n171, CK 
                           => clk, RB => resetn, Q => in_buf_109_port);
   in_buf_reg_4_11 : DFERPQ1 port map( D => siso_data_in(11), CEB => n171, CK 
                           => clk, RB => resetn, Q => in_buf_107_port);
   in_buf_reg_4_9 : DFERPQ1 port map( D => siso_data_in(9), CEB => n171, CK => 
                           clk, RB => resetn, Q => in_buf_105_port);
   in_buf_reg_4_7 : DFERPQ1 port map( D => siso_data_in(7), CEB => n171, CK => 
                           clk, RB => resetn, Q => in_buf_103_port);
   in_buf_reg_4_5 : DFERPQ1 port map( D => siso_data_in(5), CEB => n171, CK => 
                           clk, RB => resetn, Q => in_buf_101_port);
   in_buf_reg_4_3 : DFERPQ1 port map( D => siso_data_in(3), CEB => n171, CK => 
                           clk, RB => resetn, Q => in_buf_99_port);
   in_buf_reg_4_1 : DFERPQ1 port map( D => siso_data_in(1), CEB => n171, CK => 
                           clk, RB => resetn, Q => in_buf_97_port);
   in_buf_reg_7_30 : DFERPQ1 port map( D => siso_data_in(14), CEB => n176, CK 
                           => clk, RB => resetn, Q => in_buf_30_port);
   in_buf_reg_7_28 : DFERPQ1 port map( D => siso_data_in(12), CEB => n176, CK 
                           => clk, RB => resetn, Q => in_buf_28_port);
   in_buf_reg_7_26 : DFERPQ1 port map( D => siso_data_in(10), CEB => n176, CK 
                           => clk, RB => resetn, Q => in_buf_26_port);
   in_buf_reg_7_24 : DFERPQ1 port map( D => siso_data_in(8), CEB => n176, CK =>
                           clk, RB => resetn, Q => in_buf_24_port);
   in_buf_reg_7_22 : DFERPQ1 port map( D => siso_data_in(6), CEB => n176, CK =>
                           clk, RB => resetn, Q => in_buf_22_port);
   in_buf_reg_7_20 : DFERPQ1 port map( D => siso_data_in(4), CEB => n176, CK =>
                           clk, RB => resetn, Q => in_buf_20_port);
   in_buf_reg_7_18 : DFERPQ1 port map( D => siso_data_in(2), CEB => n176, CK =>
                           clk, RB => resetn, Q => in_buf_18_port);
   in_buf_reg_7_16 : DFERPQ1 port map( D => siso_data_in(0), CEB => n176, CK =>
                           clk, RB => resetn, Q => in_buf_16_port);
   in_buf_reg_7_14 : DFERPQ1 port map( D => siso_data_in(14), CEB => n177, CK 
                           => clk, RB => resetn, Q => in_buf_14_port);
   in_buf_reg_7_12 : DFERPQ1 port map( D => siso_data_in(12), CEB => n177, CK 
                           => clk, RB => resetn, Q => in_buf_12_port);
   in_buf_reg_7_10 : DFERPQ1 port map( D => siso_data_in(10), CEB => n177, CK 
                           => clk, RB => resetn, Q => in_buf_10_port);
   in_buf_reg_7_8 : DFERPQ1 port map( D => siso_data_in(8), CEB => n177, CK => 
                           clk, RB => resetn, Q => in_buf_8_port);
   in_buf_reg_7_6 : DFERPQ1 port map( D => siso_data_in(6), CEB => n177, CK => 
                           clk, RB => resetn, Q => in_buf_6_port);
   in_buf_reg_7_4 : DFERPQ1 port map( D => siso_data_in(4), CEB => n177, CK => 
                           clk, RB => resetn, Q => in_buf_4_port);
   in_buf_reg_7_2 : DFERPQ1 port map( D => siso_data_in(2), CEB => n177, CK => 
                           clk, RB => resetn, Q => in_buf_2_port);
   in_trigger_reg : DFFRPQ1 port map( D => n241, CK => clk, RB => resetn, Q => 
                           in_trigger);
   in_buf_reg_3_30 : DFERPQ1 port map( D => siso_data_in(14), CEB => n168, CK 
                           => clk, RB => resetn, Q => in_buf_158_port);
   in_buf_reg_3_28 : DFERPQ1 port map( D => siso_data_in(12), CEB => n168, CK 
                           => clk, RB => resetn, Q => in_buf_156_port);
   in_buf_reg_3_26 : DFERPQ1 port map( D => siso_data_in(10), CEB => n168, CK 
                           => clk, RB => resetn, Q => in_buf_154_port);
   in_buf_reg_3_24 : DFERPQ1 port map( D => siso_data_in(8), CEB => n168, CK =>
                           clk, RB => resetn, Q => in_buf_152_port);
   in_buf_reg_3_22 : DFERPQ1 port map( D => siso_data_in(6), CEB => n168, CK =>
                           clk, RB => resetn, Q => in_buf_150_port);
   in_buf_reg_3_20 : DFERPQ1 port map( D => siso_data_in(4), CEB => n168, CK =>
                           clk, RB => resetn, Q => in_buf_148_port);
   in_buf_reg_3_18 : DFERPQ1 port map( D => siso_data_in(2), CEB => n168, CK =>
                           clk, RB => resetn, Q => in_buf_146_port);
   in_buf_reg_3_16 : DFERPQ1 port map( D => siso_data_in(0), CEB => n168, CK =>
                           clk, RB => resetn, Q => in_buf_144_port);
   in_buf_reg_3_14 : DFERPQ1 port map( D => siso_data_in(14), CEB => n169, CK 
                           => clk, RB => resetn, Q => in_buf_142_port);
   in_buf_reg_3_12 : DFERPQ1 port map( D => siso_data_in(12), CEB => n169, CK 
                           => clk, RB => resetn, Q => in_buf_140_port);
   in_buf_reg_3_10 : DFERPQ1 port map( D => siso_data_in(10), CEB => n169, CK 
                           => clk, RB => resetn, Q => in_buf_138_port);
   in_buf_reg_3_8 : DFERPQ1 port map( D => siso_data_in(8), CEB => n169, CK => 
                           clk, RB => resetn, Q => in_buf_136_port);
   in_buf_reg_3_6 : DFERPQ1 port map( D => siso_data_in(6), CEB => n169, CK => 
                           clk, RB => resetn, Q => in_buf_134_port);
   in_buf_reg_3_4 : DFERPQ1 port map( D => siso_data_in(4), CEB => n169, CK => 
                           clk, RB => resetn, Q => in_buf_132_port);
   in_buf_reg_3_2 : DFERPQ1 port map( D => siso_data_in(2), CEB => n169, CK => 
                           clk, RB => resetn, Q => in_buf_130_port);
   in_buf_reg_2_30 : DFERPQ1 port map( D => siso_data_in(14), CEB => n166, CK 
                           => clk, RB => resetn, Q => in_buf_190_port);
   in_buf_reg_2_28 : DFERPQ1 port map( D => siso_data_in(12), CEB => n166, CK 
                           => clk, RB => resetn, Q => in_buf_188_port);
   in_buf_reg_2_26 : DFERPQ1 port map( D => siso_data_in(10), CEB => n166, CK 
                           => clk, RB => resetn, Q => in_buf_186_port);
   in_buf_reg_2_24 : DFERPQ1 port map( D => siso_data_in(8), CEB => n166, CK =>
                           clk, RB => resetn, Q => in_buf_184_port);
   in_buf_reg_2_22 : DFERPQ1 port map( D => siso_data_in(6), CEB => n166, CK =>
                           clk, RB => resetn, Q => in_buf_182_port);
   in_buf_reg_2_20 : DFERPQ1 port map( D => siso_data_in(4), CEB => n166, CK =>
                           clk, RB => resetn, Q => in_buf_180_port);
   in_buf_reg_2_18 : DFERPQ1 port map( D => siso_data_in(2), CEB => n166, CK =>
                           clk, RB => resetn, Q => in_buf_178_port);
   in_buf_reg_2_16 : DFERPQ1 port map( D => siso_data_in(0), CEB => n166, CK =>
                           clk, RB => resetn, Q => in_buf_176_port);
   in_buf_reg_6_30 : DFERPQ1 port map( D => siso_data_in(14), CEB => n174, CK 
                           => clk, RB => resetn, Q => in_buf_62_port);
   in_buf_reg_6_28 : DFERPQ1 port map( D => siso_data_in(12), CEB => n174, CK 
                           => clk, RB => resetn, Q => in_buf_60_port);
   in_buf_reg_6_26 : DFERPQ1 port map( D => siso_data_in(10), CEB => n174, CK 
                           => clk, RB => resetn, Q => in_buf_58_port);
   in_buf_reg_6_24 : DFERPQ1 port map( D => siso_data_in(8), CEB => n174, CK =>
                           clk, RB => resetn, Q => in_buf_56_port);
   in_buf_reg_6_22 : DFERPQ1 port map( D => siso_data_in(6), CEB => n174, CK =>
                           clk, RB => resetn, Q => in_buf_54_port);
   in_buf_reg_6_20 : DFERPQ1 port map( D => siso_data_in(4), CEB => n174, CK =>
                           clk, RB => resetn, Q => in_buf_52_port);
   in_buf_reg_6_18 : DFERPQ1 port map( D => siso_data_in(2), CEB => n174, CK =>
                           clk, RB => resetn, Q => in_buf_50_port);
   in_buf_reg_6_16 : DFERPQ1 port map( D => siso_data_in(0), CEB => n174, CK =>
                           clk, RB => resetn, Q => in_buf_48_port);
   in_buf_reg_2_14 : DFERPQ1 port map( D => siso_data_in(14), CEB => n167, CK 
                           => clk, RB => resetn, Q => in_buf_174_port);
   in_buf_reg_2_12 : DFERPQ1 port map( D => siso_data_in(12), CEB => n167, CK 
                           => clk, RB => resetn, Q => in_buf_172_port);
   in_buf_reg_2_10 : DFERPQ1 port map( D => siso_data_in(10), CEB => n167, CK 
                           => clk, RB => resetn, Q => in_buf_170_port);
   in_buf_reg_2_8 : DFERPQ1 port map( D => siso_data_in(8), CEB => n167, CK => 
                           clk, RB => resetn, Q => in_buf_168_port);
   in_buf_reg_2_6 : DFERPQ1 port map( D => siso_data_in(6), CEB => n167, CK => 
                           clk, RB => resetn, Q => in_buf_166_port);
   in_buf_reg_2_4 : DFERPQ1 port map( D => siso_data_in(4), CEB => n167, CK => 
                           clk, RB => resetn, Q => in_buf_164_port);
   in_buf_reg_2_2 : DFERPQ1 port map( D => siso_data_in(2), CEB => n167, CK => 
                           clk, RB => resetn, Q => in_buf_162_port);
   in_buf_reg_6_14 : DFERPQ1 port map( D => siso_data_in(14), CEB => n175, CK 
                           => clk, RB => resetn, Q => in_buf_46_port);
   in_buf_reg_6_12 : DFERPQ1 port map( D => siso_data_in(12), CEB => n175, CK 
                           => clk, RB => resetn, Q => in_buf_44_port);
   in_buf_reg_6_10 : DFERPQ1 port map( D => siso_data_in(10), CEB => n175, CK 
                           => clk, RB => resetn, Q => in_buf_42_port);
   in_buf_reg_6_8 : DFERPQ1 port map( D => siso_data_in(8), CEB => n175, CK => 
                           clk, RB => resetn, Q => in_buf_40_port);
   in_buf_reg_6_6 : DFERPQ1 port map( D => siso_data_in(6), CEB => n175, CK => 
                           clk, RB => resetn, Q => in_buf_38_port);
   in_buf_reg_6_4 : DFERPQ1 port map( D => siso_data_in(4), CEB => n175, CK => 
                           clk, RB => resetn, Q => in_buf_36_port);
   in_buf_reg_6_2 : DFERPQ1 port map( D => siso_data_in(2), CEB => n175, CK => 
                           clk, RB => resetn, Q => in_buf_34_port);
   in_buf_reg_5_30 : DFERPQ1 port map( D => siso_data_in(14), CEB => n172, CK 
                           => clk, RB => resetn, Q => in_buf_94_port);
   in_buf_reg_5_28 : DFERPQ1 port map( D => siso_data_in(12), CEB => n172, CK 
                           => clk, RB => resetn, Q => in_buf_92_port);
   in_buf_reg_5_26 : DFERPQ1 port map( D => siso_data_in(10), CEB => n172, CK 
                           => clk, RB => resetn, Q => in_buf_90_port);
   in_buf_reg_5_24 : DFERPQ1 port map( D => siso_data_in(8), CEB => n172, CK =>
                           clk, RB => resetn, Q => in_buf_88_port);
   in_buf_reg_5_22 : DFERPQ1 port map( D => siso_data_in(6), CEB => n172, CK =>
                           clk, RB => resetn, Q => in_buf_86_port);
   in_buf_reg_5_20 : DFERPQ1 port map( D => siso_data_in(4), CEB => n172, CK =>
                           clk, RB => resetn, Q => in_buf_84_port);
   in_buf_reg_5_18 : DFERPQ1 port map( D => siso_data_in(2), CEB => n172, CK =>
                           clk, RB => resetn, Q => in_buf_82_port);
   in_buf_reg_5_16 : DFERPQ1 port map( D => siso_data_in(0), CEB => n172, CK =>
                           clk, RB => resetn, Q => in_buf_80_port);
   in_buf_reg_5_14 : DFERPQ1 port map( D => siso_data_in(14), CEB => n173, CK 
                           => clk, RB => resetn, Q => in_buf_78_port);
   in_buf_reg_5_12 : DFERPQ1 port map( D => siso_data_in(12), CEB => n173, CK 
                           => clk, RB => resetn, Q => in_buf_76_port);
   in_buf_reg_5_10 : DFERPQ1 port map( D => siso_data_in(10), CEB => n173, CK 
                           => clk, RB => resetn, Q => in_buf_74_port);
   in_buf_reg_5_8 : DFERPQ1 port map( D => siso_data_in(8), CEB => n173, CK => 
                           clk, RB => resetn, Q => in_buf_72_port);
   in_buf_reg_5_6 : DFERPQ1 port map( D => siso_data_in(6), CEB => n173, CK => 
                           clk, RB => resetn, Q => in_buf_70_port);
   in_buf_reg_5_4 : DFERPQ1 port map( D => siso_data_in(4), CEB => n173, CK => 
                           clk, RB => resetn, Q => in_buf_68_port);
   in_buf_reg_5_2 : DFERPQ1 port map( D => siso_data_in(2), CEB => n173, CK => 
                           clk, RB => resetn, Q => in_buf_66_port);
   in_buf_reg_7_0 : DFERPQ1 port map( D => siso_data_in(0), CEB => n177, CK => 
                           clk, RB => resetn, Q => in_buf_0_port);
   in_buf_reg_1_30 : DFERPQ1 port map( D => siso_data_in(14), CEB => n164, CK 
                           => clk, RB => resetn, Q => in_buf_222_port);
   in_buf_reg_1_28 : DFERPQ1 port map( D => siso_data_in(12), CEB => n164, CK 
                           => clk, RB => resetn, Q => in_buf_220_port);
   in_buf_reg_1_26 : DFERPQ1 port map( D => siso_data_in(10), CEB => n164, CK 
                           => clk, RB => resetn, Q => in_buf_218_port);
   in_buf_reg_1_24 : DFERPQ1 port map( D => siso_data_in(8), CEB => n164, CK =>
                           clk, RB => resetn, Q => in_buf_216_port);
   in_buf_reg_1_22 : DFERPQ1 port map( D => siso_data_in(6), CEB => n164, CK =>
                           clk, RB => resetn, Q => in_buf_214_port);
   in_buf_reg_1_20 : DFERPQ1 port map( D => siso_data_in(4), CEB => n164, CK =>
                           clk, RB => resetn, Q => in_buf_212_port);
   in_buf_reg_1_18 : DFERPQ1 port map( D => siso_data_in(2), CEB => n164, CK =>
                           clk, RB => resetn, Q => in_buf_210_port);
   in_buf_reg_1_16 : DFERPQ1 port map( D => siso_data_in(0), CEB => n164, CK =>
                           clk, RB => resetn, Q => in_buf_208_port);
   in_buf_reg_1_14 : DFERPQ1 port map( D => siso_data_in(14), CEB => n165, CK 
                           => clk, RB => resetn, Q => in_buf_206_port);
   in_buf_reg_1_12 : DFERPQ1 port map( D => siso_data_in(12), CEB => n165, CK 
                           => clk, RB => resetn, Q => in_buf_204_port);
   in_buf_reg_1_10 : DFERPQ1 port map( D => siso_data_in(10), CEB => n165, CK 
                           => clk, RB => resetn, Q => in_buf_202_port);
   in_buf_reg_1_8 : DFERPQ1 port map( D => siso_data_in(8), CEB => n165, CK => 
                           clk, RB => resetn, Q => in_buf_200_port);
   in_buf_reg_1_6 : DFERPQ1 port map( D => siso_data_in(6), CEB => n165, CK => 
                           clk, RB => resetn, Q => in_buf_198_port);
   in_buf_reg_1_4 : DFERPQ1 port map( D => siso_data_in(4), CEB => n165, CK => 
                           clk, RB => resetn, Q => in_buf_196_port);
   in_buf_reg_1_2 : DFERPQ1 port map( D => siso_data_in(2), CEB => n165, CK => 
                           clk, RB => resetn, Q => in_buf_194_port);
   in_buf_reg_4_30 : DFERPQ1 port map( D => siso_data_in(14), CEB => n170, CK 
                           => clk, RB => resetn, Q => in_buf_126_port);
   in_buf_reg_4_28 : DFERPQ1 port map( D => siso_data_in(12), CEB => n170, CK 
                           => clk, RB => resetn, Q => in_buf_124_port);
   in_buf_reg_4_26 : DFERPQ1 port map( D => siso_data_in(10), CEB => n170, CK 
                           => clk, RB => resetn, Q => in_buf_122_port);
   in_buf_reg_4_24 : DFERPQ1 port map( D => siso_data_in(8), CEB => n170, CK =>
                           clk, RB => resetn, Q => in_buf_120_port);
   in_buf_reg_4_22 : DFERPQ1 port map( D => siso_data_in(6), CEB => n170, CK =>
                           clk, RB => resetn, Q => in_buf_118_port);
   in_buf_reg_4_20 : DFERPQ1 port map( D => siso_data_in(4), CEB => n170, CK =>
                           clk, RB => resetn, Q => in_buf_116_port);
   in_buf_reg_4_18 : DFERPQ1 port map( D => siso_data_in(2), CEB => n170, CK =>
                           clk, RB => resetn, Q => in_buf_114_port);
   in_buf_reg_4_16 : DFERPQ1 port map( D => siso_data_in(0), CEB => n170, CK =>
                           clk, RB => resetn, Q => in_buf_112_port);
   in_buf_reg_0_30 : DFERPQ1 port map( D => siso_data_in(14), CEB => n162, CK 
                           => clk, RB => resetn, Q => in_buf_254_port);
   in_buf_reg_0_28 : DFERPQ1 port map( D => siso_data_in(12), CEB => n162, CK 
                           => clk, RB => resetn, Q => in_buf_252_port);
   in_buf_reg_0_26 : DFERPQ1 port map( D => siso_data_in(10), CEB => n162, CK 
                           => clk, RB => resetn, Q => in_buf_250_port);
   in_buf_reg_0_24 : DFERPQ1 port map( D => siso_data_in(8), CEB => n162, CK =>
                           clk, RB => resetn, Q => in_buf_248_port);
   in_buf_reg_0_22 : DFERPQ1 port map( D => siso_data_in(6), CEB => n162, CK =>
                           clk, RB => resetn, Q => in_buf_246_port);
   in_buf_reg_0_20 : DFERPQ1 port map( D => siso_data_in(4), CEB => n162, CK =>
                           clk, RB => resetn, Q => in_buf_244_port);
   in_buf_reg_0_18 : DFERPQ1 port map( D => siso_data_in(2), CEB => n162, CK =>
                           clk, RB => resetn, Q => in_buf_242_port);
   in_buf_reg_0_16 : DFERPQ1 port map( D => siso_data_in(0), CEB => n162, CK =>
                           clk, RB => resetn, Q => in_buf_240_port);
   in_buf_reg_0_14 : DFERPQ1 port map( D => siso_data_in(14), CEB => n163, CK 
                           => clk, RB => resetn, Q => in_buf_238_port);
   in_buf_reg_0_12 : DFERPQ1 port map( D => siso_data_in(12), CEB => n163, CK 
                           => clk, RB => resetn, Q => in_buf_236_port);
   in_buf_reg_0_10 : DFERPQ1 port map( D => siso_data_in(10), CEB => n163, CK 
                           => clk, RB => resetn, Q => in_buf_234_port);
   in_buf_reg_0_8 : DFERPQ1 port map( D => siso_data_in(8), CEB => n163, CK => 
                           clk, RB => resetn, Q => in_buf_232_port);
   in_buf_reg_0_6 : DFERPQ1 port map( D => siso_data_in(6), CEB => n163, CK => 
                           clk, RB => resetn, Q => in_buf_230_port);
   in_buf_reg_0_4 : DFERPQ1 port map( D => siso_data_in(4), CEB => n163, CK => 
                           clk, RB => resetn, Q => in_buf_228_port);
   in_buf_reg_0_2 : DFERPQ1 port map( D => siso_data_in(2), CEB => n163, CK => 
                           clk, RB => resetn, Q => in_buf_226_port);
   in_buf_reg_4_14 : DFERPQ1 port map( D => siso_data_in(14), CEB => n171, CK 
                           => clk, RB => resetn, Q => in_buf_110_port);
   in_buf_reg_4_12 : DFERPQ1 port map( D => siso_data_in(12), CEB => n171, CK 
                           => clk, RB => resetn, Q => in_buf_108_port);
   in_buf_reg_4_10 : DFERPQ1 port map( D => siso_data_in(10), CEB => n171, CK 
                           => clk, RB => resetn, Q => in_buf_106_port);
   in_buf_reg_4_8 : DFERPQ1 port map( D => siso_data_in(8), CEB => n171, CK => 
                           clk, RB => resetn, Q => in_buf_104_port);
   in_buf_reg_4_6 : DFERPQ1 port map( D => siso_data_in(6), CEB => n171, CK => 
                           clk, RB => resetn, Q => in_buf_102_port);
   in_buf_reg_4_4 : DFERPQ1 port map( D => siso_data_in(4), CEB => n171, CK => 
                           clk, RB => resetn, Q => in_buf_100_port);
   in_buf_reg_4_2 : DFERPQ1 port map( D => siso_data_in(2), CEB => n171, CK => 
                           clk, RB => resetn, Q => in_buf_98_port);
   in_buf_reg_3_0 : DFERPQ1 port map( D => siso_data_in(0), CEB => n169, CK => 
                           clk, RB => resetn, Q => in_buf_128_port);
   in_buf_reg_2_0 : DFERPQ1 port map( D => siso_data_in(0), CEB => n167, CK => 
                           clk, RB => resetn, Q => in_buf_160_port);
   in_buf_reg_6_0 : DFERPQ1 port map( D => siso_data_in(0), CEB => n175, CK => 
                           clk, RB => resetn, Q => in_buf_32_port);
   in_buf_reg_5_0 : DFERPQ1 port map( D => siso_data_in(0), CEB => n173, CK => 
                           clk, RB => resetn, Q => in_buf_64_port);
   out_buf_reg_7_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => n245, CK
                           => clk, RB => resetn, Q => out_buf_15_port);
   out_buf_reg_7_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => n245, CK
                           => clk, RB => resetn, Q => out_buf_14_port);
   out_buf_reg_7_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => n245, CK
                           => clk, RB => resetn, Q => out_buf_13_port);
   out_buf_reg_7_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => n245, CK
                           => clk, RB => resetn, Q => out_buf_12_port);
   out_buf_reg_7_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => n245, CK
                           => clk, RB => resetn, Q => out_buf_11_port);
   out_buf_reg_7_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => n245, CK
                           => clk, RB => resetn, Q => out_buf_10_port);
   out_buf_reg_7_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n245, CK 
                           => clk, RB => resetn, Q => out_buf_9_port);
   out_buf_reg_7_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n245, CK 
                           => clk, RB => resetn, Q => out_buf_8_port);
   out_buf_reg_7_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n245, CK 
                           => clk, RB => resetn, Q => out_buf_7_port);
   out_buf_reg_7_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n245, CK 
                           => clk, RB => resetn, Q => out_buf_6_port);
   out_buf_reg_7_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n245, CK 
                           => clk, RB => resetn, Q => out_buf_5_port);
   out_buf_reg_7_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n245, CK 
                           => clk, RB => resetn, Q => out_buf_4_port);
   out_buf_reg_7_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n245, CK 
                           => clk, RB => resetn, Q => out_buf_3_port);
   out_buf_reg_7_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n245, CK 
                           => clk, RB => resetn, Q => out_buf_2_port);
   out_buf_reg_7_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n245, CK 
                           => clk, RB => resetn, Q => out_buf_1_port);
   out_buf_reg_7_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n245, CK 
                           => clk, RB => resetn, Q => out_buf_0_port);
   in_buf_reg_1_0 : DFERPQ1 port map( D => siso_data_in(0), CEB => n165, CK => 
                           clk, RB => resetn, Q => in_buf_192_port);
   out_buf_reg_3_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_143_port);
   out_buf_reg_3_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_142_port);
   out_buf_reg_3_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_141_port);
   out_buf_reg_3_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_140_port);
   out_buf_reg_3_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_139_port);
   out_buf_reg_3_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_138_port);
   out_buf_reg_3_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n252, CK 
                           => clk, RB => resetn, Q => out_buf_137_port);
   out_buf_reg_3_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n252, CK 
                           => clk, RB => resetn, Q => out_buf_136_port);
   out_buf_reg_3_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n252, CK 
                           => clk, RB => resetn, Q => out_buf_135_port);
   out_buf_reg_3_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n252, CK 
                           => clk, RB => resetn, Q => out_buf_134_port);
   out_buf_reg_3_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n252, CK 
                           => clk, RB => resetn, Q => out_buf_133_port);
   out_buf_reg_3_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n252, CK 
                           => clk, RB => resetn, Q => out_buf_132_port);
   out_buf_reg_3_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n252, CK 
                           => clk, RB => resetn, Q => out_buf_131_port);
   out_buf_reg_3_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n252, CK 
                           => clk, RB => resetn, Q => out_buf_130_port);
   out_buf_reg_3_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n252, CK 
                           => clk, RB => resetn, Q => out_buf_129_port);
   out_buf_reg_3_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n252, CK 
                           => clk, RB => resetn, Q => out_buf_128_port);
   in_buf_reg_0_0 : DFERPQ1 port map( D => siso_data_in(0), CEB => n163, CK => 
                           clk, RB => resetn, Q => in_buf_224_port);
   in_buf_reg_4_0 : DFERPQ1 port map( D => siso_data_in(0), CEB => n171, CK => 
                           clk, RB => resetn, Q => in_buf_96_port);
   out_buf_reg_2_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_175_port);
   out_buf_reg_2_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_174_port);
   out_buf_reg_2_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_173_port);
   out_buf_reg_2_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_172_port);
   out_buf_reg_2_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_171_port);
   out_buf_reg_2_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_170_port);
   out_buf_reg_2_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n251, CK 
                           => clk, RB => resetn, Q => out_buf_169_port);
   out_buf_reg_2_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n251, CK 
                           => clk, RB => resetn, Q => out_buf_168_port);
   out_buf_reg_2_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n251, CK 
                           => clk, RB => resetn, Q => out_buf_167_port);
   out_buf_reg_2_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n251, CK 
                           => clk, RB => resetn, Q => out_buf_166_port);
   out_buf_reg_2_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n251, CK 
                           => clk, RB => resetn, Q => out_buf_165_port);
   out_buf_reg_2_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n251, CK 
                           => clk, RB => resetn, Q => out_buf_164_port);
   out_buf_reg_2_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n251, CK 
                           => clk, RB => resetn, Q => out_buf_163_port);
   out_buf_reg_2_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n251, CK 
                           => clk, RB => resetn, Q => out_buf_162_port);
   out_buf_reg_2_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n251, CK 
                           => clk, RB => resetn, Q => out_buf_161_port);
   out_buf_reg_2_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n251, CK 
                           => clk, RB => resetn, Q => out_buf_160_port);
   out_buf_reg_6_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_47_port);
   out_buf_reg_6_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_46_port);
   out_buf_reg_6_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_45_port);
   out_buf_reg_6_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_44_port);
   out_buf_reg_6_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_43_port);
   out_buf_reg_6_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_42_port);
   out_buf_reg_6_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n250, CK 
                           => clk, RB => resetn, Q => out_buf_41_port);
   out_buf_reg_6_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n250, CK 
                           => clk, RB => resetn, Q => out_buf_40_port);
   out_buf_reg_6_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n250, CK 
                           => clk, RB => resetn, Q => out_buf_39_port);
   out_buf_reg_6_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n250, CK 
                           => clk, RB => resetn, Q => out_buf_38_port);
   out_buf_reg_6_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n250, CK 
                           => clk, RB => resetn, Q => out_buf_37_port);
   out_buf_reg_6_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n250, CK 
                           => clk, RB => resetn, Q => out_buf_36_port);
   out_buf_reg_6_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n250, CK 
                           => clk, RB => resetn, Q => out_buf_35_port);
   out_buf_reg_6_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n250, CK 
                           => clk, RB => resetn, Q => out_buf_34_port);
   out_buf_reg_6_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n250, CK 
                           => clk, RB => resetn, Q => out_buf_33_port);
   out_buf_reg_6_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n250, CK 
                           => clk, RB => resetn, Q => out_buf_32_port);
   out_buf_reg_7_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => n245, CK
                           => clk, RB => resetn, Q => out_buf_31_port);
   out_buf_reg_7_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => n245, CK
                           => clk, RB => resetn, Q => out_buf_30_port);
   out_buf_reg_7_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => n245, CK
                           => clk, RB => resetn, Q => out_buf_29_port);
   out_buf_reg_7_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => n245, CK
                           => clk, RB => resetn, Q => out_buf_28_port);
   out_buf_reg_7_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => n245, CK
                           => clk, RB => resetn, Q => out_buf_27_port);
   out_buf_reg_7_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => n245, CK
                           => clk, RB => resetn, Q => out_buf_26_port);
   out_buf_reg_7_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => n245, CK
                           => clk, RB => resetn, Q => out_buf_25_port);
   out_buf_reg_7_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => n245, CK
                           => clk, RB => resetn, Q => out_buf_24_port);
   out_buf_reg_7_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => n245, CK
                           => clk, RB => resetn, Q => out_buf_23_port);
   out_buf_reg_7_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => n245, CK
                           => clk, RB => resetn, Q => out_buf_22_port);
   out_buf_reg_7_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => n245, CK
                           => clk, RB => resetn, Q => out_buf_21_port);
   out_buf_reg_7_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => n245, CK
                           => clk, RB => resetn, Q => out_buf_20_port);
   out_buf_reg_7_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => n245, CK
                           => clk, RB => resetn, Q => out_buf_19_port);
   out_buf_reg_7_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => n245, CK
                           => clk, RB => resetn, Q => out_buf_18_port);
   out_buf_reg_7_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => n245, CK
                           => clk, RB => resetn, Q => out_buf_17_port);
   out_buf_reg_7_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => n245, CK
                           => clk, RB => resetn, Q => out_buf_16_port);
   out_buf_reg_5_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_79_port);
   out_buf_reg_5_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_78_port);
   out_buf_reg_5_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_77_port);
   out_buf_reg_5_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_76_port);
   out_buf_reg_5_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_75_port);
   out_buf_reg_5_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_74_port);
   out_buf_reg_5_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n249, CK 
                           => clk, RB => resetn, Q => out_buf_73_port);
   out_buf_reg_5_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n249, CK 
                           => clk, RB => resetn, Q => out_buf_72_port);
   out_buf_reg_5_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n249, CK 
                           => clk, RB => resetn, Q => out_buf_71_port);
   out_buf_reg_5_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n249, CK 
                           => clk, RB => resetn, Q => out_buf_70_port);
   out_buf_reg_5_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n249, CK 
                           => clk, RB => resetn, Q => out_buf_69_port);
   out_buf_reg_5_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n249, CK 
                           => clk, RB => resetn, Q => out_buf_68_port);
   out_buf_reg_5_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n249, CK 
                           => clk, RB => resetn, Q => out_buf_67_port);
   out_buf_reg_5_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n249, CK 
                           => clk, RB => resetn, Q => out_buf_66_port);
   out_buf_reg_5_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n249, CK 
                           => clk, RB => resetn, Q => out_buf_65_port);
   out_buf_reg_5_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n249, CK 
                           => clk, RB => resetn, Q => out_buf_64_port);
   out_buf_reg_3_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_159_port);
   out_buf_reg_3_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_158_port);
   out_buf_reg_3_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_157_port);
   out_buf_reg_3_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_156_port);
   out_buf_reg_3_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_155_port);
   out_buf_reg_3_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_154_port);
   out_buf_reg_3_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_153_port);
   out_buf_reg_3_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_152_port);
   out_buf_reg_3_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_151_port);
   out_buf_reg_3_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_150_port);
   out_buf_reg_3_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_149_port);
   out_buf_reg_3_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_148_port);
   out_buf_reg_3_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_147_port);
   out_buf_reg_3_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_146_port);
   out_buf_reg_3_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_145_port);
   out_buf_reg_3_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => n252, CK
                           => clk, RB => resetn, Q => out_buf_144_port);
   out_buf_reg_1_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_207_port);
   out_buf_reg_1_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_206_port);
   out_buf_reg_1_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_205_port);
   out_buf_reg_1_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_204_port);
   out_buf_reg_1_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_203_port);
   out_buf_reg_1_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_202_port);
   out_buf_reg_1_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n248, CK 
                           => clk, RB => resetn, Q => out_buf_201_port);
   out_buf_reg_1_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n248, CK 
                           => clk, RB => resetn, Q => out_buf_200_port);
   out_buf_reg_1_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n248, CK 
                           => clk, RB => resetn, Q => out_buf_199_port);
   out_buf_reg_1_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n248, CK 
                           => clk, RB => resetn, Q => out_buf_198_port);
   out_buf_reg_1_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n248, CK 
                           => clk, RB => resetn, Q => out_buf_197_port);
   out_buf_reg_1_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n248, CK 
                           => clk, RB => resetn, Q => out_buf_196_port);
   out_buf_reg_1_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n248, CK 
                           => clk, RB => resetn, Q => out_buf_195_port);
   out_buf_reg_1_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n248, CK 
                           => clk, RB => resetn, Q => out_buf_194_port);
   out_buf_reg_1_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n248, CK 
                           => clk, RB => resetn, Q => out_buf_193_port);
   out_buf_reg_1_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n248, CK 
                           => clk, RB => resetn, Q => out_buf_192_port);
   out_buf_reg_2_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_191_port);
   out_buf_reg_2_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_190_port);
   out_buf_reg_2_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_189_port);
   out_buf_reg_2_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_188_port);
   out_buf_reg_2_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_187_port);
   out_buf_reg_2_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_186_port);
   out_buf_reg_2_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_185_port);
   out_buf_reg_2_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_184_port);
   out_buf_reg_2_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_183_port);
   out_buf_reg_2_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_182_port);
   out_buf_reg_2_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_181_port);
   out_buf_reg_2_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_180_port);
   out_buf_reg_2_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_179_port);
   out_buf_reg_2_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_178_port);
   out_buf_reg_2_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_177_port);
   out_buf_reg_2_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => n251, CK
                           => clk, RB => resetn, Q => out_buf_176_port);
   out_buf_reg_6_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_63_port);
   out_buf_reg_6_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_62_port);
   out_buf_reg_6_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_61_port);
   out_buf_reg_6_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_60_port);
   out_buf_reg_6_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_59_port);
   out_buf_reg_6_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_58_port);
   out_buf_reg_6_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_57_port);
   out_buf_reg_6_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_56_port);
   out_buf_reg_6_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_55_port);
   out_buf_reg_6_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_54_port);
   out_buf_reg_6_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_53_port);
   out_buf_reg_6_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_52_port);
   out_buf_reg_6_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_51_port);
   out_buf_reg_6_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_50_port);
   out_buf_reg_6_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_49_port);
   out_buf_reg_6_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => n250, CK
                           => clk, RB => resetn, Q => out_buf_48_port);
   out_buf_reg_0_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_239_port);
   out_buf_reg_0_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_238_port);
   out_buf_reg_0_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_237_port);
   out_buf_reg_0_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_236_port);
   out_buf_reg_0_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_235_port);
   out_buf_reg_0_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_234_port);
   out_buf_reg_0_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n247, CK 
                           => clk, RB => resetn, Q => out_buf_233_port);
   out_buf_reg_0_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n247, CK 
                           => clk, RB => resetn, Q => out_buf_232_port);
   out_buf_reg_0_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n247, CK 
                           => clk, RB => resetn, Q => out_buf_231_port);
   out_buf_reg_0_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n247, CK 
                           => clk, RB => resetn, Q => out_buf_230_port);
   out_buf_reg_0_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n247, CK 
                           => clk, RB => resetn, Q => out_buf_229_port);
   out_buf_reg_0_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n247, CK 
                           => clk, RB => resetn, Q => out_buf_228_port);
   out_buf_reg_0_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n247, CK 
                           => clk, RB => resetn, Q => out_buf_227_port);
   out_buf_reg_0_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n247, CK 
                           => clk, RB => resetn, Q => out_buf_226_port);
   out_buf_reg_0_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n247, CK 
                           => clk, RB => resetn, Q => out_buf_225_port);
   out_buf_reg_0_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n247, CK 
                           => clk, RB => resetn, Q => out_buf_224_port);
   out_buf_reg_4_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_111_port);
   out_buf_reg_4_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_110_port);
   out_buf_reg_4_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_109_port);
   out_buf_reg_4_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_108_port);
   out_buf_reg_4_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_107_port);
   out_buf_reg_4_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_106_port);
   out_buf_reg_4_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n246, CK 
                           => clk, RB => resetn, Q => out_buf_105_port);
   out_buf_reg_4_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n246, CK 
                           => clk, RB => resetn, Q => out_buf_104_port);
   out_buf_reg_4_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n246, CK 
                           => clk, RB => resetn, Q => out_buf_103_port);
   out_buf_reg_4_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n246, CK 
                           => clk, RB => resetn, Q => out_buf_102_port);
   out_buf_reg_4_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n246, CK 
                           => clk, RB => resetn, Q => out_buf_101_port);
   out_buf_reg_4_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n246, CK 
                           => clk, RB => resetn, Q => out_buf_100_port);
   out_buf_reg_4_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n246, CK 
                           => clk, RB => resetn, Q => out_buf_99_port);
   out_buf_reg_4_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n246, CK 
                           => clk, RB => resetn, Q => out_buf_98_port);
   out_buf_reg_4_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n246, CK 
                           => clk, RB => resetn, Q => out_buf_97_port);
   out_buf_reg_4_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n246, CK 
                           => clk, RB => resetn, Q => out_buf_96_port);
   out_buf_reg_5_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_95_port);
   out_buf_reg_5_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_94_port);
   out_buf_reg_5_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_93_port);
   out_buf_reg_5_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_92_port);
   out_buf_reg_5_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_91_port);
   out_buf_reg_5_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_90_port);
   out_buf_reg_5_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_89_port);
   out_buf_reg_5_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_88_port);
   out_buf_reg_5_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_87_port);
   out_buf_reg_5_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_86_port);
   out_buf_reg_5_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_85_port);
   out_buf_reg_5_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_84_port);
   out_buf_reg_5_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_83_port);
   out_buf_reg_5_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_82_port);
   out_buf_reg_5_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_81_port);
   out_buf_reg_5_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => n249, CK
                           => clk, RB => resetn, Q => out_buf_80_port);
   out_buf_reg_1_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_223_port);
   out_buf_reg_1_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_222_port);
   out_buf_reg_1_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_221_port);
   out_buf_reg_1_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_220_port);
   out_buf_reg_1_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_219_port);
   out_buf_reg_1_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_218_port);
   out_buf_reg_1_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_217_port);
   out_buf_reg_1_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_216_port);
   out_buf_reg_1_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_215_port);
   out_buf_reg_1_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_214_port);
   out_buf_reg_1_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_213_port);
   out_buf_reg_1_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_212_port);
   out_buf_reg_1_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_211_port);
   out_buf_reg_1_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_210_port);
   out_buf_reg_1_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_209_port);
   out_buf_reg_1_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => n248, CK
                           => clk, RB => resetn, Q => out_buf_208_port);
   out_buf_reg_0_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_255_port);
   out_buf_reg_0_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_254_port);
   out_buf_reg_0_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_253_port);
   out_buf_reg_0_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_252_port);
   out_buf_reg_0_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_251_port);
   out_buf_reg_0_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_250_port);
   out_buf_reg_0_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_249_port);
   out_buf_reg_0_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_248_port);
   out_buf_reg_0_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_247_port);
   out_buf_reg_0_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_246_port);
   out_buf_reg_0_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_245_port);
   out_buf_reg_0_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_244_port);
   out_buf_reg_0_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_243_port);
   out_buf_reg_0_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_242_port);
   out_buf_reg_0_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_241_port);
   out_buf_reg_0_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => n247, CK
                           => clk, RB => resetn, Q => out_buf_240_port);
   out_buf_reg_4_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_127_port);
   out_buf_reg_4_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_126_port);
   out_buf_reg_4_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_125_port);
   out_buf_reg_4_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_124_port);
   out_buf_reg_4_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_123_port);
   out_buf_reg_4_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_122_port);
   out_buf_reg_4_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_121_port);
   out_buf_reg_4_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_120_port);
   out_buf_reg_4_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_119_port);
   out_buf_reg_4_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_118_port);
   out_buf_reg_4_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_117_port);
   out_buf_reg_4_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_116_port);
   out_buf_reg_4_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_115_port);
   out_buf_reg_4_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_114_port);
   out_buf_reg_4_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_113_port);
   out_buf_reg_4_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => n246, CK
                           => clk, RB => resetn, Q => out_buf_112_port);
   out_trigger_reg : DFFRPQ1 port map( D => n240, CK => clk, RB => resetn, Q =>
                           out_trigger);
   read_comp_res_reg : DFERPQ1 port map( D => avs_writedata(2), CEB => n179, CK
                           => clk, RB => resetn, Q => read_comp_res);
   in_counter_reg_0 : DFERPQ1 port map( D => n155, CEB => n683, CK => clk, RB 
                           => resetn, Q => in_counter_0_port);
   in_counter_reg_2 : DFFRPQ1 port map( D => n238, CK => clk, RB => resetn, Q 
                           => in_counter_2_port);
   in_counter_reg_1 : DFFRPQ1 port map( D => n237, CK => clk, RB => resetn, Q 
                           => in_counter_1_port);
   in_busy_reg : DFFRPQ1 port map( D => n239, CK => clk, RB => resetn, Q => 
                           in_busy);
   odd_reg : DFFRPQ1 port map( D => n156, CK => clk, RB => resetn, Q => odd);
   out_busy_reg : DFFRPQ1 port map( D => n234, CK => clk, RB => resetn, Q => 
                           out_busy);
   odd_reg2 : DFFRPQ1 port map( D => n154, CK => clk, RB => resetn, Q => odd1);
   operand_load_reg : DFERPQ1 port map( D => avs_writedata(1), CEB => n179, CK 
                           => clk, RB => resetn, Q => operand_load);
   coeff_load_reg : DFERPQ1 port map( D => avs_writedata(0), CEB => n179, CK =>
                           clk, RB => resetn, Q => coeff_load);
   out_counter_reg_0 : DFFRPQ1 port map( D => n236, CK => clk, RB => resetn, Q 
                           => N62);
   out_counter_reg_2 : DFFRPQ1 port map( D => n235, CK => clk, RB => resetn, Q 
                           => N64);
   out_counter_reg_1 : DFFRPQ1 port map( D => n201, CK => clk, RB => resetn, Q 
                           => N63);
   operand_regs_reg_3_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_159_port);
   operand_regs_reg_5_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_95_port);
   operand_regs_reg_1_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_223_port);
   coeff_memory_reg_1_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_31);
   coeff_memory_reg_2_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_31);
   coeff_memory_reg_3_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_31);
   coeff_memory_reg_0_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_31);
   coeff_memory_reg_4_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_31);
   operand_regs_reg_2_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_191_port);
   operand_regs_reg_4_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_127_port);
   operand_regs_reg_6_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_63_port);
   operand_regs_reg_7_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_31_port);
   operand_regs_reg_3_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_158_port);
   operand_regs_reg_5_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_94_port);
   operand_regs_reg_0_31 : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_255_port);
   operand_regs_reg_3_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_157_port);
   operand_regs_reg_5_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_93_port);
   coeff_memory_reg_1_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_30);
   coeff_memory_reg_2_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_30);
   coeff_memory_reg_3_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_30);
   coeff_memory_reg_0_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_30);
   coeff_memory_reg_4_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_30);
   operand_regs_reg_2_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_190_port);
   operand_regs_reg_4_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_126_port);
   operand_regs_reg_6_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_62_port);
   operand_regs_reg_1_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_222_port);
   operand_regs_reg_7_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_30_port);
   operand_regs_reg_0_30 : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_254_port);
   operand_regs_reg_1_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_221_port);
   operand_regs_reg_3_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_156_port);
   operand_regs_reg_5_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_92_port);
   operand_regs_reg_1_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_220_port);
   coeff_memory_reg_1_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_29);
   coeff_memory_reg_2_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_29);
   coeff_memory_reg_3_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_29);
   operand_regs_reg_3_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_155_port);
   operand_regs_reg_5_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_91_port);
   coeff_memory_reg_0_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_29);
   coeff_memory_reg_4_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_29);
   operand_regs_reg_2_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_189_port);
   operand_regs_reg_4_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_125_port);
   operand_regs_reg_6_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_61_port);
   operand_regs_reg_7_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_29_port);
   operand_regs_reg_0_29 : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_253_port);
   coeff_memory_reg_1_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_28);
   coeff_memory_reg_2_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_28);
   coeff_memory_reg_3_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_28);
   coeff_memory_reg_0_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_28);
   coeff_memory_reg_4_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_28);
   operand_regs_reg_2_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_188_port);
   operand_regs_reg_4_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_124_port);
   operand_regs_reg_6_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_60_port);
   operand_regs_reg_7_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_28_port);
   operand_regs_reg_0_28 : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_252_port);
   operand_regs_reg_1_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_219_port);
   coeff_memory_reg_1_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_27);
   coeff_memory_reg_2_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_27);
   coeff_memory_reg_3_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_27);
   operand_regs_reg_3_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_154_port);
   operand_regs_reg_5_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_90_port);
   coeff_memory_reg_0_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_27);
   coeff_memory_reg_4_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_27);
   operand_regs_reg_2_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_187_port);
   operand_regs_reg_4_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_123_port);
   operand_regs_reg_6_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_59_port);
   operand_regs_reg_7_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_27_port);
   operand_regs_reg_0_27 : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_251_port);
   coeff_memory_reg_1_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_26);
   coeff_memory_reg_2_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_26);
   coeff_memory_reg_3_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_26);
   coeff_memory_reg_0_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_26);
   coeff_memory_reg_4_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_26);
   operand_regs_reg_2_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_186_port);
   operand_regs_reg_4_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_122_port);
   operand_regs_reg_6_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_58_port);
   operand_regs_reg_7_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_26_port);
   operand_regs_reg_1_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_218_port);
   operand_regs_reg_0_26 : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_250_port);
   operand_regs_reg_3_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_153_port);
   operand_regs_reg_5_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_89_port);
   operand_regs_reg_1_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_217_port);
   coeff_memory_reg_1_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_25);
   coeff_memory_reg_2_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_25);
   coeff_memory_reg_3_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_25);
   coeff_memory_reg_0_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_25);
   coeff_memory_reg_4_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_25);
   operand_regs_reg_2_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_185_port);
   operand_regs_reg_4_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_121_port);
   operand_regs_reg_6_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_57_port);
   operand_regs_reg_7_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_25_port);
   operand_regs_reg_0_25 : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_249_port);
   operand_regs_reg_3_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_152_port);
   operand_regs_reg_5_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_88_port);
   coeff_memory_reg_1_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_24);
   coeff_memory_reg_2_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_24);
   coeff_memory_reg_3_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_24);
   coeff_memory_reg_0_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_24);
   coeff_memory_reg_4_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_24);
   operand_regs_reg_2_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_184_port);
   operand_regs_reg_4_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_120_port);
   operand_regs_reg_6_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_56_port);
   operand_regs_reg_0_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_248_port);
   operand_regs_reg_7_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_24_port);
   operand_regs_reg_1_24 : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_216_port);
   operand_regs_reg_3_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_151_port);
   operand_regs_reg_5_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_87_port);
   operand_regs_reg_1_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_215_port);
   coeff_memory_reg_1_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_23);
   coeff_memory_reg_2_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_23);
   coeff_memory_reg_3_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_23);
   coeff_memory_reg_0_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_23);
   coeff_memory_reg_4_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_23);
   operand_regs_reg_2_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_183_port);
   operand_regs_reg_4_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_119_port);
   operand_regs_reg_6_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_55_port);
   operand_regs_reg_7_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_23_port);
   operand_regs_reg_0_23 : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_247_port);
   operand_regs_reg_3_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_150_port);
   operand_regs_reg_5_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_86_port);
   operand_regs_reg_3_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_149_port);
   operand_regs_reg_5_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_85_port);
   coeff_memory_reg_1_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_22);
   coeff_memory_reg_2_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_22);
   coeff_memory_reg_3_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_22);
   coeff_memory_reg_0_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_22);
   coeff_memory_reg_4_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_22);
   operand_regs_reg_2_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_182_port);
   operand_regs_reg_4_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_118_port);
   operand_regs_reg_6_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_54_port);
   operand_regs_reg_0_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_246_port);
   operand_regs_reg_7_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_22_port);
   operand_regs_reg_1_22 : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_214_port);
   operand_regs_reg_1_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_213_port);
   coeff_memory_reg_1_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_21);
   coeff_memory_reg_2_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_21);
   coeff_memory_reg_3_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_21);
   operand_regs_reg_3_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_148_port);
   operand_regs_reg_5_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_84_port);
   operand_regs_reg_3_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_147_port);
   operand_regs_reg_5_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_83_port);
   coeff_memory_reg_0_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_21);
   coeff_memory_reg_4_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_21);
   operand_regs_reg_2_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_181_port);
   operand_regs_reg_4_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_117_port);
   operand_regs_reg_6_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_53_port);
   operand_regs_reg_7_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_21_port);
   operand_regs_reg_0_21 : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_245_port);
   coeff_memory_reg_1_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_20);
   coeff_memory_reg_2_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_20);
   coeff_memory_reg_3_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_20);
   coeff_memory_reg_0_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_20);
   coeff_memory_reg_4_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_20);
   operand_regs_reg_2_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_180_port);
   operand_regs_reg_4_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_116_port);
   operand_regs_reg_6_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_52_port);
   operand_regs_reg_0_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_244_port);
   operand_regs_reg_7_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_20_port);
   operand_regs_reg_1_20 : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_212_port);
   operand_regs_reg_1_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_211_port);
   operand_regs_reg_5_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_82_port);
   operand_regs_reg_3_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_146_port);
   operand_regs_reg_3_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_145_port);
   operand_regs_reg_5_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_81_port);
   operand_regs_reg_1_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_210_port);
   coeff_memory_reg_1_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_19);
   coeff_memory_reg_2_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_19);
   coeff_memory_reg_3_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_19);
   coeff_memory_reg_0_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_19);
   coeff_memory_reg_4_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_19);
   operand_regs_reg_2_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_179_port);
   operand_regs_reg_4_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_115_port);
   operand_regs_reg_6_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_51_port);
   operand_regs_reg_7_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_19_port);
   operand_regs_reg_0_19 : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_243_port);
   operand_regs_reg_1_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_209_port);
   coeff_memory_reg_1_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_18);
   coeff_memory_reg_2_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_18);
   coeff_memory_reg_3_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_18);
   coeff_memory_reg_0_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_18);
   coeff_memory_reg_4_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_18);
   operand_regs_reg_2_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_178_port);
   operand_regs_reg_4_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_114_port);
   operand_regs_reg_6_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_50_port);
   operand_regs_reg_7_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_18_port);
   operand_regs_reg_0_18 : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_242_port);
   operand_regs_reg_3_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_144_port);
   operand_regs_reg_5_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_80_port);
   coeff_memory_reg_1_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_17);
   coeff_memory_reg_2_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_17);
   coeff_memory_reg_3_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_17);
   coeff_memory_reg_0_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_17);
   coeff_memory_reg_4_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_17);
   operand_regs_reg_2_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_177_port);
   operand_regs_reg_4_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_113_port);
   operand_regs_reg_6_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_49_port);
   operand_regs_reg_7_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_17_port);
   operand_regs_reg_0_17 : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_241_port);
   coeff_memory_reg_1_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_16);
   coeff_memory_reg_2_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_16);
   coeff_memory_reg_3_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_16);
   coeff_memory_reg_0_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_16);
   coeff_memory_reg_4_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_16);
   operand_regs_reg_2_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_176_port);
   operand_regs_reg_4_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_112_port);
   operand_regs_reg_6_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_48_port);
   operand_regs_reg_7_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_16_port);
   operand_regs_reg_0_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_240_port);
   operand_regs_reg_1_16 : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_208_port);
   operand_regs_reg_3_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_143_port);
   operand_regs_reg_5_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_79_port);
   coeff_memory_reg_1_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_15);
   coeff_memory_reg_2_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_15);
   coeff_memory_reg_3_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_15);
   coeff_memory_reg_0_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_15);
   coeff_memory_reg_4_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_15);
   operand_regs_reg_2_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_175_port);
   operand_regs_reg_4_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_111_port);
   operand_regs_reg_6_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_47_port);
   operand_regs_reg_0_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_239_port);
   operand_regs_reg_3_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_142_port);
   operand_regs_reg_5_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_78_port);
   operand_regs_reg_7_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_15_port);
   operand_regs_reg_3_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_141_port);
   operand_regs_reg_5_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_77_port);
   operand_regs_reg_1_15 : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_207_port);
   coeff_memory_reg_1_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_14);
   coeff_memory_reg_2_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_14);
   coeff_memory_reg_3_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_14);
   coeff_memory_reg_0_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_14);
   coeff_memory_reg_4_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_14);
   operand_regs_reg_2_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_174_port);
   operand_regs_reg_4_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_110_port);
   operand_regs_reg_6_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_46_port);
   operand_regs_reg_0_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_238_port);
   operand_regs_reg_7_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_14_port);
   operand_regs_reg_1_14 : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_206_port);
   operand_regs_reg_1_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_205_port);
   coeff_memory_reg_1_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_13);
   coeff_memory_reg_2_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_13);
   coeff_memory_reg_3_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_13);
   coeff_memory_reg_0_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_13);
   coeff_memory_reg_4_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_13);
   operand_regs_reg_2_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_173_port);
   operand_regs_reg_4_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_109_port);
   operand_regs_reg_6_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_45_port);
   operand_regs_reg_7_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_13_port);
   operand_regs_reg_0_13 : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_237_port);
   operand_regs_reg_3_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_140_port);
   operand_regs_reg_5_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_76_port);
   operand_regs_reg_3_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_139_port);
   operand_regs_reg_5_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_75_port);
   coeff_memory_reg_1_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_12);
   coeff_memory_reg_2_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_12);
   coeff_memory_reg_3_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_12);
   coeff_memory_reg_0_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_12);
   coeff_memory_reg_4_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_12);
   operand_regs_reg_2_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_172_port);
   operand_regs_reg_4_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_108_port);
   operand_regs_reg_6_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_44_port);
   operand_regs_reg_0_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_236_port);
   operand_regs_reg_3_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_138_port);
   operand_regs_reg_5_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_74_port);
   operand_regs_reg_7_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_12_port);
   operand_regs_reg_1_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_203_port);
   operand_regs_reg_1_12 : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_204_port);
   coeff_memory_reg_1_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_11);
   coeff_memory_reg_2_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_11);
   coeff_memory_reg_3_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_11);
   coeff_memory_reg_0_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_11);
   coeff_memory_reg_4_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_11);
   operand_regs_reg_2_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_171_port);
   operand_regs_reg_4_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_107_port);
   operand_regs_reg_6_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_43_port);
   operand_regs_reg_7_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_11_port);
   operand_regs_reg_0_11 : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_235_port);
   operand_regs_reg_3_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n255,
                           CK => clk, RB => resetn, Q => operand_regs_137_port)
                           ;
   operand_regs_reg_5_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n260,
                           CK => clk, RB => resetn, Q => operand_regs_73_port);
   coeff_memory_reg_1_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_10);
   coeff_memory_reg_2_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n262, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_10);
   coeff_memory_reg_3_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_10);
   coeff_memory_reg_0_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_10);
   coeff_memory_reg_4_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_10);
   operand_regs_reg_2_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n254, CK => clk, RB => resetn, Q => 
                           operand_regs_170_port);
   operand_regs_reg_4_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_106_port);
   operand_regs_reg_6_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_42_port);
   operand_regs_reg_7_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n253, CK => clk, RB => resetn, Q => 
                           operand_regs_10_port);
   operand_regs_reg_1_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_202_port);
   operand_regs_reg_0_10 : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_234_port);
   coeff_memory_reg_1_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n264,
                           CK => clk, RB => resetn, Q => coeff_memory_1_9);
   coeff_memory_reg_2_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n262,
                           CK => clk, RB => resetn, Q => coeff_memory_2_9);
   coeff_memory_reg_3_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n261,
                           CK => clk, RB => resetn, Q => coeff_memory_3_9);
   operand_regs_reg_1_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n257,
                           CK => clk, RB => resetn, Q => operand_regs_201_port)
                           ;
   coeff_memory_reg_0_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n263,
                           CK => clk, RB => resetn, Q => coeff_memory_0_9);
   coeff_memory_reg_4_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n265,
                           CK => clk, RB => resetn, Q => coeff_memory_4_9);
   operand_regs_reg_2_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n254,
                           CK => clk, RB => resetn, Q => operand_regs_169_port)
                           ;
   operand_regs_reg_4_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n258,
                           CK => clk, RB => resetn, Q => operand_regs_105_port)
                           ;
   operand_regs_reg_6_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n259,
                           CK => clk, RB => resetn, Q => operand_regs_41_port);
   operand_regs_reg_7_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n253,
                           CK => clk, RB => resetn, Q => operand_regs_9_port);
   operand_regs_reg_0_9 : DFERPQ1 port map( D => avs_writedata(9), CEB => n256,
                           CK => clk, RB => resetn, Q => operand_regs_233_port)
                           ;
   operand_regs_reg_3_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n255,
                           CK => clk, RB => resetn, Q => operand_regs_135_port)
                           ;
   operand_regs_reg_5_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n260,
                           CK => clk, RB => resetn, Q => operand_regs_71_port);
   operand_regs_reg_3_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n255,
                           CK => clk, RB => resetn, Q => operand_regs_136_port)
                           ;
   operand_regs_reg_5_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n260,
                           CK => clk, RB => resetn, Q => operand_regs_72_port);
   coeff_memory_reg_1_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n264,
                           CK => clk, RB => resetn, Q => coeff_memory_1_8);
   coeff_memory_reg_2_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n262,
                           CK => clk, RB => resetn, Q => coeff_memory_2_8);
   coeff_memory_reg_3_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n261,
                           CK => clk, RB => resetn, Q => coeff_memory_3_8);
   coeff_memory_reg_0_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n263,
                           CK => clk, RB => resetn, Q => coeff_memory_0_8);
   coeff_memory_reg_4_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n265,
                           CK => clk, RB => resetn, Q => coeff_memory_4_8);
   operand_regs_reg_2_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n254,
                           CK => clk, RB => resetn, Q => operand_regs_168_port)
                           ;
   operand_regs_reg_4_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n258,
                           CK => clk, RB => resetn, Q => operand_regs_104_port)
                           ;
   operand_regs_reg_6_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n259,
                           CK => clk, RB => resetn, Q => operand_regs_40_port);
   operand_regs_reg_0_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n256,
                           CK => clk, RB => resetn, Q => operand_regs_232_port)
                           ;
   operand_regs_reg_7_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n253,
                           CK => clk, RB => resetn, Q => operand_regs_8_port);
   operand_regs_reg_3_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n255,
                           CK => clk, RB => resetn, Q => operand_regs_134_port)
                           ;
   operand_regs_reg_5_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n260,
                           CK => clk, RB => resetn, Q => operand_regs_70_port);
   operand_regs_reg_1_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n257,
                           CK => clk, RB => resetn, Q => operand_regs_199_port)
                           ;
   operand_regs_reg_1_8 : DFERPQ1 port map( D => avs_writedata(8), CEB => n257,
                           CK => clk, RB => resetn, Q => operand_regs_200_port)
                           ;
   operand_regs_reg_1_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n257,
                           CK => clk, RB => resetn, Q => operand_regs_198_port)
                           ;
   coeff_memory_reg_1_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n264,
                           CK => clk, RB => resetn, Q => coeff_memory_1_7);
   coeff_memory_reg_2_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n262,
                           CK => clk, RB => resetn, Q => coeff_memory_2_7);
   coeff_memory_reg_3_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n261,
                           CK => clk, RB => resetn, Q => coeff_memory_3_7);
   operand_regs_reg_3_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n255,
                           CK => clk, RB => resetn, Q => operand_regs_133_port)
                           ;
   operand_regs_reg_5_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n260,
                           CK => clk, RB => resetn, Q => operand_regs_69_port);
   coeff_memory_reg_0_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n263,
                           CK => clk, RB => resetn, Q => coeff_memory_0_7);
   coeff_memory_reg_4_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n265,
                           CK => clk, RB => resetn, Q => coeff_memory_4_7);
   operand_regs_reg_2_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n254,
                           CK => clk, RB => resetn, Q => operand_regs_167_port)
                           ;
   operand_regs_reg_4_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n258,
                           CK => clk, RB => resetn, Q => operand_regs_103_port)
                           ;
   operand_regs_reg_6_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n259,
                           CK => clk, RB => resetn, Q => operand_regs_39_port);
   operand_regs_reg_7_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n253,
                           CK => clk, RB => resetn, Q => operand_regs_7_port);
   operand_regs_reg_0_7 : DFERPQ1 port map( D => avs_writedata(7), CEB => n256,
                           CK => clk, RB => resetn, Q => operand_regs_231_port)
                           ;
   operand_regs_reg_1_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n257,
                           CK => clk, RB => resetn, Q => operand_regs_197_port)
                           ;
   coeff_memory_reg_1_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n264,
                           CK => clk, RB => resetn, Q => coeff_memory_1_6);
   coeff_memory_reg_2_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n262,
                           CK => clk, RB => resetn, Q => coeff_memory_2_6);
   coeff_memory_reg_3_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n261,
                           CK => clk, RB => resetn, Q => coeff_memory_3_6);
   coeff_memory_reg_0_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n263,
                           CK => clk, RB => resetn, Q => coeff_memory_0_6);
   coeff_memory_reg_4_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n265,
                           CK => clk, RB => resetn, Q => coeff_memory_4_6);
   operand_regs_reg_2_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n254,
                           CK => clk, RB => resetn, Q => operand_regs_166_port)
                           ;
   operand_regs_reg_4_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n258,
                           CK => clk, RB => resetn, Q => operand_regs_102_port)
                           ;
   operand_regs_reg_6_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n259,
                           CK => clk, RB => resetn, Q => operand_regs_38_port);
   operand_regs_reg_7_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n253,
                           CK => clk, RB => resetn, Q => operand_regs_6_port);
   operand_regs_reg_0_6 : DFERPQ1 port map( D => avs_writedata(6), CEB => n256,
                           CK => clk, RB => resetn, Q => operand_regs_230_port)
                           ;
   coeff_memory_reg_1_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n264,
                           CK => clk, RB => resetn, Q => coeff_memory_1_5);
   coeff_memory_reg_2_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n262,
                           CK => clk, RB => resetn, Q => coeff_memory_2_5);
   coeff_memory_reg_3_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n261,
                           CK => clk, RB => resetn, Q => coeff_memory_3_5);
   coeff_memory_reg_0_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n263,
                           CK => clk, RB => resetn, Q => coeff_memory_0_5);
   coeff_memory_reg_4_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n265,
                           CK => clk, RB => resetn, Q => coeff_memory_4_5);
   operand_regs_reg_2_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n254,
                           CK => clk, RB => resetn, Q => operand_regs_165_port)
                           ;
   operand_regs_reg_4_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n258,
                           CK => clk, RB => resetn, Q => operand_regs_101_port)
                           ;
   operand_regs_reg_6_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n259,
                           CK => clk, RB => resetn, Q => operand_regs_37_port);
   operand_regs_reg_7_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n253,
                           CK => clk, RB => resetn, Q => operand_regs_5_port);
   operand_regs_reg_0_5 : DFERPQ1 port map( D => avs_writedata(5), CEB => n256,
                           CK => clk, RB => resetn, Q => operand_regs_229_port)
                           ;
   operand_regs_reg_3_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n255,
                           CK => clk, RB => resetn, Q => operand_regs_132_port)
                           ;
   operand_regs_reg_5_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n260,
                           CK => clk, RB => resetn, Q => operand_regs_68_port);
   operand_regs_reg_3_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n255,
                           CK => clk, RB => resetn, Q => operand_regs_131_port)
                           ;
   operand_regs_reg_5_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n260,
                           CK => clk, RB => resetn, Q => operand_regs_67_port);
   coeff_memory_reg_1_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n264,
                           CK => clk, RB => resetn, Q => coeff_memory_1_4);
   coeff_memory_reg_2_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n262,
                           CK => clk, RB => resetn, Q => coeff_memory_2_4);
   coeff_memory_reg_3_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n261,
                           CK => clk, RB => resetn, Q => coeff_memory_3_4);
   coeff_memory_reg_0_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n263,
                           CK => clk, RB => resetn, Q => coeff_memory_0_4);
   coeff_memory_reg_4_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n265,
                           CK => clk, RB => resetn, Q => coeff_memory_4_4);
   operand_regs_reg_2_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n254,
                           CK => clk, RB => resetn, Q => operand_regs_164_port)
                           ;
   operand_regs_reg_4_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n258,
                           CK => clk, RB => resetn, Q => operand_regs_100_port)
                           ;
   operand_regs_reg_6_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n259,
                           CK => clk, RB => resetn, Q => operand_regs_36_port);
   operand_regs_reg_7_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n253,
                           CK => clk, RB => resetn, Q => operand_regs_4_port);
   operand_regs_reg_0_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n256,
                           CK => clk, RB => resetn, Q => operand_regs_228_port)
                           ;
   operand_regs_reg_1_4 : DFERPQ1 port map( D => avs_writedata(4), CEB => n257,
                           CK => clk, RB => resetn, Q => operand_regs_196_port)
                           ;
   operand_regs_reg_1_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n257,
                           CK => clk, RB => resetn, Q => operand_regs_195_port)
                           ;
   coeff_memory_reg_1_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n264,
                           CK => clk, RB => resetn, Q => coeff_memory_1_3);
   coeff_memory_reg_2_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n262,
                           CK => clk, RB => resetn, Q => coeff_memory_2_3);
   coeff_memory_reg_3_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n261,
                           CK => clk, RB => resetn, Q => coeff_memory_3_3);
   coeff_memory_reg_0_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n263,
                           CK => clk, RB => resetn, Q => coeff_memory_0_3);
   coeff_memory_reg_4_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n265,
                           CK => clk, RB => resetn, Q => coeff_memory_4_3);
   operand_regs_reg_2_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n254,
                           CK => clk, RB => resetn, Q => operand_regs_163_port)
                           ;
   operand_regs_reg_4_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n258,
                           CK => clk, RB => resetn, Q => operand_regs_99_port);
   operand_regs_reg_6_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n259,
                           CK => clk, RB => resetn, Q => operand_regs_35_port);
   operand_regs_reg_7_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n253,
                           CK => clk, RB => resetn, Q => operand_regs_3_port);
   operand_regs_reg_3_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n255,
                           CK => clk, RB => resetn, Q => operand_regs_128_port)
                           ;
   operand_regs_reg_5_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n260,
                           CK => clk, RB => resetn, Q => operand_regs_64_port);
   operand_regs_reg_0_3 : DFERPQ1 port map( D => avs_writedata(3), CEB => n256,
                           CK => clk, RB => resetn, Q => operand_regs_227_port)
                           ;
   coeff_memory_reg_1_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n264,
                           CK => clk, RB => resetn, Q => coeff_memory_1_2);
   coeff_memory_reg_2_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n262,
                           CK => clk, RB => resetn, Q => coeff_memory_2_2);
   coeff_memory_reg_3_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n261,
                           CK => clk, RB => resetn, Q => coeff_memory_3_2);
   coeff_memory_reg_0_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n263,
                           CK => clk, RB => resetn, Q => coeff_memory_0_2);
   coeff_memory_reg_4_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n265,
                           CK => clk, RB => resetn, Q => coeff_memory_4_2);
   operand_regs_reg_2_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n254,
                           CK => clk, RB => resetn, Q => operand_regs_162_port)
                           ;
   operand_regs_reg_4_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n258,
                           CK => clk, RB => resetn, Q => operand_regs_98_port);
   operand_regs_reg_6_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n259,
                           CK => clk, RB => resetn, Q => operand_regs_34_port);
   operand_regs_reg_3_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n255,
                           CK => clk, RB => resetn, Q => operand_regs_129_port)
                           ;
   operand_regs_reg_5_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n260,
                           CK => clk, RB => resetn, Q => operand_regs_65_port);
   operand_regs_reg_3_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n255,
                           CK => clk, RB => resetn, Q => operand_regs_130_port)
                           ;
   operand_regs_reg_5_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n260,
                           CK => clk, RB => resetn, Q => operand_regs_66_port);
   operand_regs_reg_1_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n257,
                           CK => clk, RB => resetn, Q => operand_regs_192_port)
                           ;
   operand_regs_reg_0_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n256,
                           CK => clk, RB => resetn, Q => operand_regs_226_port)
                           ;
   operand_regs_reg_7_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n253,
                           CK => clk, RB => resetn, Q => operand_regs_2_port);
   operand_regs_reg_1_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n257,
                           CK => clk, RB => resetn, Q => operand_regs_193_port)
                           ;
   operand_regs_reg_1_2 : DFERPQ1 port map( D => avs_writedata(2), CEB => n257,
                           CK => clk, RB => resetn, Q => operand_regs_194_port)
                           ;
   coeff_memory_reg_1_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n264,
                           CK => clk, RB => resetn, Q => coeff_memory_1_1);
   coeff_memory_reg_2_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n262,
                           CK => clk, RB => resetn, Q => coeff_memory_2_1);
   coeff_memory_reg_3_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n261,
                           CK => clk, RB => resetn, Q => coeff_memory_3_1);
   coeff_memory_reg_0_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n263,
                           CK => clk, RB => resetn, Q => coeff_memory_0_1);
   coeff_memory_reg_4_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n265,
                           CK => clk, RB => resetn, Q => coeff_memory_4_1);
   operand_regs_reg_2_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n254,
                           CK => clk, RB => resetn, Q => operand_regs_161_port)
                           ;
   operand_regs_reg_4_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n258,
                           CK => clk, RB => resetn, Q => operand_regs_97_port);
   operand_regs_reg_6_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n259,
                           CK => clk, RB => resetn, Q => operand_regs_33_port);
   operand_regs_reg_7_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n253,
                           CK => clk, RB => resetn, Q => operand_regs_1_port);
   operand_regs_reg_0_1 : DFERPQ1 port map( D => avs_writedata(1), CEB => n256,
                           CK => clk, RB => resetn, Q => operand_regs_225_port)
                           ;
   coeff_memory_reg_1_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n264,
                           CK => clk, RB => resetn, Q => coeff_memory_1_0);
   coeff_memory_reg_2_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n262,
                           CK => clk, RB => resetn, Q => coeff_memory_2_0);
   coeff_memory_reg_3_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n261,
                           CK => clk, RB => resetn, Q => coeff_memory_3_0);
   coeff_memory_reg_0_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n263,
                           CK => clk, RB => resetn, Q => coeff_memory_0_0);
   coeff_memory_reg_4_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n265,
                           CK => clk, RB => resetn, Q => coeff_memory_4_0);
   operand_regs_reg_2_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n254,
                           CK => clk, RB => resetn, Q => operand_regs_160_port)
                           ;
   operand_regs_reg_4_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n258,
                           CK => clk, RB => resetn, Q => operand_regs_96_port);
   operand_regs_reg_6_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n259,
                           CK => clk, RB => resetn, Q => operand_regs_32_port);
   operand_regs_reg_7_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n253,
                           CK => clk, RB => resetn, Q => operand_regs_0_port);
   operand_regs_reg_0_0 : DFERPQ1 port map( D => avs_writedata(0), CEB => n256,
                           CK => clk, RB => resetn, Q => operand_regs_224_port)
                           ;
   filt_mult_inputs_reg : DFERPQ1 port map( D => avs_writedata(0), CEB => n178,
                           CK => clk, RB => resetn, Q => filt_mult_inputs);
   avs_readdata_reg_30 : DFFSPQ1 port map( D => n203, CK => clk, SB => resetn, 
                           Q => avs_readdata_30_port);
   avs_readdata_reg_28 : DFFSPQ1 port map( D => n205, CK => clk, SB => resetn, 
                           Q => avs_readdata_28_port);
   avs_readdata_reg_26 : DFFSPQ1 port map( D => n207, CK => clk, SB => resetn, 
                           Q => avs_readdata_26_port);
   avs_readdata_reg_24 : DFFSPQ1 port map( D => n209, CK => clk, SB => resetn, 
                           Q => avs_readdata_24_port);
   avs_readdata_reg_22 : DFFSPQ1 port map( D => n211, CK => clk, SB => resetn, 
                           Q => avs_readdata_22_port);
   avs_readdata_reg_20 : DFFSPQ1 port map( D => n213, CK => clk, SB => resetn, 
                           Q => avs_readdata_20_port);
   avs_readdata_reg_18 : DFFSPQ1 port map( D => n215, CK => clk, SB => resetn, 
                           Q => avs_readdata_18_port);
   avs_readdata_reg_16 : DFFSPQ1 port map( D => n217, CK => clk, SB => resetn, 
                           Q => avs_readdata_16_port);
   avs_readdata_reg_14 : DFFSPQ1 port map( D => n219, CK => clk, SB => resetn, 
                           Q => avs_readdata_14_port);
   avs_readdata_reg_12 : DFFSPQ1 port map( D => n221, CK => clk, SB => resetn, 
                           Q => avs_readdata_12_port);
   avs_readdata_reg_10 : DFFSPQ1 port map( D => n223, CK => clk, SB => resetn, 
                           Q => avs_readdata_10_port);
   avs_readdata_reg_8 : DFFSPQ1 port map( D => n225, CK => clk, SB => resetn, Q
                           => avs_readdata_8_port);
   avs_readdata_reg_6 : DFFSPQ1 port map( D => n227, CK => clk, SB => resetn, Q
                           => avs_readdata_6_port);
   avs_readdata_reg_4 : DFFSPQ1 port map( D => n229, CK => clk, SB => resetn, Q
                           => avs_readdata_4_port);
   avs_readdata_reg_2 : DFFSPQ1 port map( D => n231, CK => clk, SB => resetn, Q
                           => avs_readdata_2_port);
   avs_readdata_reg_0 : DFFSPQ1 port map( D => n233, CK => clk, SB => resetn, Q
                           => avs_readdata_0_port);
   avs_readdata_reg_31 : DFFRPQ1 port map( D => n202, CK => clk, RB => resetn, 
                           Q => avs_readdata_31_port);
   avs_readdata_reg_29 : DFFRPQ1 port map( D => n204, CK => clk, RB => resetn, 
                           Q => avs_readdata_29_port);
   avs_readdata_reg_27 : DFFRPQ1 port map( D => n206, CK => clk, RB => resetn, 
                           Q => avs_readdata_27_port);
   avs_readdata_reg_25 : DFFRPQ1 port map( D => n208, CK => clk, RB => resetn, 
                           Q => avs_readdata_25_port);
   avs_readdata_reg_23 : DFFRPQ1 port map( D => n210, CK => clk, RB => resetn, 
                           Q => avs_readdata_23_port);
   avs_readdata_reg_21 : DFFRPQ1 port map( D => n212, CK => clk, RB => resetn, 
                           Q => avs_readdata_21_port);
   avs_readdata_reg_19 : DFFRPQ1 port map( D => n214, CK => clk, RB => resetn, 
                           Q => avs_readdata_19_port);
   avs_readdata_reg_17 : DFFRPQ1 port map( D => n216, CK => clk, RB => resetn, 
                           Q => avs_readdata_17_port);
   avs_readdata_reg_15 : DFFRPQ1 port map( D => n218, CK => clk, RB => resetn, 
                           Q => avs_readdata_15_port);
   avs_readdata_reg_13 : DFFRPQ1 port map( D => n220, CK => clk, RB => resetn, 
                           Q => avs_readdata_13_port);
   avs_readdata_reg_11 : DFFRPQ1 port map( D => n222, CK => clk, RB => resetn, 
                           Q => avs_readdata_11_port);
   avs_readdata_reg_9 : DFFRPQ1 port map( D => n224, CK => clk, RB => resetn, Q
                           => avs_readdata_9_port);
   avs_readdata_reg_7 : DFFRPQ1 port map( D => n226, CK => clk, RB => resetn, Q
                           => avs_readdata_7_port);
   avs_readdata_reg_5 : DFFRPQ1 port map( D => n228, CK => clk, RB => resetn, Q
                           => avs_readdata_5_port);
   avs_readdata_reg_3 : DFFRPQ1 port map( D => n230, CK => clk, RB => resetn, Q
                           => avs_readdata_3_port);
   avs_readdata_reg_1 : DFFRPQ1 port map( D => n232, CK => clk, RB => resetn, Q
                           => avs_readdata_1_port);
   stop_sim_reg : DFFRPQ1 port map( D => n157, CK => clk, RB => resetn, Q => 
                           stop_sim_port);
   siso_req_reg : DFERPQ1 port map( D => n690, CEB => n161, CK => clk, RB => 
                           resetn, Q => siso_req);
   siso_data_out_reg_0 : DFERPQ1 port map( D => N2888, CEB => n695, CK => clk, 
                           RB => resetn, Q => siso_data_out(0));
   siso_data_out_reg_15 : DFERPQ1 port map( D => N2903, CEB => n695, CK => clk,
                           RB => resetn, Q => siso_data_out(15));
   siso_data_out_reg_14 : DFERPQ1 port map( D => N2902, CEB => n695, CK => clk,
                           RB => resetn, Q => siso_data_out(14));
   siso_data_out_reg_13 : DFERPQ1 port map( D => N2901, CEB => n695, CK => clk,
                           RB => resetn, Q => siso_data_out(13));
   siso_data_out_reg_12 : DFERPQ1 port map( D => N2900, CEB => n695, CK => clk,
                           RB => resetn, Q => siso_data_out(12));
   siso_data_out_reg_11 : DFERPQ1 port map( D => N2899, CEB => n695, CK => clk,
                           RB => resetn, Q => siso_data_out(11));
   siso_data_out_reg_10 : DFERPQ1 port map( D => N2898, CEB => n695, CK => clk,
                           RB => resetn, Q => siso_data_out(10));
   siso_data_out_reg_9 : DFERPQ1 port map( D => N2897, CEB => n695, CK => clk, 
                           RB => resetn, Q => siso_data_out(9));
   siso_data_out_reg_8 : DFERPQ1 port map( D => N2896, CEB => n695, CK => clk, 
                           RB => resetn, Q => siso_data_out(8));
   siso_data_out_reg_7 : DFERPQ1 port map( D => N2895, CEB => n695, CK => clk, 
                           RB => resetn, Q => siso_data_out(7));
   siso_data_out_reg_6 : DFERPQ1 port map( D => N2894, CEB => n695, CK => clk, 
                           RB => resetn, Q => siso_data_out(6));
   siso_data_out_reg_5 : DFERPQ1 port map( D => N2893, CEB => n695, CK => clk, 
                           RB => resetn, Q => siso_data_out(5));
   siso_data_out_reg_4 : DFERPQ1 port map( D => N2892, CEB => n695, CK => clk, 
                           RB => resetn, Q => siso_data_out(4));
   siso_data_out_reg_3 : DFERPQ1 port map( D => N2891, CEB => n695, CK => clk, 
                           RB => resetn, Q => siso_data_out(3));
   siso_data_out_reg_2 : DFERPQ1 port map( D => N2890, CEB => n695, CK => clk, 
                           RB => resetn, Q => siso_data_out(2));
   siso_data_out_reg_1 : DFERPQ1 port map( D => N2889, CEB => n695, CK => clk, 
                           RB => resetn, Q => siso_data_out(1));
   siso_ready_reg : DFFRPQ1 port map( D => out_busy, CK => clk, RB => resetn, Q
                           => siso_ready);
   U642 : AND2D1 port map( A1 => n289, A2 => avs_addr(0), Z => n242);
   U643 : AND2D1 port map( A1 => n536, A2 => N62, Z => n243);
   U644 : AND2D1 port map( A1 => n538, A2 => N62, Z => n244);
   U645 : NAN3D1 port map( A1 => n106, A2 => avs_addr(0), A3 => n110, Z => n245
                           );
   U646 : NAN2D1 port map( A1 => n110, A2 => n99, Z => n246);
   U647 : NAN2D1 port map( A1 => n110, A2 => n97, Z => n247);
   U648 : NAN2D1 port map( A1 => n110, A2 => n93, Z => n248);
   U649 : NAN2D1 port map( A1 => n110, A2 => n109, Z => n249);
   U650 : NAN2D1 port map( A1 => n110, A2 => n108, Z => n250);
   U651 : NAN2D1 port map( A1 => n110, A2 => n69, Z => n251);
   U652 : NAN2D1 port map( A1 => n110, A2 => n68, Z => n252);
   U653 : NAN3D1 port map( A1 => n106, A2 => avs_addr(0), A3 => n107, Z => n253
                           );
   U654 : NAN2D1 port map( A1 => n107, A2 => n69, Z => n254);
   U655 : NAN2D1 port map( A1 => n107, A2 => n68, Z => n255);
   U656 : NAN2D1 port map( A1 => n107, A2 => n97, Z => n256);
   U657 : NAN2D1 port map( A1 => n107, A2 => n93, Z => n257);
   U658 : NAN2D1 port map( A1 => n107, A2 => n99, Z => n258);
   U659 : NAN2D1 port map( A1 => n108, A2 => n107, Z => n259);
   U660 : NAN2D1 port map( A1 => n109, A2 => n107, Z => n260);
   U661 : NAN2D1 port map( A1 => n103, A2 => n68, Z => n261);
   U662 : NAN2D1 port map( A1 => n103, A2 => n69, Z => n262);
   U663 : NAN2D1 port map( A1 => n103, A2 => n97, Z => n263);
   U664 : NAN2D1 port map( A1 => n103, A2 => n93, Z => n264);
   U665 : NAN2D1 port map( A1 => n103, A2 => n99, Z => n265);
   U666 : AND2D1 port map( A1 => n288, A2 => avs_addr(0), Z => n266);
   U667 : AND3D1 port map( A1 => N66, A2 => n270, A3 => read_comp_res, Z => 
                           n267);
   U668 : AND2D1 port map( A1 => n535, A2 => N62, Z => n268);
   U669 : AND2D1 port map( A1 => n537, A2 => N62, Z => n269);
   U670 : BUFBD2 port map( A => filt_mult_inputs, Z => n673);
   U671 : INVD1 port map( A => n528, Z => n529);
   U672 : INVD1 port map( A => n533, Z => n534);
   U673 : INVD1 port map( A => n530, Z => n532);
   U674 : INVD1 port map( A => n530, Z => n531);
   U675 : INVD1 port map( A => n526, Z => n527);
   U676 : INVD1 port map( A => n523, Z => n524);
   U677 : INVD1 port map( A => n523, Z => n525);
   U678 : INVD1 port map( A => n74, Z => n677);
   U679 : INVD1 port map( A => n96, Z => n678);
   U680 : NAN2D1 port map( A1 => n118, A2 => n691, Z => n176);
   U681 : NAN2D1 port map( A1 => n689, A2 => n118, Z => n174);
   U682 : NOR2M1D1 port map( A1 => n104, A2 => n686, Z => n103);
   U683 : INVD1 port map( A => n270, Z => n676);
   U684 : INVD1 port map( A => n516, Z => n528);
   U685 : INVD1 port map( A => n518, Z => n533);
   U686 : INVD1 port map( A => n517, Z => n530);
   U687 : INVD1 port map( A => n675, Z => n674);
   U688 : INVD1 port map( A => n513, Z => n523);
   U689 : INVD1 port map( A => n514, Z => n526);
   U690 : NAN2D1 port map( A1 => n93, A2 => n679, Z => n74);
   U691 : OAI211D1 port map( A1 => n6300, A2 => n6400, B => n270, C => n65, Z 
                           => n14);
   U692 : NOR2D1 port map( A1 => n68, A2 => n69, Z => n6300);
   U693 : NOR3D1 port map( A1 => n677, A2 => N66, A3 => n678, Z => n65);
   U694 : AND2D1 port map( A1 => n111, A2 => n681, Z => n99);
   U695 : INVD1 port map( A => n6400, Z => n679);
   U696 : NAN2D1 port map( A1 => n97, A2 => n679, Z => n96);
   U697 : AND2D1 port map( A1 => n106, A2 => n681, Z => n108);
   U698 : INVD1 port map( A => n673, Z => n276);
   U699 : INVD1 port map( A => n673, Z => n278);
   U700 : INVD1 port map( A => n673, Z => n279);
   U701 : INVD1 port map( A => n673, Z => n275);
   U702 : INVD1 port map( A => n673, Z => n281);
   U703 : INVD1 port map( A => n673, Z => n272);
   U704 : INVD1 port map( A => n673, Z => n285);
   U705 : INVD1 port map( A => n673, Z => n284);
   U706 : INVD1 port map( A => n673, Z => n280);
   U707 : INVD1 port map( A => n673, Z => n286);
   U708 : INVD1 port map( A => n673, Z => n271);
   U709 : INVD1 port map( A => n673, Z => n273);
   U710 : INVD1 port map( A => n673, Z => n274);
   U711 : INVD1 port map( A => n673, Z => n282);
   U712 : INVD1 port map( A => n673, Z => n277);
   U713 : INVD1 port map( A => n673, Z => n283);
   U714 : INVD1 port map( A => n673, Z => n287);
   U715 : NOR3D1 port map( A1 => n697, A2 => n694, A3 => n671, Z => n78);
   U716 : INVD1 port map( A => n81, Z => n684);
   U717 : INVD1 port map( A => n672, Z => n696);
   U718 : NOR2D1 port map( A1 => n693, A2 => n687, Z => n118);
   U719 : INVD1 port map( A => n88, Z => n691);
   U720 : NOR2D1 port map( A1 => n683, A2 => n91, Z => n89);
   U721 : INVD1 port map( A => n84, Z => n683);
   U722 : INVD1 port map( A => n155, Z => n688);
   U723 : NAN2D1 port map( A1 => n119, A2 => n115, Z => n171);
   U724 : NAN2D1 port map( A1 => n119, A2 => n101, Z => n162);
   U725 : NAN2D1 port map( A1 => n119, A2 => n118, Z => n170);
   U726 : NAN2D1 port map( A1 => n120, A2 => n119, Z => n163);
   U727 : NAN2D1 port map( A1 => n87, A2 => n84, Z => n86);
   U728 : NAN2D1 port map( A1 => n689, A2 => n115, Z => n175);
   U729 : NAN2D1 port map( A1 => n120, A2 => n689, Z => n167);
   U730 : NAN2D1 port map( A1 => n689, A2 => n101, Z => n166);
   U731 : INVD1 port map( A => n85, Z => n689);
   U732 : NAN2D1 port map( A1 => n87, A2 => n101, Z => n164);
   U733 : NAN2D1 port map( A1 => n115, A2 => n87, Z => n173);
   U734 : NAN2D1 port map( A1 => n120, A2 => n87, Z => n165);
   U735 : NAN2D1 port map( A1 => n118, A2 => n87, Z => n172);
   U736 : NAN2D1 port map( A1 => n691, A2 => n101, Z => n168);
   U737 : NAN2D1 port map( A1 => n115, A2 => n691, Z => n177);
   U738 : NAN2D1 port map( A1 => n120, A2 => n691, Z => n169);
   U739 : NOR3M1D1 port map( A1 => n104, A2 => coeff_load, A3 => operand_load, 
                           Z => n110);
   U740 : AND2D1 port map( A1 => N66, A2 => avs_write, Z => n104);
   U741 : AND3D1 port map( A1 => n686, A2 => n104, A3 => operand_load, Z => 
                           n107);
   U742 : NAN4D1 port map( A1 => n5900, A2 => n14, A3 => n6000, A4 => n6100, Z 
                           => n233);
   U743 : NAN2M1D1 port map( A1 => n70, A2 => n270, Z => n5900);
   U744 : NAN2D1 port map( A1 => N2009, A2 => n267, Z => n6000);
   U745 : INVD1 port map( A => n12, Z => n675);
   U746 : NOR3M1D1 port map( A1 => N66, A2 => n676, A3 => read_comp_res, Z => 
                           n12);
   U747 : INVD1 port map( A => avs_write, Z => n682);
   U748 : AND2D1 port map( A1 => avs_read, A2 => n682, Z => n270);
   U749 : NAN3D1 port map( A1 => n56, A2 => n14, A3 => n57, Z => n231);
   U750 : NAN2D1 port map( A1 => N2007, A2 => n267, Z => n56);
   U751 : NAN3D1 port map( A1 => n427, A2 => n426, A3 => n428, Z => N2007);
   U752 : NAN3D1 port map( A1 => n53, A2 => n14, A3 => n54, Z => n229);
   U753 : NAN2D1 port map( A1 => N2005, A2 => n267, Z => n53);
   U754 : NAN3D1 port map( A1 => n433, A2 => n432, A3 => n434, Z => N2005);
   U755 : NAN3D1 port map( A1 => n50, A2 => n14, A3 => n51, Z => n227);
   U756 : NAN2D1 port map( A1 => N2003, A2 => n267, Z => n50);
   U757 : NAN3D1 port map( A1 => n439, A2 => n438, A3 => n440, Z => N2003);
   U758 : NAN3D1 port map( A1 => n47, A2 => n14, A3 => n48, Z => n225);
   U759 : NAN2D1 port map( A1 => N2001, A2 => n267, Z => n47);
   U760 : NAN3D1 port map( A1 => n445, A2 => n444, A3 => n446, Z => N2001);
   U761 : NAN3D1 port map( A1 => n44, A2 => n14, A3 => n45, Z => n223);
   U762 : NAN2D1 port map( A1 => N1999, A2 => n267, Z => n44);
   U763 : NAN3D1 port map( A1 => n451, A2 => n450, A3 => n452, Z => N1999);
   U764 : NAN3D1 port map( A1 => n41, A2 => n14, A3 => n42, Z => n221);
   U765 : NAN2D1 port map( A1 => N1997, A2 => n267, Z => n41);
   U766 : NAN3D1 port map( A1 => n457, A2 => n456, A3 => n458, Z => N1997);
   U767 : NAN3D1 port map( A1 => n38, A2 => n14, A3 => n39, Z => n219);
   U768 : NAN2D1 port map( A1 => N1995, A2 => n267, Z => n38);
   U769 : NAN3D1 port map( A1 => n463, A2 => n462, A3 => n464, Z => N1995);
   U770 : NAN3D1 port map( A1 => n35, A2 => n14, A3 => n36, Z => n217);
   U771 : NAN2D1 port map( A1 => N1993, A2 => n267, Z => n35);
   U772 : NAN3D1 port map( A1 => n469, A2 => n468, A3 => n470, Z => N1993);
   U773 : NAN3D1 port map( A1 => n13, A2 => n14, A3 => n15, Z => n203);
   U774 : NAN2D1 port map( A1 => N1979, A2 => n267, Z => n13);
   U775 : NAN3D1 port map( A1 => n511, A2 => n510, A3 => n512, Z => N1979);
   U776 : INVD1 port map( A => avs_addr(2), Z => n522);
   U777 : NAN3D1 port map( A1 => n32, A2 => n14, A3 => n33, Z => n215);
   U778 : NAN2D1 port map( A1 => N1991, A2 => n267, Z => n32);
   U779 : NAN3D1 port map( A1 => n475, A2 => n474, A3 => n476, Z => N1991);
   U780 : NAN3D1 port map( A1 => n29, A2 => n14, A3 => n30, Z => n213);
   U781 : NAN2D1 port map( A1 => N1989, A2 => n267, Z => n29);
   U782 : NAN3D1 port map( A1 => n481, A2 => n480, A3 => n482, Z => N1989);
   U783 : NAN3D1 port map( A1 => n26, A2 => n14, A3 => n27, Z => n211);
   U784 : NAN2D1 port map( A1 => N1987, A2 => n267, Z => n26);
   U785 : NAN3D1 port map( A1 => n487, A2 => n486, A3 => n488, Z => N1987);
   U786 : NAN3D1 port map( A1 => n23, A2 => n14, A3 => n24, Z => n209);
   U787 : NAN2D1 port map( A1 => N1985, A2 => n267, Z => n23);
   U788 : NAN3D1 port map( A1 => n493, A2 => n492, A3 => n494, Z => N1985);
   U789 : NAN3D1 port map( A1 => n20, A2 => n14, A3 => n21, Z => n207);
   U790 : NAN2D1 port map( A1 => N1983, A2 => n267, Z => n20);
   U791 : NAN3D1 port map( A1 => n499, A2 => n498, A3 => n500, Z => N1983);
   U792 : NAN3D1 port map( A1 => n17, A2 => n14, A3 => n18, Z => n205);
   U793 : NAN2D1 port map( A1 => N1981, A2 => n267, Z => n17);
   U794 : NAN3D1 port map( A1 => n505, A2 => n504, A3 => n506, Z => N1981);
   U795 : OAI21M20D1 port map( A1 => avs_readdata_1_port, A2 => n676, B => n58,
                           Z => n232);
   U796 : NAN3D1 port map( A1 => n424, A2 => n423, A3 => n425, Z => N2008);
   U797 : OAI21M20D1 port map( A1 => avs_readdata_3_port, A2 => n676, B => n55,
                           Z => n230);
   U798 : NAN3D1 port map( A1 => n430, A2 => n429, A3 => n431, Z => N2006);
   U799 : OAI21M20D1 port map( A1 => avs_readdata_5_port, A2 => n676, B => n52,
                           Z => n228);
   U800 : NAN3D1 port map( A1 => n436, A2 => n435, A3 => n437, Z => N2004);
   U801 : OAI21M20D1 port map( A1 => avs_readdata_7_port, A2 => n676, B => n49,
                           Z => n226);
   U802 : NAN3D1 port map( A1 => n442, A2 => n441, A3 => n443, Z => N2002);
   U803 : OAI21M20D1 port map( A1 => avs_readdata_15_port, A2 => n676, B => n37
                           , Z => n218);
   U804 : NAN3D1 port map( A1 => n466, A2 => n465, A3 => n467, Z => N1994);
   U805 : OAI21M20D1 port map( A1 => avs_readdata_17_port, A2 => n676, B => n34
                           , Z => n216);
   U806 : NAN3D1 port map( A1 => n472, A2 => n471, A3 => n473, Z => N1992);
   U807 : OAI21M20D1 port map( A1 => avs_readdata_19_port, A2 => n676, B => n31
                           , Z => n214);
   U808 : NAN3D1 port map( A1 => n478, A2 => n477, A3 => n479, Z => N1990);
   U809 : OAI21M20D1 port map( A1 => avs_readdata_21_port, A2 => n676, B => n28
                           , Z => n212);
   U810 : NAN3D1 port map( A1 => n484, A2 => n483, A3 => n485, Z => N1988);
   U811 : OAI21M20D1 port map( A1 => avs_readdata_23_port, A2 => n676, B => n25
                           , Z => n210);
   U812 : NAN3D1 port map( A1 => n490, A2 => n489, A3 => n491, Z => N1986);
   U813 : OAI21M20D1 port map( A1 => avs_readdata_25_port, A2 => n676, B => n22
                           , Z => n208);
   U814 : NAN3D1 port map( A1 => n496, A2 => n495, A3 => n497, Z => N1984);
   U815 : OAI21M20D1 port map( A1 => avs_readdata_27_port, A2 => n676, B => n19
                           , Z => n206);
   U816 : NAN3D1 port map( A1 => n502, A2 => n501, A3 => n503, Z => N1982);
   U817 : OAI21M20D1 port map( A1 => avs_readdata_29_port, A2 => n676, B => n16
                           , Z => n204);
   U818 : NAN3D1 port map( A1 => n508, A2 => n507, A3 => n509, Z => N1980);
   U819 : OAI21M20D1 port map( A1 => avs_readdata_31_port, A2 => n676, B => n10
                           , Z => n202);
   U820 : OAI21M20D1 port map( A1 => avs_readdata_9_port, A2 => n676, B => n46,
                           Z => n224);
   U821 : NAN3D1 port map( A1 => n448, A2 => n447, A3 => n449, Z => N2000);
   U822 : OAI21M20D1 port map( A1 => avs_readdata_11_port, A2 => n676, B => n43
                           , Z => n222);
   U823 : NAN3D1 port map( A1 => n454, A2 => n453, A3 => n455, Z => N1998);
   U824 : OAI21M20D1 port map( A1 => avs_readdata_13_port, A2 => n676, B => n40
                           , Z => n220);
   U825 : NAN3D1 port map( A1 => n460, A2 => n459, A3 => n461, Z => N1996);
   U826 : NAN3D1 port map( A1 => n520, A2 => n519, A3 => n521, Z => N1978);
   U827 : NAN2D1 port map( A1 => comp_res_31_port, A2 => n529, Z => n520);
   U828 : AOI22M10D1 port map( B1 => in_buf_63_port, B2 => n515, A1 => n528, A2
                           => in_buf_127_port, Z => n417);
   U829 : NAN3D1 port map( A1 => n421, A2 => n420, A3 => n422, Z => N2009);
   U830 : NAN2D1 port map( A1 => comp_res_0_port, A2 => n529, Z => n421);
   U831 : NAN2D1 port map( A1 => comp_res_25_port, A2 => n529, Z => n496);
   U832 : NAN2D1 port map( A1 => comp_res_27_port, A2 => n529, Z => n502);
   U833 : NAN2D1 port map( A1 => comp_res_29_port, A2 => n529, Z => n508);
   U834 : NAN2D1 port map( A1 => comp_res_1_port, A2 => n529, Z => n424);
   U835 : NAN2D1 port map( A1 => comp_res_3_port, A2 => n529, Z => n430);
   U836 : NAN2D1 port map( A1 => comp_res_5_port, A2 => n529, Z => n436);
   U837 : NAN2D1 port map( A1 => comp_res_7_port, A2 => n529, Z => n442);
   U838 : NAN2D1 port map( A1 => comp_res_9_port, A2 => n529, Z => n448);
   U839 : NAN2D1 port map( A1 => comp_res_11_port, A2 => n529, Z => n454);
   U840 : NAN2D1 port map( A1 => comp_res_13_port, A2 => n529, Z => n460);
   U841 : NAN2D1 port map( A1 => comp_res_15_port, A2 => n529, Z => n466);
   U842 : NAN2D1 port map( A1 => comp_res_17_port, A2 => n516, Z => n472);
   U843 : NAN2D1 port map( A1 => comp_res_19_port, A2 => n529, Z => n478);
   U844 : NAN2D1 port map( A1 => comp_res_21_port, A2 => n516, Z => n484);
   U845 : NAN2D1 port map( A1 => comp_res_23_port, A2 => n516, Z => n490);
   U846 : NAN2D1 port map( A1 => comp_res_24_port, A2 => n529, Z => n493);
   U847 : NAN2D1 port map( A1 => comp_res_26_port, A2 => n529, Z => n499);
   U848 : NAN2D1 port map( A1 => comp_res_28_port, A2 => n529, Z => n505);
   U849 : NAN2D1 port map( A1 => comp_res_30_port, A2 => n529, Z => n511);
   U850 : NAN2D1 port map( A1 => comp_res_2_port, A2 => n516, Z => n427);
   U851 : NAN2D1 port map( A1 => comp_res_4_port, A2 => n516, Z => n433);
   U852 : NAN2D1 port map( A1 => comp_res_6_port, A2 => n516, Z => n439);
   U853 : NAN2D1 port map( A1 => comp_res_8_port, A2 => n516, Z => n445);
   U854 : NAN2D1 port map( A1 => comp_res_10_port, A2 => n516, Z => n451);
   U855 : NAN2D1 port map( A1 => comp_res_12_port, A2 => n516, Z => n457);
   U856 : NAN2D1 port map( A1 => comp_res_14_port, A2 => n516, Z => n463);
   U857 : NAN2D1 port map( A1 => comp_res_16_port, A2 => n516, Z => n469);
   U858 : NAN2D1 port map( A1 => comp_res_18_port, A2 => n516, Z => n475);
   U859 : NAN2D1 port map( A1 => comp_res_20_port, A2 => n516, Z => n481);
   U860 : NAN2D1 port map( A1 => comp_res_22_port, A2 => n516, Z => n487);
   U861 : NOR3D1 port map( A1 => avs_addr(1), A2 => avs_addr(2), A3 => n681, Z 
                           => n93);
   U862 : INVD1 port map( A => avs_addr(0), Z => n681);
   U863 : NOR3D1 port map( A1 => n681, A2 => avs_addr(2), A3 => n680, Z => n68)
                           ;
   U864 : INVD1 port map( A => avs_addr(1), Z => n680);
   U865 : NOR3D1 port map( A1 => avs_addr(0), A2 => avs_addr(2), A3 => n680, Z 
                           => n69);
   U866 : AND2D1 port map( A1 => avs_addr(2), A2 => n680, Z => n111);
   U867 : AND2D1 port map( A1 => n111, A2 => avs_addr(0), Z => n109);
   U868 : NAN2D1 port map( A1 => n114, A2 => avs_addr(3), Z => n6400);
   U869 : NOR2D1 port map( A1 => avs_addr(5), A2 => avs_addr(4), Z => n114);
   U870 : AND2D1 port map( A1 => avs_addr(2), A2 => avs_addr(1), Z => n106);
   U871 : NOR3D1 port map( A1 => avs_addr(1), A2 => avs_addr(2), A3 => 
                           avs_addr(0), Z => n97);
   U872 : NOR2D1 port map( A1 => n92, A2 => n682, Z => n240);
   U873 : NOR2D1 port map( A1 => n95, A2 => n682, Z => n241);
   U874 : NAN3D1 port map( A1 => avs_write, A2 => n679, A3 => n109, Z => n179);
   U875 : AO31D1 port map( A1 => avs_write, A2 => n679, A3 => n99, B => 
                           stop_sim_port, Z => n157);
   U876 : NAN3D1 port map( A1 => avs_write, A2 => n679, A3 => n108, Z => n178);
   U877 : AO22D1 port map( A1 => operand_regs_32_port, A2 => n278, B1 => 
                           coeff_memory_3_0, B2 => n673, Z => N3009);
   U878 : AO22D1 port map( A1 => operand_regs_96_port, A2 => n279, B1 => 
                           coeff_memory_2_0, B2 => n673, Z => N2977);
   U879 : AO22D1 port map( A1 => operand_regs_160_port, A2 => n276, B1 => 
                           coeff_memory_1_0, B2 => n673, Z => N2945);
   U880 : AO22D1 port map( A1 => coeff_memory_4_0, A2 => n673, B1 => n275, B2 
                           => operand_regs_0_port, Z => N3041);
   U881 : AO22D1 port map( A1 => coeff_memory_0_0, A2 => n673, B1 => n275, B2 
                           => operand_regs_224_port, Z => N2913);
   U882 : AO22D1 port map( A1 => operand_regs_33_port, A2 => n276, B1 => 
                           coeff_memory_3_1, B2 => n673, Z => N3010);
   U883 : AO22D1 port map( A1 => operand_regs_97_port, A2 => n278, B1 => 
                           coeff_memory_2_1, B2 => n673, Z => N2978);
   U884 : AO22D1 port map( A1 => operand_regs_161_port, A2 => n281, B1 => 
                           coeff_memory_1_1, B2 => n673, Z => N2946);
   U885 : AO22D1 port map( A1 => coeff_memory_4_1, A2 => n673, B1 => n275, B2 
                           => operand_regs_1_port, Z => N3042);
   U886 : AO22D1 port map( A1 => coeff_memory_0_1, A2 => n673, B1 => n272, B2 
                           => operand_regs_225_port, Z => N2914);
   U887 : AO22D1 port map( A1 => n673, A2 => operand_regs_194_port, B1 => n272,
                           B2 => operand_regs_2_port, Z => N3203);
   U888 : AO22D1 port map( A1 => n673, A2 => operand_regs_193_port, B1 => n272,
                           B2 => operand_regs_1_port, Z => N3202);
   U889 : OAI21M20D1 port map( A1 => operand_regs_66_port, A2 => n285, B => 
                           n151, Z => N3139);
   U890 : OAI21M20D1 port map( A1 => operand_regs_130_port, A2 => n285, B => 
                           n151, Z => N3107);
   U891 : OAI21M20D1 port map( A1 => operand_regs_65_port, A2 => n285, B => 
                           n152, Z => N3138);
   U892 : OAI21M20D1 port map( A1 => operand_regs_129_port, A2 => n284, B => 
                           n152, Z => N3106);
   U893 : AO22D1 port map( A1 => operand_regs_34_port, A2 => n278, B1 => 
                           coeff_memory_3_2, B2 => n673, Z => N3011);
   U894 : AO22D1 port map( A1 => operand_regs_98_port, A2 => n280, B1 => 
                           coeff_memory_2_2, B2 => n673, Z => N2979);
   U895 : AO22D1 port map( A1 => operand_regs_162_port, A2 => n281, B1 => 
                           coeff_memory_1_2, B2 => n673, Z => N2947);
   U896 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_194_port, B => 
                           n151, Z => N3075);
   U897 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_193_port, B => 
                           n152, Z => N3074);
   U898 : AO22D1 port map( A1 => n673, A2 => operand_regs_192_port, B1 => n271,
                           B2 => operand_regs_0_port, Z => N3201);
   U899 : AO22D1 port map( A1 => coeff_memory_4_2, A2 => n673, B1 => n275, B2 
                           => operand_regs_2_port, Z => N3043);
   U900 : AO22D1 port map( A1 => coeff_memory_0_2, A2 => n673, B1 => n271, B2 
                           => operand_regs_226_port, Z => N2915);
   U901 : OAI21M20D1 port map( A1 => operand_regs_64_port, A2 => n285, B => 
                           n153, Z => N3137);
   U902 : OAI21M20D1 port map( A1 => operand_regs_128_port, A2 => n284, B => 
                           n153, Z => N3105);
   U903 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_192_port, B => 
                           n153, Z => N3073);
   U904 : AO22D1 port map( A1 => operand_regs_35_port, A2 => n276, B1 => 
                           coeff_memory_3_3, B2 => n673, Z => N3012);
   U905 : AO22D1 port map( A1 => operand_regs_99_port, A2 => n280, B1 => 
                           coeff_memory_2_3, B2 => n673, Z => N2980);
   U906 : AO22D1 port map( A1 => operand_regs_163_port, A2 => n281, B1 => 
                           coeff_memory_1_3, B2 => n673, Z => N2948);
   U907 : AO22D1 port map( A1 => coeff_memory_4_3, A2 => n673, B1 => n275, B2 
                           => operand_regs_3_port, Z => N3044);
   U908 : AO22D1 port map( A1 => coeff_memory_0_3, A2 => n673, B1 => n272, B2 
                           => operand_regs_227_port, Z => N2916);
   U909 : AO22D1 port map( A1 => operand_regs_36_port, A2 => n278, B1 => 
                           coeff_memory_3_4, B2 => n673, Z => N3013);
   U910 : AO22D1 port map( A1 => operand_regs_100_port, A2 => n280, B1 => 
                           coeff_memory_2_4, B2 => n673, Z => N2981);
   U911 : AO22D1 port map( A1 => operand_regs_164_port, A2 => n281, B1 => 
                           coeff_memory_1_4, B2 => n673, Z => N2949);
   U912 : AO22D1 port map( A1 => n673, A2 => operand_regs_195_port, B1 => n273,
                           B2 => operand_regs_3_port, Z => N3204);
   U913 : AO22D1 port map( A1 => coeff_memory_4_4, A2 => n673, B1 => n275, B2 
                           => operand_regs_4_port, Z => N3045);
   U914 : AO22D1 port map( A1 => coeff_memory_0_4, A2 => n673, B1 => n272, B2 
                           => operand_regs_228_port, Z => N2917);
   U915 : AO22D1 port map( A1 => n673, A2 => operand_regs_196_port, B1 => n272,
                           B2 => operand_regs_4_port, Z => N3205);
   U916 : NAN2D1 port map( A1 => operand_regs_226_port, A2 => n673, Z => n151);
   U917 : NAN2D1 port map( A1 => operand_regs_225_port, A2 => n673, Z => n152);
   U918 : OAI21M20D1 port map( A1 => operand_regs_67_port, A2 => n285, B => 
                           n150, Z => N3140);
   U919 : OAI21M20D1 port map( A1 => operand_regs_131_port, A2 => n285, B => 
                           n150, Z => N3108);
   U920 : OAI21M20D1 port map( A1 => operand_regs_68_port, A2 => n285, B => 
                           n149, Z => N3141);
   U921 : OAI21M20D1 port map( A1 => operand_regs_132_port, A2 => n285, B => 
                           n149, Z => N3109);
   U922 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_195_port, B => 
                           n150, Z => N3076);
   U923 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_196_port, B => 
                           n149, Z => N3077);
   U924 : AO22D1 port map( A1 => operand_regs_37_port, A2 => n276, B1 => 
                           coeff_memory_3_5, B2 => n673, Z => N3014);
   U925 : AO22D1 port map( A1 => operand_regs_101_port, A2 => n280, B1 => 
                           coeff_memory_2_5, B2 => n673, Z => N2982);
   U926 : AO22D1 port map( A1 => operand_regs_165_port, A2 => n281, B1 => 
                           coeff_memory_1_5, B2 => n673, Z => N2950);
   U927 : NAN2D1 port map( A1 => operand_regs_224_port, A2 => n673, Z => n153);
   U928 : AO22D1 port map( A1 => coeff_memory_4_5, A2 => n673, B1 => n274, B2 
                           => operand_regs_5_port, Z => N3046);
   U929 : AO22D1 port map( A1 => coeff_memory_0_5, A2 => n673, B1 => n272, B2 
                           => operand_regs_229_port, Z => N2918);
   U930 : AO22D1 port map( A1 => operand_regs_38_port, A2 => n278, B1 => 
                           coeff_memory_3_6, B2 => n673, Z => N3015);
   U931 : AO22D1 port map( A1 => operand_regs_102_port, A2 => n280, B1 => 
                           coeff_memory_2_6, B2 => n673, Z => N2983);
   U932 : AO22D1 port map( A1 => operand_regs_166_port, A2 => n281, B1 => 
                           coeff_memory_1_6, B2 => n673, Z => N2951);
   U933 : AO22D1 port map( A1 => coeff_memory_4_6, A2 => n673, B1 => n274, B2 
                           => operand_regs_6_port, Z => N3047);
   U934 : AO22D1 port map( A1 => coeff_memory_0_6, A2 => n673, B1 => n272, B2 
                           => operand_regs_230_port, Z => N2919);
   U935 : NAN2D1 port map( A1 => operand_regs_227_port, A2 => n673, Z => n150);
   U936 : NAN2D1 port map( A1 => operand_regs_228_port, A2 => n673, Z => n149);
   U937 : AO22D1 port map( A1 => n673, A2 => operand_regs_197_port, B1 => n271,
                           B2 => operand_regs_5_port, Z => N3206);
   U938 : AO22D1 port map( A1 => operand_regs_39_port, A2 => n277, B1 => 
                           coeff_memory_3_7, B2 => n673, Z => N3016);
   U939 : AO22D1 port map( A1 => operand_regs_103_port, A2 => n280, B1 => 
                           coeff_memory_2_7, B2 => n673, Z => N2984);
   U940 : AO22D1 port map( A1 => operand_regs_167_port, A2 => n282, B1 => 
                           coeff_memory_1_7, B2 => n673, Z => N2952);
   U941 : OAI21M20D1 port map( A1 => operand_regs_69_port, A2 => n285, B => 
                           n148, Z => N3142);
   U942 : OAI21M20D1 port map( A1 => operand_regs_133_port, A2 => n284, B => 
                           n148, Z => N3110);
   U943 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_197_port, B => 
                           n148, Z => N3078);
   U944 : AO22D1 port map( A1 => coeff_memory_4_7, A2 => n673, B1 => n274, B2 
                           => operand_regs_7_port, Z => N3048);
   U945 : AO22D1 port map( A1 => coeff_memory_0_7, A2 => n673, B1 => n272, B2 
                           => operand_regs_231_port, Z => N2920);
   U946 : AO22D1 port map( A1 => n673, A2 => operand_regs_198_port, B1 => n272,
                           B2 => operand_regs_6_port, Z => N3207);
   U947 : OAI21M20D1 port map( A1 => operand_regs_134_port, A2 => n283, B => 
                           n147, Z => N3111);
   U948 : OAI21M20D1 port map( A1 => operand_regs_70_port, A2 => n285, B => 
                           n147, Z => N3143);
   U949 : NAN2D1 port map( A1 => operand_regs_229_port, A2 => n673, Z => n148);
   U950 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_198_port, B => 
                           n147, Z => N3079);
   U951 : AO22D1 port map( A1 => n673, A2 => operand_regs_200_port, B1 => n271,
                           B2 => operand_regs_8_port, Z => N3209);
   U952 : AO22D1 port map( A1 => n673, A2 => operand_regs_199_port, B1 => n273,
                           B2 => operand_regs_7_port, Z => N3208);
   U953 : AO22D1 port map( A1 => operand_regs_40_port, A2 => n278, B1 => 
                           coeff_memory_3_8, B2 => n673, Z => N3017);
   U954 : AO22D1 port map( A1 => operand_regs_104_port, A2 => n280, B1 => 
                           coeff_memory_2_8, B2 => n673, Z => N2985);
   U955 : AO22D1 port map( A1 => operand_regs_168_port, A2 => n282, B1 => 
                           coeff_memory_1_8, B2 => n673, Z => N2953);
   U956 : AO22D1 port map( A1 => coeff_memory_4_8, A2 => n673, B1 => n274, B2 
                           => operand_regs_8_port, Z => N3049);
   U957 : AO22D1 port map( A1 => coeff_memory_0_8, A2 => n673, B1 => n273, B2 
                           => operand_regs_232_port, Z => N2921);
   U958 : OAI21M20D1 port map( A1 => operand_regs_136_port, A2 => n283, B => 
                           n145, Z => N3113);
   U959 : OAI21M20D1 port map( A1 => operand_regs_72_port, A2 => n285, B => 
                           n145, Z => N3145);
   U960 : OAI21M20D1 port map( A1 => operand_regs_71_port, A2 => n285, B => 
                           n146, Z => N3144);
   U961 : OAI21M20D1 port map( A1 => operand_regs_135_port, A2 => n284, B => 
                           n146, Z => N3112);
   U962 : OAI21M20D1 port map( A1 => n283, A2 => operand_regs_199_port, B => 
                           n146, Z => N3080);
   U963 : OAI21M20D1 port map( A1 => n287, A2 => operand_regs_200_port, B => 
                           n145, Z => N3081);
   U964 : NAN2D1 port map( A1 => operand_regs_230_port, A2 => n673, Z => n147);
   U965 : AO22D1 port map( A1 => operand_regs_41_port, A2 => n276, B1 => 
                           coeff_memory_3_9, B2 => n673, Z => N3018);
   U966 : AO22D1 port map( A1 => operand_regs_105_port, A2 => n280, B1 => 
                           coeff_memory_2_9, B2 => n673, Z => N2986);
   U967 : AO22D1 port map( A1 => operand_regs_169_port, A2 => n282, B1 => 
                           coeff_memory_1_9, B2 => n673, Z => N2954);
   U968 : AO22D1 port map( A1 => coeff_memory_4_9, A2 => n673, B1 => n274, B2 
                           => operand_regs_9_port, Z => N3050);
   U969 : AO22D1 port map( A1 => coeff_memory_0_9, A2 => n673, B1 => n273, B2 
                           => operand_regs_233_port, Z => N2922);
   U970 : NAN2D1 port map( A1 => operand_regs_232_port, A2 => n673, Z => n145);
   U971 : NAN2D1 port map( A1 => operand_regs_231_port, A2 => n673, Z => n146);
   U972 : AO22D1 port map( A1 => n673, A2 => operand_regs_201_port, B1 => n271,
                           B2 => operand_regs_9_port, Z => N3210);
   U973 : AO22D1 port map( A1 => operand_regs_42_port, A2 => n277, B1 => 
                           coeff_memory_3_10, B2 => n673, Z => N3019);
   U974 : AO22D1 port map( A1 => operand_regs_106_port, A2 => n280, B1 => 
                           coeff_memory_2_10, B2 => n673, Z => N2987);
   U975 : AO22D1 port map( A1 => operand_regs_170_port, A2 => n282, B1 => 
                           coeff_memory_1_10, B2 => n673, Z => N2955);
   U976 : AO22D1 port map( A1 => coeff_memory_4_10, A2 => n673, B1 => n274, B2 
                           => operand_regs_10_port, Z => N3051);
   U977 : AO22D1 port map( A1 => coeff_memory_0_10, A2 => n673, B1 => n273, B2 
                           => operand_regs_234_port, Z => N2923);
   U978 : AO22D1 port map( A1 => n673, A2 => operand_regs_202_port, B1 => n271,
                           B2 => operand_regs_10_port, Z => N3211);
   U979 : OAI21M20D1 port map( A1 => operand_regs_73_port, A2 => n285, B => 
                           n144, Z => N3146);
   U980 : OAI21M20D1 port map( A1 => operand_regs_137_port, A2 => n284, B => 
                           n144, Z => N3114);
   U981 : OAI21M20D1 port map( A1 => n287, A2 => operand_regs_201_port, B => 
                           n144, Z => N3082);
   U982 : AO22D1 port map( A1 => operand_regs_43_port, A2 => n276, B1 => 
                           coeff_memory_3_11, B2 => n673, Z => N3020);
   U983 : AO22D1 port map( A1 => operand_regs_107_port, A2 => n280, B1 => 
                           coeff_memory_2_11, B2 => n673, Z => N2988);
   U984 : AO22D1 port map( A1 => operand_regs_171_port, A2 => n282, B1 => 
                           coeff_memory_1_11, B2 => n673, Z => N2956);
   U985 : AO22D1 port map( A1 => coeff_memory_4_11, A2 => n673, B1 => n271, B2 
                           => operand_regs_11_port, Z => N3052);
   U986 : AO22D1 port map( A1 => coeff_memory_0_11, A2 => n673, B1 => n273, B2 
                           => operand_regs_235_port, Z => N2924);
   U987 : AO22D1 port map( A1 => n673, A2 => operand_regs_204_port, B1 => n271,
                           B2 => operand_regs_12_port, Z => N3213);
   U988 : AO22D1 port map( A1 => n673, A2 => operand_regs_203_port, B1 => n271,
                           B2 => operand_regs_11_port, Z => N3212);
   U989 : NAN2D1 port map( A1 => operand_regs_233_port, A2 => n673, Z => n144);
   U990 : OAI21M20D1 port map( A1 => operand_regs_74_port, A2 => n285, B => 
                           n143, Z => N3147);
   U991 : OAI21M20D1 port map( A1 => operand_regs_138_port, A2 => n284, B => 
                           n143, Z => N3115);
   U992 : OAI21M20D1 port map( A1 => n287, A2 => operand_regs_202_port, B => 
                           n143, Z => N3083);
   U993 : AO22D1 port map( A1 => operand_regs_44_port, A2 => n281, B1 => 
                           coeff_memory_3_12, B2 => n673, Z => N3021);
   U994 : AO22D1 port map( A1 => operand_regs_108_port, A2 => n280, B1 => 
                           coeff_memory_2_12, B2 => n673, Z => N2989);
   U995 : AO22D1 port map( A1 => operand_regs_172_port, A2 => n282, B1 => 
                           coeff_memory_1_12, B2 => n673, Z => N2957);
   U996 : AO22D1 port map( A1 => coeff_memory_4_12, A2 => n673, B1 => n287, B2 
                           => operand_regs_12_port, Z => N3053);
   U997 : AO22D1 port map( A1 => coeff_memory_0_12, A2 => n673, B1 => n273, B2 
                           => operand_regs_236_port, Z => N2925);
   U998 : NAN2D1 port map( A1 => operand_regs_234_port, A2 => n673, Z => n143);
   U999 : OAI21M20D1 port map( A1 => operand_regs_75_port, A2 => n287, B => 
                           n142, Z => N3148);
   U1000 : OAI21M20D1 port map( A1 => operand_regs_139_port, A2 => n284, B => 
                           n142, Z => N3116);
   U1001 : OAI21M20D1 port map( A1 => operand_regs_76_port, A2 => n287, B => 
                           n141, Z => N3149);
   U1002 : OAI21M20D1 port map( A1 => operand_regs_140_port, A2 => n284, B => 
                           n141, Z => N3117);
   U1003 : OAI21M20D1 port map( A1 => n287, A2 => operand_regs_203_port, B => 
                           n142, Z => N3084);
   U1004 : OAI21M20D1 port map( A1 => n287, A2 => operand_regs_204_port, B => 
                           n141, Z => N3085);
   U1005 : AO22D1 port map( A1 => operand_regs_45_port, A2 => n276, B1 => 
                           coeff_memory_3_13, B2 => n673, Z => N3022);
   U1006 : AO22D1 port map( A1 => operand_regs_109_port, A2 => n280, B1 => 
                           coeff_memory_2_13, B2 => n673, Z => N2990);
   U1007 : AO22D1 port map( A1 => operand_regs_173_port, A2 => n282, B1 => 
                           coeff_memory_1_13, B2 => n673, Z => N2958);
   U1008 : AO22D1 port map( A1 => coeff_memory_4_13, A2 => n673, B1 => n275, B2
                           => operand_regs_13_port, Z => N3054);
   U1009 : AO22D1 port map( A1 => coeff_memory_0_13, A2 => n673, B1 => n273, B2
                           => operand_regs_237_port, Z => N2926);
   U1010 : NAN2D1 port map( A1 => operand_regs_235_port, A2 => n673, Z => n142)
                           ;
   U1011 : NAN2D1 port map( A1 => operand_regs_236_port, A2 => n673, Z => n141)
                           ;
   U1012 : AO22D1 port map( A1 => n673, A2 => operand_regs_205_port, B1 => n287
                           , B2 => operand_regs_13_port, Z => N3214);
   U1013 : AO22D1 port map( A1 => n673, A2 => operand_regs_206_port, B1 => n271
                           , B2 => operand_regs_14_port, Z => N3215);
   U1014 : AO22D1 port map( A1 => operand_regs_46_port, A2 => n278, B1 => 
                           coeff_memory_3_14, B2 => n673, Z => N3023);
   U1015 : AO22D1 port map( A1 => operand_regs_110_port, A2 => n279, B1 => 
                           coeff_memory_2_14, B2 => n673, Z => N2991);
   U1016 : AO22D1 port map( A1 => operand_regs_174_port, A2 => n282, B1 => 
                           coeff_memory_1_14, B2 => n673, Z => N2959);
   U1017 : AO22D1 port map( A1 => coeff_memory_4_14, A2 => n673, B1 => n276, B2
                           => operand_regs_14_port, Z => N3055);
   U1018 : AO22D1 port map( A1 => coeff_memory_0_14, A2 => n673, B1 => n287, B2
                           => operand_regs_238_port, Z => N2927);
   U1019 : OAI21M20D1 port map( A1 => operand_regs_77_port, A2 => n287, B => 
                           n140, Z => N3150);
   U1020 : OAI21M20D1 port map( A1 => operand_regs_141_port, A2 => n284, B => 
                           n140, Z => N3118);
   U1021 : OAI21M20D1 port map( A1 => operand_regs_78_port, A2 => n287, B => 
                           n139, Z => N3151);
   U1022 : OAI21M20D1 port map( A1 => operand_regs_142_port, A2 => n284, B => 
                           n139, Z => N3119);
   U1023 : OAI21M20D1 port map( A1 => n287, A2 => operand_regs_205_port, B => 
                           n140, Z => N3086);
   U1024 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_206_port, B => 
                           n139, Z => N3087);
   U1025 : AO22D1 port map( A1 => operand_regs_47_port, A2 => n278, B1 => 
                           coeff_memory_3_15, B2 => n673, Z => N3024);
   U1026 : AO22D1 port map( A1 => operand_regs_111_port, A2 => n277, B1 => 
                           coeff_memory_2_15, B2 => n673, Z => N2992);
   U1027 : AO22D1 port map( A1 => operand_regs_175_port, A2 => n278, B1 => 
                           coeff_memory_1_15, B2 => n673, Z => N2960);
   U1028 : AO22D1 port map( A1 => n673, A2 => operand_regs_207_port, B1 => n272
                           , B2 => operand_regs_15_port, Z => N3216);
   U1029 : AO22D1 port map( A1 => coeff_memory_4_15, A2 => n673, B1 => n275, B2
                           => operand_regs_15_port, Z => N3056);
   U1030 : AO22D1 port map( A1 => coeff_memory_0_15, A2 => n673, B1 => n287, B2
                           => operand_regs_239_port, Z => N2928);
   U1031 : NAN2D1 port map( A1 => operand_regs_237_port, A2 => n673, Z => n140)
                           ;
   U1032 : NAN2D1 port map( A1 => operand_regs_238_port, A2 => n673, Z => n139)
                           ;
   U1033 : OAI21M20D1 port map( A1 => operand_regs_79_port, A2 => n287, B => 
                           n138, Z => N3152);
   U1034 : OAI21M20D1 port map( A1 => operand_regs_143_port, A2 => n284, B => 
                           n138, Z => N3120);
   U1035 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_207_port, B => 
                           n138, Z => N3088);
   U1036 : AO22D1 port map( A1 => operand_regs_48_port, A2 => n281, B1 => 
                           coeff_memory_3_16, B2 => n673, Z => N3025);
   U1037 : AO22D1 port map( A1 => operand_regs_112_port, A2 => n277, B1 => 
                           coeff_memory_2_16, B2 => n673, Z => N2993);
   U1038 : AO22D1 port map( A1 => operand_regs_176_port, A2 => n282, B1 => 
                           coeff_memory_1_16, B2 => n673, Z => N2961);
   U1039 : AO22D1 port map( A1 => coeff_memory_4_16, A2 => n673, B1 => n276, B2
                           => operand_regs_16_port, Z => N3057);
   U1040 : AO22D1 port map( A1 => coeff_memory_0_16, A2 => n673, B1 => n287, B2
                           => operand_regs_240_port, Z => N2929);
   U1041 : AO22D1 port map( A1 => n673, A2 => operand_regs_208_port, B1 => n271
                           , B2 => operand_regs_16_port, Z => N3217);
   U1042 : NAN2D1 port map( A1 => operand_regs_239_port, A2 => n673, Z => n138)
                           ;
   U1043 : AO22D1 port map( A1 => operand_regs_49_port, A2 => n281, B1 => 
                           coeff_memory_3_17, B2 => n673, Z => N3026);
   U1044 : AO22D1 port map( A1 => operand_regs_113_port, A2 => n277, B1 => 
                           coeff_memory_2_17, B2 => n673, Z => N2994);
   U1045 : AO22D1 port map( A1 => operand_regs_177_port, A2 => n282, B1 => 
                           coeff_memory_1_17, B2 => n673, Z => N2962);
   U1046 : AO22D1 port map( A1 => coeff_memory_4_17, A2 => n673, B1 => n276, B2
                           => operand_regs_17_port, Z => N3058);
   U1047 : AO22D1 port map( A1 => coeff_memory_0_17, A2 => n673, B1 => n287, B2
                           => operand_regs_241_port, Z => N2930);
   U1048 : OAI21M20D1 port map( A1 => operand_regs_80_port, A2 => n287, B => 
                           n137, Z => N3153);
   U1049 : OAI21M20D1 port map( A1 => operand_regs_144_port, A2 => n284, B => 
                           n137, Z => N3121);
   U1050 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_208_port, B => 
                           n137, Z => N3089);
   U1051 : AO22D1 port map( A1 => operand_regs_50_port, A2 => n281, B1 => 
                           coeff_memory_3_18, B2 => n673, Z => N3027);
   U1052 : AO22D1 port map( A1 => operand_regs_114_port, A2 => n277, B1 => 
                           coeff_memory_2_18, B2 => n673, Z => N2995);
   U1053 : AO22D1 port map( A1 => operand_regs_178_port, A2 => n282, B1 => 
                           coeff_memory_1_18, B2 => n673, Z => N2963);
   U1054 : AO22D1 port map( A1 => coeff_memory_4_18, A2 => n673, B1 => n275, B2
                           => operand_regs_18_port, Z => N3059);
   U1055 : AO22D1 port map( A1 => coeff_memory_0_18, A2 => n673, B1 => n283, B2
                           => operand_regs_242_port, Z => N2931);
   U1056 : AO22D1 port map( A1 => n673, A2 => operand_regs_209_port, B1 => n272
                           , B2 => operand_regs_17_port, Z => N3218);
   U1057 : AO22D1 port map( A1 => operand_regs_51_port, A2 => n281, B1 => 
                           coeff_memory_3_19, B2 => n673, Z => N3028);
   U1058 : AO22D1 port map( A1 => operand_regs_115_port, A2 => n277, B1 => 
                           coeff_memory_2_19, B2 => n673, Z => N2996);
   U1059 : AO22D1 port map( A1 => operand_regs_179_port, A2 => n282, B1 => 
                           coeff_memory_1_19, B2 => n673, Z => N2964);
   U1060 : NAN2D1 port map( A1 => operand_regs_240_port, A2 => n673, Z => n137)
                           ;
   U1061 : AO22D1 port map( A1 => coeff_memory_0_19, A2 => n673, B1 => n274, B2
                           => operand_regs_243_port, Z => N2932);
   U1062 : AO22D1 port map( A1 => coeff_memory_4_19, A2 => n673, B1 => n276, B2
                           => operand_regs_19_port, Z => N3060);
   U1063 : OAI21M20D1 port map( A1 => operand_regs_81_port, A2 => n287, B => 
                           n136, Z => N3154);
   U1064 : OAI21M20D1 port map( A1 => operand_regs_145_port, A2 => n284, B => 
                           n136, Z => N3122);
   U1065 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_209_port, B => 
                           n136, Z => N3090);
   U1066 : AO22D1 port map( A1 => n673, A2 => operand_regs_210_port, B1 => n271
                           , B2 => operand_regs_18_port, Z => N3219);
   U1067 : NAN2D1 port map( A1 => operand_regs_241_port, A2 => n673, Z => n136)
                           ;
   U1068 : OAI21M20D1 port map( A1 => operand_regs_82_port, A2 => n282, B => 
                           n135, Z => N3155);
   U1069 : OAI21M20D1 port map( A1 => operand_regs_146_port, A2 => n287, B => 
                           n135, Z => N3123);
   U1070 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_210_port, B => 
                           n135, Z => N3091);
   U1071 : AO22D1 port map( A1 => n673, A2 => operand_regs_211_port, B1 => n277
                           , B2 => operand_regs_19_port, Z => N3220);
   U1072 : AO22D1 port map( A1 => n673, A2 => operand_regs_212_port, B1 => n271
                           , B2 => operand_regs_20_port, Z => N3221);
   U1073 : AO22D1 port map( A1 => operand_regs_52_port, A2 => n281, B1 => 
                           coeff_memory_3_20, B2 => n673, Z => N3029);
   U1074 : AO22D1 port map( A1 => operand_regs_116_port, A2 => n277, B1 => 
                           coeff_memory_2_20, B2 => n673, Z => N2997);
   U1075 : AO22D1 port map( A1 => operand_regs_180_port, A2 => n282, B1 => 
                           coeff_memory_1_20, B2 => n673, Z => N2965);
   U1076 : AO22D1 port map( A1 => coeff_memory_4_20, A2 => n673, B1 => n276, B2
                           => operand_regs_20_port, Z => N3061);
   U1077 : AO22D1 port map( A1 => coeff_memory_0_20, A2 => n673, B1 => n274, B2
                           => operand_regs_244_port, Z => N2933);
   U1078 : NAN2D1 port map( A1 => operand_regs_242_port, A2 => n673, Z => n135)
                           ;
   U1079 : OAI21M20D1 port map( A1 => operand_regs_83_port, A2 => n287, B => 
                           n134, Z => N3156);
   U1080 : OAI21M20D1 port map( A1 => operand_regs_147_port, A2 => n287, B => 
                           n134, Z => N3124);
   U1081 : OAI21M20D1 port map( A1 => operand_regs_84_port, A2 => n283, B => 
                           n133, Z => N3157);
   U1082 : OAI21M20D1 port map( A1 => operand_regs_148_port, A2 => n277, B => 
                           n133, Z => N3125);
   U1083 : AO22D1 port map( A1 => operand_regs_53_port, A2 => n281, B1 => 
                           coeff_memory_3_21, B2 => n673, Z => N3030);
   U1084 : AO22D1 port map( A1 => operand_regs_117_port, A2 => n277, B1 => 
                           coeff_memory_2_21, B2 => n673, Z => N2998);
   U1085 : AO22D1 port map( A1 => operand_regs_181_port, A2 => n279, B1 => 
                           coeff_memory_1_21, B2 => n673, Z => N2966);
   U1086 : OAI21M20D1 port map( A1 => n287, A2 => operand_regs_211_port, B => 
                           n134, Z => N3092);
   U1087 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_212_port, B => 
                           n133, Z => N3093);
   U1088 : AO22D1 port map( A1 => coeff_memory_4_21, A2 => n673, B1 => n275, B2
                           => operand_regs_21_port, Z => N3062);
   U1089 : AO22D1 port map( A1 => coeff_memory_0_21, A2 => n673, B1 => n274, B2
                           => operand_regs_245_port, Z => N2934);
   U1090 : NAN2D1 port map( A1 => operand_regs_243_port, A2 => n673, Z => n134)
                           ;
   U1091 : NAN2D1 port map( A1 => operand_regs_244_port, A2 => n673, Z => n133)
                           ;
   U1092 : AO22D1 port map( A1 => n673, A2 => operand_regs_213_port, B1 => n273
                           , B2 => operand_regs_21_port, Z => N3222);
   U1093 : AO22D1 port map( A1 => n673, A2 => operand_regs_214_port, B1 => n273
                           , B2 => operand_regs_22_port, Z => N3223);
   U1094 : AO22D1 port map( A1 => operand_regs_54_port, A2 => n283, B1 => 
                           coeff_memory_3_22, B2 => n673, Z => N3031);
   U1095 : AO22D1 port map( A1 => operand_regs_118_port, A2 => n277, B1 => 
                           coeff_memory_2_22, B2 => n673, Z => N2999);
   U1096 : AO22D1 port map( A1 => operand_regs_182_port, A2 => n279, B1 => 
                           coeff_memory_1_22, B2 => n673, Z => N2967);
   U1097 : AO22D1 port map( A1 => coeff_memory_4_22, A2 => n673, B1 => n275, B2
                           => operand_regs_22_port, Z => N3063);
   U1098 : AO22D1 port map( A1 => coeff_memory_0_22, A2 => n673, B1 => n274, B2
                           => operand_regs_246_port, Z => N2935);
   U1099 : OAI21M20D1 port map( A1 => operand_regs_85_port, A2 => n282, B => 
                           n132, Z => N3158);
   U1100 : OAI21M20D1 port map( A1 => operand_regs_149_port, A2 => n287, B => 
                           n132, Z => N3126);
   U1101 : OAI21M20D1 port map( A1 => operand_regs_86_port, A2 => n287, B => 
                           n131, Z => N3159);
   U1102 : OAI21M20D1 port map( A1 => operand_regs_150_port, A2 => n283, B => 
                           n131, Z => N3127);
   U1103 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_213_port, B => 
                           n132, Z => N3094);
   U1104 : OAI21M20D1 port map( A1 => n286, A2 => operand_regs_214_port, B => 
                           n131, Z => N3095);
   U1105 : AO22D1 port map( A1 => operand_regs_55_port, A2 => n283, B1 => 
                           coeff_memory_3_23, B2 => n673, Z => N3032);
   U1106 : AO22D1 port map( A1 => operand_regs_119_port, A2 => n277, B1 => 
                           coeff_memory_2_23, B2 => n673, Z => N3000);
   U1107 : AO22D1 port map( A1 => operand_regs_183_port, A2 => n279, B1 => 
                           coeff_memory_1_23, B2 => n673, Z => N2968);
   U1108 : AO22D1 port map( A1 => coeff_memory_4_23, A2 => n673, B1 => n275, B2
                           => operand_regs_23_port, Z => N3064);
   U1109 : AO22D1 port map( A1 => coeff_memory_0_23, A2 => n673, B1 => n274, B2
                           => operand_regs_247_port, Z => N2936);
   U1110 : AO22D1 port map( A1 => n673, A2 => operand_regs_215_port, B1 => n287
                           , B2 => operand_regs_23_port, Z => N3224);
   U1111 : NAN2D1 port map( A1 => operand_regs_245_port, A2 => n673, Z => n132)
                           ;
   U1112 : NAN2D1 port map( A1 => operand_regs_246_port, A2 => n673, Z => n131)
                           ;
   U1113 : OAI21M20D1 port map( A1 => operand_regs_87_port, A2 => n283, B => 
                           n130, Z => N3160);
   U1114 : OAI21M20D1 port map( A1 => operand_regs_151_port, A2 => n287, B => 
                           n130, Z => N3128);
   U1115 : OAI21M20D1 port map( A1 => n283, A2 => operand_regs_215_port, B => 
                           n130, Z => N3096);
   U1116 : AO22D1 port map( A1 => operand_regs_56_port, A2 => n283, B1 => 
                           coeff_memory_3_24, B2 => n673, Z => N3033);
   U1117 : AO22D1 port map( A1 => operand_regs_120_port, A2 => n277, B1 => 
                           coeff_memory_2_24, B2 => n673, Z => N3001);
   U1118 : AO22D1 port map( A1 => operand_regs_184_port, A2 => n279, B1 => 
                           coeff_memory_1_24, B2 => n673, Z => N2969);
   U1119 : AO22D1 port map( A1 => n673, A2 => operand_regs_216_port, B1 => n273
                           , B2 => operand_regs_24_port, Z => N3225);
   U1120 : AO22D1 port map( A1 => coeff_memory_4_24, A2 => n673, B1 => n287, B2
                           => operand_regs_24_port, Z => N3065);
   U1121 : AO22D1 port map( A1 => coeff_memory_0_24, A2 => n673, B1 => n274, B2
                           => operand_regs_248_port, Z => N2937);
   U1122 : NAN2D1 port map( A1 => operand_regs_247_port, A2 => n673, Z => n130)
                           ;
   U1123 : OAI21M20D1 port map( A1 => operand_regs_88_port, A2 => n282, B => 
                           n129, Z => N3161);
   U1124 : OAI21M20D1 port map( A1 => operand_regs_152_port, A2 => n287, B => 
                           n129, Z => N3129);
   U1125 : OAI21M20D1 port map( A1 => n287, A2 => operand_regs_216_port, B => 
                           n129, Z => N3097);
   U1126 : AO22D1 port map( A1 => operand_regs_57_port, A2 => n283, B1 => 
                           coeff_memory_3_25, B2 => n673, Z => N3034);
   U1127 : AO22D1 port map( A1 => operand_regs_121_port, A2 => n277, B1 => 
                           coeff_memory_2_25, B2 => n673, Z => N3002);
   U1128 : AO22D1 port map( A1 => operand_regs_185_port, A2 => n279, B1 => 
                           coeff_memory_1_25, B2 => n673, Z => N2970);
   U1129 : AO22D1 port map( A1 => coeff_memory_4_25, A2 => n673, B1 => n277, B2
                           => operand_regs_25_port, Z => N3066);
   U1130 : AO22D1 port map( A1 => coeff_memory_0_25, A2 => n673, B1 => n274, B2
                           => operand_regs_249_port, Z => N2938);
   U1131 : AO22D1 port map( A1 => n673, A2 => operand_regs_217_port, B1 => n283
                           , B2 => operand_regs_25_port, Z => N3226);
   U1132 : NAN2D1 port map( A1 => operand_regs_248_port, A2 => n673, Z => n129)
                           ;
   U1133 : OAI21M20D1 port map( A1 => operand_regs_89_port, A2 => n277, B => 
                           n128, Z => N3162);
   U1134 : OAI21M20D1 port map( A1 => operand_regs_153_port, A2 => n287, B => 
                           n128, Z => N3130);
   U1135 : OAI21M20D1 port map( A1 => n282, A2 => operand_regs_217_port, B => 
                           n128, Z => N3098);
   U1136 : AO22D1 port map( A1 => operand_regs_58_port, A2 => n283, B1 => 
                           coeff_memory_3_26, B2 => n673, Z => N3035);
   U1137 : AO22D1 port map( A1 => operand_regs_122_port, A2 => n276, B1 => 
                           coeff_memory_2_26, B2 => n673, Z => N3003);
   U1138 : AO22D1 port map( A1 => operand_regs_186_port, A2 => n279, B1 => 
                           coeff_memory_1_26, B2 => n673, Z => N2971);
   U1139 : AO22D1 port map( A1 => coeff_memory_4_26, A2 => n673, B1 => n283, B2
                           => operand_regs_26_port, Z => N3067);
   U1140 : AO22D1 port map( A1 => coeff_memory_0_26, A2 => n673, B1 => n287, B2
                           => operand_regs_250_port, Z => N2939);
   U1141 : AO22D1 port map( A1 => n673, A2 => operand_regs_218_port, B1 => n273
                           , B2 => operand_regs_26_port, Z => N3227);
   U1142 : NAN2D1 port map( A1 => operand_regs_249_port, A2 => n673, Z => n128)
                           ;
   U1143 : AO22D1 port map( A1 => operand_regs_59_port, A2 => n283, B1 => 
                           coeff_memory_3_27, B2 => n673, Z => N3036);
   U1144 : AO22D1 port map( A1 => operand_regs_123_port, A2 => n278, B1 => 
                           coeff_memory_2_27, B2 => n673, Z => N3004);
   U1145 : AO22D1 port map( A1 => operand_regs_187_port, A2 => n279, B1 => 
                           coeff_memory_1_27, B2 => n673, Z => N2972);
   U1146 : OAI21M20D1 port map( A1 => operand_regs_90_port, A2 => n287, B => 
                           n127, Z => N3163);
   U1147 : OAI21M20D1 port map( A1 => operand_regs_154_port, A2 => n287, B => 
                           n127, Z => N3131);
   U1148 : OAI21M20D1 port map( A1 => n283, A2 => operand_regs_218_port, B => 
                           n127, Z => N3099);
   U1149 : AO22D1 port map( A1 => coeff_memory_4_27, A2 => n673, B1 => n287, B2
                           => operand_regs_27_port, Z => N3068);
   U1150 : AO22D1 port map( A1 => coeff_memory_0_27, A2 => n673, B1 => n283, B2
                           => operand_regs_251_port, Z => N2940);
   U1151 : AO22D1 port map( A1 => operand_regs_60_port, A2 => n283, B1 => 
                           coeff_memory_3_28, B2 => n673, Z => N3037);
   U1152 : AO22D1 port map( A1 => operand_regs_124_port, A2 => n278, B1 => 
                           coeff_memory_2_28, B2 => n673, Z => N3005);
   U1153 : AO22D1 port map( A1 => operand_regs_188_port, A2 => n279, B1 => 
                           coeff_memory_1_28, B2 => n673, Z => N2973);
   U1154 : NAN2D1 port map( A1 => operand_regs_250_port, A2 => n673, Z => n127)
                           ;
   U1155 : AO22D1 port map( A1 => n673, A2 => operand_regs_219_port, B1 => n277
                           , B2 => operand_regs_27_port, Z => N3228);
   U1156 : AO22D1 port map( A1 => coeff_memory_4_28, A2 => n673, B1 => n283, B2
                           => operand_regs_28_port, Z => N3069);
   U1157 : AO22D1 port map( A1 => coeff_memory_0_28, A2 => n673, B1 => n282, B2
                           => operand_regs_252_port, Z => N2941);
   U1158 : OAI21M20D1 port map( A1 => operand_regs_91_port, A2 => n283, B => 
                           n126, Z => N3164);
   U1159 : OAI21M20D1 port map( A1 => operand_regs_155_port, A2 => n283, B => 
                           n126, Z => N3132);
   U1160 : AO22D1 port map( A1 => operand_regs_61_port, A2 => n283, B1 => 
                           coeff_memory_3_29, B2 => n673, Z => N3038);
   U1161 : AO22D1 port map( A1 => operand_regs_125_port, A2 => n278, B1 => 
                           coeff_memory_2_29, B2 => n673, Z => N3006);
   U1162 : AO22D1 port map( A1 => operand_regs_189_port, A2 => n279, B1 => 
                           coeff_memory_1_29, B2 => n673, Z => N2974);
   U1163 : OAI21M20D1 port map( A1 => n287, A2 => operand_regs_219_port, B => 
                           n126, Z => N3100);
   U1164 : AO22D1 port map( A1 => coeff_memory_4_29, A2 => n673, B1 => n287, B2
                           => operand_regs_29_port, Z => N3070);
   U1165 : AO22D1 port map( A1 => coeff_memory_0_29, A2 => n673, B1 => n287, B2
                           => operand_regs_253_port, Z => N2942);
   U1166 : AO22D1 port map( A1 => n673, A2 => operand_regs_220_port, B1 => n273
                           , B2 => operand_regs_28_port, Z => N3229);
   U1167 : NAN2D1 port map( A1 => operand_regs_251_port, A2 => n673, Z => n126)
                           ;
   U1168 : OAI21M20D1 port map( A1 => operand_regs_92_port, A2 => n287, B => 
                           n125, Z => N3165);
   U1169 : OAI21M20D1 port map( A1 => operand_regs_156_port, A2 => n277, B => 
                           n125, Z => N3133);
   U1170 : OAI21M20D1 port map( A1 => n283, A2 => operand_regs_220_port, B => 
                           n125, Z => N3101);
   U1171 : AO22D1 port map( A1 => operand_regs_62_port, A2 => n283, B1 => 
                           coeff_memory_3_30, B2 => n673, Z => N3039);
   U1172 : AO22D1 port map( A1 => operand_regs_126_port, A2 => n278, B1 => 
                           coeff_memory_2_30, B2 => n673, Z => N3007);
   U1173 : AO22D1 port map( A1 => operand_regs_190_port, A2 => n279, B1 => 
                           coeff_memory_1_30, B2 => n673, Z => N2975);
   U1174 : NAN2D1 port map( A1 => operand_regs_252_port, A2 => n673, Z => n125)
                           ;
   U1175 : AO22D1 port map( A1 => coeff_memory_4_30, A2 => n673, B1 => n282, B2
                           => operand_regs_30_port, Z => N3071);
   U1176 : AO22D1 port map( A1 => coeff_memory_0_30, A2 => n673, B1 => n283, B2
                           => operand_regs_254_port, Z => N2943);
   U1177 : AO22D1 port map( A1 => n673, A2 => operand_regs_221_port, B1 => n272
                           , B2 => operand_regs_29_port, Z => N3230);
   U1178 : AO22D1 port map( A1 => n673, A2 => operand_regs_222_port, B1 => n283
                           , B2 => operand_regs_30_port, Z => N3231);
   U1179 : OAI21M20D1 port map( A1 => operand_regs_93_port, A2 => n287, B => 
                           n124, Z => N3166);
   U1180 : OAI21M20D1 port map( A1 => operand_regs_157_port, A2 => n287, B => 
                           n124, Z => N3134);
   U1181 : OAI21M20D1 port map( A1 => operand_regs_94_port, A2 => n283, B => 
                           n123, Z => N3167);
   U1182 : OAI21M20D1 port map( A1 => operand_regs_158_port, A2 => n287, B => 
                           n123, Z => N3135);
   U1183 : OAI21M20D1 port map( A1 => n277, A2 => operand_regs_221_port, B => 
                           n124, Z => N3102);
   U1184 : OAI21M20D1 port map( A1 => n283, A2 => operand_regs_222_port, B => 
                           n123, Z => N3103);
   U1185 : AO22D1 port map( A1 => operand_regs_63_port, A2 => n283, B1 => 
                           coeff_memory_3_31, B2 => n673, Z => N3040);
   U1186 : AO22D1 port map( A1 => operand_regs_127_port, A2 => n280, B1 => 
                           coeff_memory_2_31, B2 => n673, Z => N3008);
   U1187 : AO22D1 port map( A1 => operand_regs_191_port, A2 => n279, B1 => 
                           coeff_memory_1_31, B2 => n673, Z => N2976);
   U1188 : AO22D1 port map( A1 => coeff_memory_4_31, A2 => n673, B1 => n287, B2
                           => operand_regs_31_port, Z => N3072);
   U1189 : AO22D1 port map( A1 => coeff_memory_0_31, A2 => n673, B1 => n282, B2
                           => operand_regs_255_port, Z => N2944);
   U1190 : NAN2D1 port map( A1 => operand_regs_253_port, A2 => n673, Z => n124)
                           ;
   U1191 : NAN2D1 port map( A1 => operand_regs_254_port, A2 => n673, Z => n123)
                           ;
   U1192 : OAI21M20D1 port map( A1 => operand_regs_95_port, A2 => n284, B => 
                           n122, Z => N3168);
   U1193 : OAI21M20D1 port map( A1 => operand_regs_159_port, A2 => n287, B => 
                           n122, Z => N3136);
   U1194 : OAI21M20D1 port map( A1 => n287, A2 => operand_regs_223_port, B => 
                           n122, Z => N3104);
   U1195 : AO22D1 port map( A1 => n673, A2 => operand_regs_223_port, B1 => n275
                           , B2 => operand_regs_31_port, Z => N3232);
   U1196 : NAN2D1 port map( A1 => operand_regs_255_port, A2 => n673, Z => n122)
                           ;
   U1197 : AO22D1 port map( A1 => N2876, A2 => n672, B1 => N2859, B2 => n696, Z
                           => N2894);
   U1198 : AO22D1 port map( A1 => N2875, A2 => n672, B1 => N2858, B2 => n696, Z
                           => N2895);
   U1199 : AO22D1 port map( A1 => N2874, A2 => n672, B1 => N2857, B2 => n696, Z
                           => N2896);
   U1200 : AO22D1 port map( A1 => N2873, A2 => n672, B1 => N2856, B2 => n696, Z
                           => N2897);
   U1201 : AO22D1 port map( A1 => N2872, A2 => n672, B1 => N2855, B2 => n696, Z
                           => N2898);
   U1202 : AO22D1 port map( A1 => N2871, A2 => n672, B1 => N2854, B2 => n696, Z
                           => N2899);
   U1203 : AO22D1 port map( A1 => N2870, A2 => n672, B1 => N2853, B2 => n696, Z
                           => N2900);
   U1204 : AO22D1 port map( A1 => N2869, A2 => n672, B1 => N2852, B2 => n696, Z
                           => N2901);
   U1205 : AO22D1 port map( A1 => N2868, A2 => n672, B1 => N2851, B2 => n696, Z
                           => N2902);
   U1206 : AO22D1 port map( A1 => N2867, A2 => n672, B1 => N2850, B2 => n696, Z
                           => N2903);
   U1207 : AO22D1 port map( A1 => N2881, A2 => n672, B1 => N2864, B2 => n696, Z
                           => N2889);
   U1208 : AO22D1 port map( A1 => N2880, A2 => n672, B1 => N2863, B2 => n696, Z
                           => N2890);
   U1209 : AO22D1 port map( A1 => N2879, A2 => n672, B1 => N2862, B2 => n696, Z
                           => N2891);
   U1210 : AO22D1 port map( A1 => N2878, A2 => n672, B1 => N2861, B2 => n696, Z
                           => N2892);
   U1211 : AO22D1 port map( A1 => N2877, A2 => n672, B1 => N2860, B2 => n696, Z
                           => N2893);
   U1212 : AO22D1 port map( A1 => N2882, A2 => n672, B1 => N2865, B2 => n696, Z
                           => N2888);
   U1213 : INVD1 port map( A => N64, Z => n671);
   U1214 : INVD1 port map( A => coeff_load, Z => n686);
   U1215 : NOR2D1 port map( A1 => n684, A2 => out_busy, Z => n79);
   U1216 : NAN3D1 port map( A1 => n81, A2 => out_busy, A3 => N62, Z => n4);
   U1217 : INVD1 port map( A => N62, Z => n694);
   U1218 : BUFD1 port map( A => odd1, Z => n672);
   U1219 : INVD1 port map( A => out_busy, Z => n695);
   U1220 : INVD1 port map( A => odd, Z => n687);
   U1221 : NAN3D1 port map( A1 => in_counter_1_port, A2 => in_busy, A3 => 
                           in_counter_0_port, Z => n88);
   U1222 : NOR2D1 port map( A1 => n690, A2 => in_counter_0_port, Z => n155);
   U1223 : OAI21M20D1 port map( A1 => n690, A2 => in_trigger, B => n100, Z => 
                           n84);
   U1224 : INVD1 port map( A => in_busy, Z => n690);
   U1225 : INVD1 port map( A => in_counter_2_port, Z => n693);
   U1226 : INVD1 port map( A => N63, Z => n697);
   U1227 : NOR2D1 port map( A1 => n688, A2 => in_counter_1_port, Z => n119);
   U1228 : NAN2D1 port map( A1 => in_counter_1_port, A2 => n155, Z => n85);
   U1229 : AND3D1 port map( A1 => in_counter_0_port, A2 => in_busy, A3 => n692,
                           Z => n87);
   U1230 : INVD1 port map( A => in_counter_1_port, Z => n692);
   U1231 : NAN2D1 port map( A1 => n78, A2 => n672, Z => n77);
   U1232 : NOR2D1 port map( A1 => n687, A2 => in_counter_2_port, Z => n101);
   U1233 : NOR2D1 port map( A1 => n693, A2 => odd, Z => n115);
   U1234 : NOR2D1 port map( A1 => odd, A2 => in_counter_2_port, Z => n120);
   U1235 : INVD1 port map( A => out_trigger, Z => n685);
   U1236 : NOR2D1 port map( A1 => n522, A2 => avs_addr(1), Z => n288);
   U1237 : NOR2D1 port map( A1 => n522, A2 => n680, Z => n289);
   U1238 : AOI22D1 port map( A1 => in_buf_64_port, A2 => n266, B1 => 
                           in_buf_0_port, B2 => n242, Z => n295);
   U1239 : NOR2D1 port map( A1 => avs_addr(1), A2 => avs_addr(2), Z => n290);
   U1240 : AND2D1 port map( A1 => n290, A2 => avs_addr(0), Z => n514);
   U1241 : NOR2D1 port map( A1 => n680, A2 => avs_addr(2), Z => n291);
   U1242 : AND2D1 port map( A1 => n291, A2 => avs_addr(0), Z => n513);
   U1243 : AOI22D1 port map( A1 => in_buf_192_port, A2 => n527, B1 => 
                           in_buf_128_port, B2 => n525, Z => n294);
   U1244 : NOR2M1D1 port map( A1 => n288, A2 => avs_addr(0), Z => n516);
   U1245 : NOR2M1D1 port map( A1 => n289, A2 => avs_addr(0), Z => n515);
   U1246 : AOI22D1 port map( A1 => in_buf_96_port, A2 => n529, B1 => 
                           in_buf_32_port, B2 => n515, Z => n293);
   U1247 : NOR2M1D1 port map( A1 => n290, A2 => avs_addr(0), Z => n518);
   U1248 : NOR2M1D1 port map( A1 => n291, A2 => avs_addr(0), Z => n517);
   U1249 : AOI22D1 port map( A1 => in_buf_224_port, A2 => n534, B1 => 
                           in_buf_160_port, B2 => n532, Z => n292);
   U1250 : NAN4D1 port map( A1 => n295, A2 => n294, A3 => n293, A4 => n292, Z 
                           => N2041);
   U1251 : AOI22D1 port map( A1 => in_buf_65_port, A2 => n266, B1 => 
                           in_buf_1_port, B2 => n242, Z => n299);
   U1252 : AOI22D1 port map( A1 => in_buf_193_port, A2 => n527, B1 => 
                           in_buf_129_port, B2 => n513, Z => n298);
   U1253 : AOI22D1 port map( A1 => in_buf_97_port, A2 => n529, B1 => 
                           in_buf_33_port, B2 => n515, Z => n297);
   U1254 : AOI22D1 port map( A1 => in_buf_225_port, A2 => n518, B1 => 
                           in_buf_161_port, B2 => n517, Z => n296);
   U1255 : NAN4D1 port map( A1 => n299, A2 => n298, A3 => n297, A4 => n296, Z 
                           => N2040);
   U1256 : AOI22D1 port map( A1 => in_buf_66_port, A2 => n266, B1 => 
                           in_buf_2_port, B2 => n242, Z => n303);
   U1257 : AOI22D1 port map( A1 => in_buf_194_port, A2 => n527, B1 => 
                           in_buf_130_port, B2 => n513, Z => n302);
   U1258 : AOI22D1 port map( A1 => in_buf_98_port, A2 => n529, B1 => 
                           in_buf_34_port, B2 => n515, Z => n301);
   U1259 : AOI22D1 port map( A1 => in_buf_226_port, A2 => n518, B1 => 
                           in_buf_162_port, B2 => n517, Z => n300);
   U1260 : NAN4D1 port map( A1 => n303, A2 => n302, A3 => n301, A4 => n300, Z 
                           => N2039);
   U1261 : AOI22D1 port map( A1 => in_buf_67_port, A2 => n266, B1 => 
                           in_buf_3_port, B2 => n242, Z => n307);
   U1262 : AOI22D1 port map( A1 => in_buf_195_port, A2 => n527, B1 => 
                           in_buf_131_port, B2 => n513, Z => n306);
   U1263 : AOI22D1 port map( A1 => in_buf_99_port, A2 => n529, B1 => 
                           in_buf_35_port, B2 => n515, Z => n305);
   U1264 : AOI22D1 port map( A1 => in_buf_227_port, A2 => n518, B1 => 
                           in_buf_163_port, B2 => n517, Z => n304);
   U1265 : NAN4D1 port map( A1 => n307, A2 => n306, A3 => n305, A4 => n304, Z 
                           => N2038);
   U1266 : AOI22D1 port map( A1 => in_buf_68_port, A2 => n266, B1 => 
                           in_buf_4_port, B2 => n242, Z => n311);
   U1267 : AOI22D1 port map( A1 => in_buf_196_port, A2 => n527, B1 => 
                           in_buf_132_port, B2 => n513, Z => n310);
   U1268 : AOI22D1 port map( A1 => in_buf_100_port, A2 => n529, B1 => 
                           in_buf_36_port, B2 => n515, Z => n309);
   U1269 : AOI22D1 port map( A1 => in_buf_228_port, A2 => n518, B1 => 
                           in_buf_164_port, B2 => n517, Z => n308);
   U1270 : NAN4D1 port map( A1 => n311, A2 => n310, A3 => n309, A4 => n308, Z 
                           => N2037);
   U1271 : AOI22D1 port map( A1 => in_buf_69_port, A2 => n266, B1 => 
                           in_buf_5_port, B2 => n242, Z => n315);
   U1272 : AOI22D1 port map( A1 => in_buf_197_port, A2 => n527, B1 => 
                           in_buf_133_port, B2 => n513, Z => n314);
   U1273 : AOI22D1 port map( A1 => in_buf_101_port, A2 => n529, B1 => 
                           in_buf_37_port, B2 => n515, Z => n313);
   U1274 : AOI22D1 port map( A1 => in_buf_229_port, A2 => n518, B1 => 
                           in_buf_165_port, B2 => n517, Z => n312);
   U1275 : NAN4D1 port map( A1 => n315, A2 => n314, A3 => n313, A4 => n312, Z 
                           => N2036);
   U1276 : AOI22D1 port map( A1 => in_buf_70_port, A2 => n266, B1 => 
                           in_buf_6_port, B2 => n242, Z => n319);
   U1277 : AOI22D1 port map( A1 => in_buf_198_port, A2 => n527, B1 => 
                           in_buf_134_port, B2 => n513, Z => n318);
   U1278 : AOI22D1 port map( A1 => in_buf_102_port, A2 => n529, B1 => 
                           in_buf_38_port, B2 => n515, Z => n317);
   U1279 : AOI22D1 port map( A1 => in_buf_230_port, A2 => n518, B1 => 
                           in_buf_166_port, B2 => n517, Z => n316);
   U1280 : NAN4D1 port map( A1 => n319, A2 => n318, A3 => n317, A4 => n316, Z 
                           => N2035);
   U1281 : AOI22D1 port map( A1 => in_buf_71_port, A2 => n266, B1 => 
                           in_buf_7_port, B2 => n242, Z => n323);
   U1282 : AOI22D1 port map( A1 => in_buf_199_port, A2 => n527, B1 => 
                           in_buf_135_port, B2 => n513, Z => n322);
   U1283 : AOI22D1 port map( A1 => in_buf_103_port, A2 => n529, B1 => 
                           in_buf_39_port, B2 => n515, Z => n321);
   U1284 : AOI22D1 port map( A1 => in_buf_231_port, A2 => n518, B1 => 
                           in_buf_167_port, B2 => n517, Z => n320);
   U1285 : NAN4D1 port map( A1 => n323, A2 => n322, A3 => n321, A4 => n320, Z 
                           => N2034);
   U1286 : AOI22D1 port map( A1 => in_buf_72_port, A2 => n266, B1 => 
                           in_buf_8_port, B2 => n242, Z => n327);
   U1287 : AOI22D1 port map( A1 => in_buf_200_port, A2 => n527, B1 => 
                           in_buf_136_port, B2 => n513, Z => n326);
   U1288 : AOI22D1 port map( A1 => in_buf_104_port, A2 => n516, B1 => 
                           in_buf_40_port, B2 => n515, Z => n325);
   U1289 : AOI22D1 port map( A1 => in_buf_232_port, A2 => n518, B1 => 
                           in_buf_168_port, B2 => n517, Z => n324);
   U1290 : NAN4D1 port map( A1 => n327, A2 => n326, A3 => n325, A4 => n324, Z 
                           => N2033);
   U1291 : AOI22D1 port map( A1 => in_buf_73_port, A2 => n266, B1 => 
                           in_buf_9_port, B2 => n242, Z => n331);
   U1292 : AOI22D1 port map( A1 => in_buf_201_port, A2 => n527, B1 => 
                           in_buf_137_port, B2 => n513, Z => n330);
   U1293 : AOI22D1 port map( A1 => in_buf_105_port, A2 => n516, B1 => 
                           in_buf_41_port, B2 => n515, Z => n329);
   U1294 : AOI22D1 port map( A1 => in_buf_233_port, A2 => n518, B1 => 
                           in_buf_169_port, B2 => n517, Z => n328);
   U1295 : NAN4D1 port map( A1 => n331, A2 => n330, A3 => n329, A4 => n328, Z 
                           => N2032);
   U1296 : AOI22D1 port map( A1 => in_buf_74_port, A2 => n266, B1 => 
                           in_buf_10_port, B2 => n242, Z => n335);
   U1297 : AOI22D1 port map( A1 => in_buf_202_port, A2 => n527, B1 => 
                           in_buf_138_port, B2 => n513, Z => n334);
   U1298 : AOI22D1 port map( A1 => in_buf_106_port, A2 => n516, B1 => 
                           in_buf_42_port, B2 => n515, Z => n333);
   U1299 : AOI22D1 port map( A1 => in_buf_234_port, A2 => n534, B1 => 
                           in_buf_170_port, B2 => n517, Z => n332);
   U1300 : NAN4D1 port map( A1 => n335, A2 => n334, A3 => n333, A4 => n332, Z 
                           => N2031);
   U1301 : AOI22D1 port map( A1 => in_buf_75_port, A2 => n266, B1 => 
                           in_buf_11_port, B2 => n242, Z => n339);
   U1302 : AOI22D1 port map( A1 => in_buf_203_port, A2 => n527, B1 => 
                           in_buf_139_port, B2 => n513, Z => n338);
   U1303 : AOI22D1 port map( A1 => in_buf_107_port, A2 => n516, B1 => 
                           in_buf_43_port, B2 => n515, Z => n337);
   U1304 : AOI22D1 port map( A1 => in_buf_235_port, A2 => n518, B1 => 
                           in_buf_171_port, B2 => n517, Z => n336);
   U1305 : NAN4D1 port map( A1 => n339, A2 => n338, A3 => n337, A4 => n336, Z 
                           => N2030);
   U1306 : AOI22D1 port map( A1 => in_buf_76_port, A2 => n266, B1 => 
                           in_buf_12_port, B2 => n242, Z => n343);
   U1307 : AOI22D1 port map( A1 => in_buf_204_port, A2 => n527, B1 => 
                           in_buf_140_port, B2 => n513, Z => n342);
   U1308 : AOI22D1 port map( A1 => in_buf_108_port, A2 => n529, B1 => 
                           in_buf_44_port, B2 => n515, Z => n341);
   U1309 : AOI22D1 port map( A1 => in_buf_236_port, A2 => n534, B1 => 
                           in_buf_172_port, B2 => n532, Z => n340);
   U1310 : NAN4D1 port map( A1 => n343, A2 => n342, A3 => n341, A4 => n340, Z 
                           => N2029);
   U1311 : AOI22D1 port map( A1 => in_buf_77_port, A2 => n266, B1 => 
                           in_buf_13_port, B2 => n242, Z => n347);
   U1312 : AOI22D1 port map( A1 => in_buf_205_port, A2 => n514, B1 => 
                           in_buf_141_port, B2 => n525, Z => n346);
   U1313 : AOI22D1 port map( A1 => in_buf_109_port, A2 => n516, B1 => 
                           in_buf_45_port, B2 => n515, Z => n345);
   U1314 : AOI22D1 port map( A1 => in_buf_237_port, A2 => n534, B1 => 
                           in_buf_173_port, B2 => n531, Z => n344);
   U1315 : NAN4D1 port map( A1 => n347, A2 => n346, A3 => n345, A4 => n344, Z 
                           => N2028);
   U1316 : AOI22D1 port map( A1 => in_buf_78_port, A2 => n266, B1 => 
                           in_buf_14_port, B2 => n242, Z => n351);
   U1317 : AOI22D1 port map( A1 => in_buf_206_port, A2 => n514, B1 => 
                           in_buf_142_port, B2 => n525, Z => n350);
   U1318 : AOI22D1 port map( A1 => in_buf_110_port, A2 => n516, B1 => 
                           in_buf_46_port, B2 => n515, Z => n349);
   U1319 : AOI22D1 port map( A1 => in_buf_238_port, A2 => n534, B1 => 
                           in_buf_174_port, B2 => n517, Z => n348);
   U1320 : NAN4D1 port map( A1 => n351, A2 => n350, A3 => n349, A4 => n348, Z 
                           => N2027);
   U1321 : AOI22D1 port map( A1 => in_buf_79_port, A2 => n266, B1 => 
                           in_buf_15_port, B2 => n242, Z => n355);
   U1322 : AOI22D1 port map( A1 => in_buf_207_port, A2 => n514, B1 => 
                           in_buf_143_port, B2 => n525, Z => n354);
   U1323 : AOI22D1 port map( A1 => in_buf_111_port, A2 => n516, B1 => 
                           in_buf_47_port, B2 => n515, Z => n353);
   U1324 : AOI22D1 port map( A1 => in_buf_239_port, A2 => n534, B1 => 
                           in_buf_175_port, B2 => n517, Z => n352);
   U1325 : NAN4D1 port map( A1 => n355, A2 => n354, A3 => n353, A4 => n352, Z 
                           => N2026);
   U1326 : AOI22D1 port map( A1 => in_buf_80_port, A2 => n266, B1 => 
                           in_buf_16_port, B2 => n242, Z => n359);
   U1327 : AOI22D1 port map( A1 => in_buf_208_port, A2 => n514, B1 => 
                           in_buf_144_port, B2 => n525, Z => n358);
   U1328 : AOI22D1 port map( A1 => in_buf_112_port, A2 => n516, B1 => 
                           in_buf_48_port, B2 => n515, Z => n357);
   U1329 : AOI22D1 port map( A1 => in_buf_240_port, A2 => n534, B1 => 
                           in_buf_176_port, B2 => n517, Z => n356);
   U1330 : NAN4D1 port map( A1 => n359, A2 => n358, A3 => n357, A4 => n356, Z 
                           => N2025);
   U1331 : AOI22D1 port map( A1 => in_buf_81_port, A2 => n266, B1 => 
                           in_buf_17_port, B2 => n242, Z => n363);
   U1332 : AOI22D1 port map( A1 => in_buf_209_port, A2 => n514, B1 => 
                           in_buf_145_port, B2 => n525, Z => n362);
   U1333 : AOI22D1 port map( A1 => in_buf_113_port, A2 => n516, B1 => 
                           in_buf_49_port, B2 => n515, Z => n361);
   U1334 : AOI22D1 port map( A1 => in_buf_241_port, A2 => n534, B1 => 
                           in_buf_177_port, B2 => n517, Z => n360);
   U1335 : NAN4D1 port map( A1 => n363, A2 => n362, A3 => n361, A4 => n360, Z 
                           => N2024);
   U1336 : AOI22D1 port map( A1 => in_buf_82_port, A2 => n266, B1 => 
                           in_buf_18_port, B2 => n242, Z => n367);
   U1337 : AOI22D1 port map( A1 => in_buf_210_port, A2 => n514, B1 => 
                           in_buf_146_port, B2 => n525, Z => n366);
   U1338 : AOI22D1 port map( A1 => in_buf_114_port, A2 => n516, B1 => 
                           in_buf_50_port, B2 => n515, Z => n365);
   U1339 : AOI22D1 port map( A1 => in_buf_242_port, A2 => n534, B1 => 
                           in_buf_178_port, B2 => n517, Z => n364);
   U1340 : NAN4D1 port map( A1 => n367, A2 => n366, A3 => n365, A4 => n364, Z 
                           => N2023);
   U1341 : AOI22D1 port map( A1 => in_buf_83_port, A2 => n266, B1 => 
                           in_buf_19_port, B2 => n242, Z => n371);
   U1342 : AOI22D1 port map( A1 => in_buf_211_port, A2 => n514, B1 => 
                           in_buf_147_port, B2 => n525, Z => n370);
   U1343 : AOI22D1 port map( A1 => in_buf_115_port, A2 => n516, B1 => 
                           in_buf_51_port, B2 => n515, Z => n369);
   U1344 : AOI22D1 port map( A1 => in_buf_243_port, A2 => n534, B1 => 
                           in_buf_179_port, B2 => n517, Z => n368);
   U1345 : NAN4D1 port map( A1 => n371, A2 => n370, A3 => n369, A4 => n368, Z 
                           => N2022);
   U1346 : AOI22D1 port map( A1 => in_buf_84_port, A2 => n266, B1 => 
                           in_buf_20_port, B2 => n242, Z => n375);
   U1347 : AOI22D1 port map( A1 => in_buf_212_port, A2 => n514, B1 => 
                           in_buf_148_port, B2 => n525, Z => n374);
   U1348 : AOI22D1 port map( A1 => in_buf_116_port, A2 => n516, B1 => 
                           in_buf_52_port, B2 => n515, Z => n373);
   U1349 : AOI22D1 port map( A1 => in_buf_244_port, A2 => n534, B1 => 
                           in_buf_180_port, B2 => n517, Z => n372);
   U1350 : NAN4D1 port map( A1 => n375, A2 => n374, A3 => n373, A4 => n372, Z 
                           => N2021);
   U1351 : AOI22D1 port map( A1 => in_buf_85_port, A2 => n266, B1 => 
                           in_buf_21_port, B2 => n242, Z => n379);
   U1352 : AOI22D1 port map( A1 => in_buf_213_port, A2 => n514, B1 => 
                           in_buf_149_port, B2 => n525, Z => n378);
   U1353 : AOI22D1 port map( A1 => in_buf_117_port, A2 => n516, B1 => 
                           in_buf_53_port, B2 => n515, Z => n377);
   U1354 : AOI22D1 port map( A1 => in_buf_245_port, A2 => n534, B1 => 
                           in_buf_181_port, B2 => n517, Z => n376);
   U1355 : NAN4D1 port map( A1 => n379, A2 => n378, A3 => n377, A4 => n376, Z 
                           => N2020);
   U1356 : AOI22D1 port map( A1 => in_buf_86_port, A2 => n266, B1 => 
                           in_buf_22_port, B2 => n242, Z => n383);
   U1357 : AOI22D1 port map( A1 => in_buf_214_port, A2 => n514, B1 => 
                           in_buf_150_port, B2 => n525, Z => n382);
   U1358 : AOI22D1 port map( A1 => in_buf_118_port, A2 => n516, B1 => 
                           in_buf_54_port, B2 => n515, Z => n381);
   U1359 : AOI22D1 port map( A1 => in_buf_246_port, A2 => n534, B1 => 
                           in_buf_182_port, B2 => n517, Z => n380);
   U1360 : NAN4D1 port map( A1 => n383, A2 => n382, A3 => n381, A4 => n380, Z 
                           => N2019);
   U1361 : AOI22D1 port map( A1 => in_buf_87_port, A2 => n266, B1 => 
                           in_buf_23_port, B2 => n242, Z => n387);
   U1362 : AOI22D1 port map( A1 => in_buf_215_port, A2 => n514, B1 => 
                           in_buf_151_port, B2 => n525, Z => n386);
   U1363 : AOI22D1 port map( A1 => in_buf_119_port, A2 => n516, B1 => 
                           in_buf_55_port, B2 => n515, Z => n385);
   U1364 : AOI22D1 port map( A1 => in_buf_247_port, A2 => n534, B1 => 
                           in_buf_183_port, B2 => n517, Z => n384);
   U1365 : NAN4D1 port map( A1 => n387, A2 => n386, A3 => n385, A4 => n384, Z 
                           => N2018);
   U1366 : AOI22D1 port map( A1 => in_buf_88_port, A2 => n266, B1 => 
                           in_buf_24_port, B2 => n242, Z => n391);
   U1367 : AOI22D1 port map( A1 => in_buf_216_port, A2 => n514, B1 => 
                           in_buf_152_port, B2 => n525, Z => n390);
   U1368 : AOI22D1 port map( A1 => in_buf_120_port, A2 => n516, B1 => 
                           in_buf_56_port, B2 => n515, Z => n389);
   U1369 : AOI22D1 port map( A1 => in_buf_248_port, A2 => n534, B1 => 
                           in_buf_184_port, B2 => n517, Z => n388);
   U1370 : NAN4D1 port map( A1 => n391, A2 => n390, A3 => n389, A4 => n388, Z 
                           => N2017);
   U1371 : AOI22D1 port map( A1 => in_buf_89_port, A2 => n266, B1 => 
                           in_buf_25_port, B2 => n242, Z => n395);
   U1372 : AOI22D1 port map( A1 => in_buf_217_port, A2 => n514, B1 => 
                           in_buf_153_port, B2 => n525, Z => n394);
   U1373 : AOI22D1 port map( A1 => in_buf_121_port, A2 => n516, B1 => 
                           in_buf_57_port, B2 => n515, Z => n393);
   U1374 : AOI22D1 port map( A1 => in_buf_249_port, A2 => n534, B1 => 
                           in_buf_185_port, B2 => n531, Z => n392);
   U1375 : NAN4D1 port map( A1 => n395, A2 => n394, A3 => n393, A4 => n392, Z 
                           => N2016);
   U1376 : AOI22D1 port map( A1 => in_buf_90_port, A2 => n266, B1 => 
                           in_buf_26_port, B2 => n242, Z => n399);
   U1377 : AOI22D1 port map( A1 => in_buf_218_port, A2 => n514, B1 => 
                           in_buf_154_port, B2 => n524, Z => n398);
   U1378 : AOI22D1 port map( A1 => in_buf_122_port, A2 => n516, B1 => 
                           in_buf_58_port, B2 => n515, Z => n397);
   U1379 : AOI22D1 port map( A1 => in_buf_250_port, A2 => n518, B1 => 
                           in_buf_186_port, B2 => n532, Z => n396);
   U1380 : NAN4D1 port map( A1 => n399, A2 => n398, A3 => n397, A4 => n396, Z 
                           => N2015);
   U1381 : AOI22D1 port map( A1 => in_buf_91_port, A2 => n266, B1 => 
                           in_buf_27_port, B2 => n242, Z => n403);
   U1382 : AOI22D1 port map( A1 => in_buf_219_port, A2 => n514, B1 => 
                           in_buf_155_port, B2 => n524, Z => n402);
   U1383 : AOI22D1 port map( A1 => in_buf_123_port, A2 => n516, B1 => 
                           in_buf_59_port, B2 => n515, Z => n401);
   U1384 : AOI22D1 port map( A1 => in_buf_251_port, A2 => n518, B1 => 
                           in_buf_187_port, B2 => n532, Z => n400);
   U1385 : NAN4D1 port map( A1 => n403, A2 => n402, A3 => n401, A4 => n400, Z 
                           => N2014);
   U1386 : AOI22D1 port map( A1 => in_buf_92_port, A2 => n266, B1 => 
                           in_buf_28_port, B2 => n242, Z => n407);
   U1387 : AOI22D1 port map( A1 => in_buf_220_port, A2 => n527, B1 => 
                           in_buf_156_port, B2 => n524, Z => n406);
   U1388 : AOI22D1 port map( A1 => in_buf_124_port, A2 => n516, B1 => 
                           in_buf_60_port, B2 => n515, Z => n405);
   U1389 : AOI22D1 port map( A1 => in_buf_252_port, A2 => n518, B1 => 
                           in_buf_188_port, B2 => n532, Z => n404);
   U1390 : NAN4D1 port map( A1 => n407, A2 => n406, A3 => n405, A4 => n404, Z 
                           => N2013);
   U1391 : AOI22D1 port map( A1 => in_buf_93_port, A2 => n266, B1 => 
                           in_buf_29_port, B2 => n242, Z => n411);
   U1392 : AOI22D1 port map( A1 => in_buf_221_port, A2 => n514, B1 => 
                           in_buf_157_port, B2 => n524, Z => n410);
   U1393 : AOI22D1 port map( A1 => in_buf_125_port, A2 => n516, B1 => 
                           in_buf_61_port, B2 => n515, Z => n409);
   U1394 : AOI22D1 port map( A1 => in_buf_253_port, A2 => n518, B1 => 
                           in_buf_189_port, B2 => n532, Z => n408);
   U1395 : NAN4D1 port map( A1 => n411, A2 => n410, A3 => n409, A4 => n408, Z 
                           => N2012);
   U1396 : AOI22D1 port map( A1 => in_buf_94_port, A2 => n266, B1 => 
                           in_buf_30_port, B2 => n242, Z => n415);
   U1397 : AOI22D1 port map( A1 => in_buf_222_port, A2 => n527, B1 => 
                           in_buf_158_port, B2 => n524, Z => n414);
   U1398 : AOI22D1 port map( A1 => in_buf_126_port, A2 => n516, B1 => 
                           in_buf_62_port, B2 => n515, Z => n413);
   U1399 : AOI22D1 port map( A1 => in_buf_254_port, A2 => n534, B1 => 
                           in_buf_190_port, B2 => n532, Z => n412);
   U1400 : NAN4D1 port map( A1 => n415, A2 => n414, A3 => n413, A4 => n412, Z 
                           => N2011);
   U1401 : AOI22D1 port map( A1 => in_buf_95_port, A2 => n266, B1 => 
                           in_buf_31_port, B2 => n242, Z => n419);
   U1402 : AOI22D1 port map( A1 => in_buf_223_port, A2 => n514, B1 => 
                           in_buf_159_port, B2 => n524, Z => n418);
   U1403 : AOI22D1 port map( A1 => in_buf_255_port, A2 => n518, B1 => 
                           in_buf_191_port, B2 => n532, Z => n416);
   U1404 : NAN4D1 port map( A1 => n419, A2 => n418, A3 => n417, A4 => n416, Z 
                           => N2010);
   U1405 : AOI22D1 port map( A1 => comp_res_96_port, A2 => n514, B1 => 
                           comp_res_32_port, B2 => n524, Z => n422);
   U1406 : AOI22D1 port map( A1 => comp_res_128_port, A2 => n518, B1 => 
                           comp_res_64_port, B2 => n532, Z => n420);
   U1407 : AOI22D1 port map( A1 => comp_res_97_port, A2 => n514, B1 => 
                           comp_res_33_port, B2 => n524, Z => n425);
   U1408 : AOI22D1 port map( A1 => comp_res_129_port, A2 => n518, B1 => 
                           comp_res_65_port, B2 => n532, Z => n423);
   U1409 : AOI22D1 port map( A1 => comp_res_98_port, A2 => n514, B1 => 
                           comp_res_34_port, B2 => n524, Z => n428);
   U1410 : AOI22D1 port map( A1 => comp_res_130_port, A2 => n518, B1 => 
                           comp_res_66_port, B2 => n532, Z => n426);
   U1411 : AOI22D1 port map( A1 => comp_res_99_port, A2 => n514, B1 => 
                           comp_res_35_port, B2 => n524, Z => n431);
   U1412 : AOI22D1 port map( A1 => comp_res_131_port, A2 => n518, B1 => 
                           comp_res_67_port, B2 => n532, Z => n429);
   U1413 : AOI22D1 port map( A1 => comp_res_100_port, A2 => n514, B1 => 
                           comp_res_36_port, B2 => n524, Z => n434);
   U1414 : AOI22D1 port map( A1 => comp_res_132_port, A2 => n518, B1 => 
                           comp_res_68_port, B2 => n532, Z => n432);
   U1415 : AOI22D1 port map( A1 => comp_res_101_port, A2 => n514, B1 => 
                           comp_res_37_port, B2 => n524, Z => n437);
   U1416 : AOI22D1 port map( A1 => comp_res_133_port, A2 => n518, B1 => 
                           comp_res_69_port, B2 => n532, Z => n435);
   U1417 : AOI22D1 port map( A1 => comp_res_102_port, A2 => n514, B1 => 
                           comp_res_38_port, B2 => n524, Z => n440);
   U1418 : AOI22D1 port map( A1 => comp_res_134_port, A2 => n518, B1 => 
                           comp_res_70_port, B2 => n532, Z => n438);
   U1419 : AOI22D1 port map( A1 => comp_res_103_port, A2 => n514, B1 => 
                           comp_res_39_port, B2 => n525, Z => n443);
   U1420 : AOI22D1 port map( A1 => comp_res_135_port, A2 => n518, B1 => 
                           comp_res_71_port, B2 => n531, Z => n441);
   U1421 : AOI22D1 port map( A1 => comp_res_104_port, A2 => n514, B1 => 
                           comp_res_40_port, B2 => n513, Z => n446);
   U1422 : AOI22D1 port map( A1 => comp_res_136_port, A2 => n534, B1 => 
                           comp_res_72_port, B2 => n517, Z => n444);
   U1423 : AOI22D1 port map( A1 => comp_res_105_port, A2 => n514, B1 => 
                           comp_res_41_port, B2 => n525, Z => n449);
   U1424 : AOI22D1 port map( A1 => comp_res_137_port, A2 => n518, B1 => 
                           comp_res_73_port, B2 => n517, Z => n447);
   U1425 : AOI22D1 port map( A1 => comp_res_106_port, A2 => n514, B1 => 
                           comp_res_42_port, B2 => n524, Z => n452);
   U1426 : AOI22D1 port map( A1 => comp_res_138_port, A2 => n534, B1 => 
                           comp_res_74_port, B2 => n517, Z => n450);
   U1427 : AOI22D1 port map( A1 => comp_res_107_port, A2 => n527, B1 => 
                           comp_res_43_port, B2 => n513, Z => n455);
   U1428 : AOI22D1 port map( A1 => comp_res_139_port, A2 => n518, B1 => 
                           comp_res_75_port, B2 => n532, Z => n453);
   U1429 : AOI22D1 port map( A1 => comp_res_108_port, A2 => n514, B1 => 
                           comp_res_44_port, B2 => n525, Z => n458);
   U1430 : AOI22D1 port map( A1 => comp_res_140_port, A2 => n534, B1 => 
                           comp_res_76_port, B2 => n517, Z => n456);
   U1431 : AOI22D1 port map( A1 => comp_res_109_port, A2 => n514, B1 => 
                           comp_res_45_port, B2 => n524, Z => n461);
   U1432 : AOI22D1 port map( A1 => comp_res_141_port, A2 => n518, B1 => 
                           comp_res_77_port, B2 => n517, Z => n459);
   U1433 : AOI22D1 port map( A1 => comp_res_110_port, A2 => n514, B1 => 
                           comp_res_46_port, B2 => n513, Z => n464);
   U1434 : AOI22D1 port map( A1 => comp_res_142_port, A2 => n534, B1 => 
                           comp_res_78_port, B2 => n532, Z => n462);
   U1435 : AOI22D1 port map( A1 => comp_res_111_port, A2 => n514, B1 => 
                           comp_res_47_port, B2 => n524, Z => n467);
   U1436 : AOI22D1 port map( A1 => comp_res_143_port, A2 => n518, B1 => 
                           comp_res_79_port, B2 => n531, Z => n465);
   U1437 : AOI22D1 port map( A1 => comp_res_112_port, A2 => n514, B1 => 
                           comp_res_48_port, B2 => n513, Z => n470);
   U1438 : AOI22D1 port map( A1 => comp_res_144_port, A2 => n518, B1 => 
                           comp_res_80_port, B2 => n517, Z => n468);
   U1439 : AOI22D1 port map( A1 => comp_res_113_port, A2 => n514, B1 => 
                           comp_res_49_port, B2 => n513, Z => n473);
   U1440 : AOI22D1 port map( A1 => comp_res_145_port, A2 => n518, B1 => 
                           comp_res_81_port, B2 => n531, Z => n471);
   U1441 : AOI22D1 port map( A1 => comp_res_114_port, A2 => n514, B1 => 
                           comp_res_50_port, B2 => n524, Z => n476);
   U1442 : AOI22D1 port map( A1 => comp_res_146_port, A2 => n534, B1 => 
                           comp_res_82_port, B2 => n531, Z => n474);
   U1443 : AOI22D1 port map( A1 => comp_res_115_port, A2 => n514, B1 => 
                           comp_res_51_port, B2 => n524, Z => n479);
   U1444 : AOI22D1 port map( A1 => comp_res_147_port, A2 => n518, B1 => 
                           comp_res_83_port, B2 => n531, Z => n477);
   U1445 : AOI22D1 port map( A1 => comp_res_116_port, A2 => n514, B1 => 
                           comp_res_52_port, B2 => n513, Z => n482);
   U1446 : AOI22D1 port map( A1 => comp_res_148_port, A2 => n518, B1 => 
                           comp_res_84_port, B2 => n531, Z => n480);
   U1447 : AOI22D1 port map( A1 => comp_res_117_port, A2 => n514, B1 => 
                           comp_res_53_port, B2 => n513, Z => n485);
   U1448 : AOI22D1 port map( A1 => comp_res_149_port, A2 => n518, B1 => 
                           comp_res_85_port, B2 => n531, Z => n483);
   U1449 : AOI22D1 port map( A1 => comp_res_118_port, A2 => n514, B1 => 
                           comp_res_54_port, B2 => n513, Z => n488);
   U1450 : AOI22D1 port map( A1 => comp_res_150_port, A2 => n518, B1 => 
                           comp_res_86_port, B2 => n531, Z => n486);
   U1451 : AOI22D1 port map( A1 => comp_res_119_port, A2 => n527, B1 => 
                           comp_res_55_port, B2 => n513, Z => n491);
   U1452 : AOI22D1 port map( A1 => comp_res_151_port, A2 => n518, B1 => 
                           comp_res_87_port, B2 => n531, Z => n489);
   U1453 : AOI22D1 port map( A1 => comp_res_120_port, A2 => n514, B1 => 
                           comp_res_56_port, B2 => n513, Z => n494);
   U1454 : AOI22D1 port map( A1 => comp_res_152_port, A2 => n518, B1 => 
                           comp_res_88_port, B2 => n531, Z => n492);
   U1455 : AOI22D1 port map( A1 => comp_res_121_port, A2 => n514, B1 => 
                           comp_res_57_port, B2 => n513, Z => n497);
   U1456 : AOI22D1 port map( A1 => comp_res_153_port, A2 => n534, B1 => 
                           comp_res_89_port, B2 => n531, Z => n495);
   U1457 : AOI22D1 port map( A1 => comp_res_122_port, A2 => n514, B1 => 
                           comp_res_58_port, B2 => n513, Z => n500);
   U1458 : AOI22D1 port map( A1 => comp_res_154_port, A2 => n518, B1 => 
                           comp_res_90_port, B2 => n531, Z => n498);
   U1459 : AOI22D1 port map( A1 => comp_res_123_port, A2 => n514, B1 => 
                           comp_res_59_port, B2 => n513, Z => n503);
   U1460 : AOI22D1 port map( A1 => comp_res_155_port, A2 => n518, B1 => 
                           comp_res_91_port, B2 => n531, Z => n501);
   U1461 : AOI22D1 port map( A1 => comp_res_124_port, A2 => n514, B1 => 
                           comp_res_60_port, B2 => n513, Z => n506);
   U1462 : AOI22D1 port map( A1 => comp_res_156_port, A2 => n534, B1 => 
                           comp_res_92_port, B2 => n531, Z => n504);
   U1463 : AOI22D1 port map( A1 => comp_res_125_port, A2 => n514, B1 => 
                           comp_res_61_port, B2 => n513, Z => n509);
   U1464 : AOI22D1 port map( A1 => comp_res_157_port, A2 => n518, B1 => 
                           comp_res_93_port, B2 => n531, Z => n507);
   U1465 : AOI22D1 port map( A1 => comp_res_126_port, A2 => n514, B1 => 
                           comp_res_62_port, B2 => n513, Z => n512);
   U1466 : AOI22D1 port map( A1 => comp_res_158_port, A2 => n534, B1 => 
                           comp_res_94_port, B2 => n531, Z => n510);
   U1467 : AOI22D1 port map( A1 => comp_res_127_port, A2 => n514, B1 => 
                           comp_res_63_port, B2 => n525, Z => n521);
   U1468 : AOI22D1 port map( A1 => comp_res_159_port, A2 => n518, B1 => 
                           comp_res_95_port, B2 => n531, Z => n519);
   U1469 : NOR2D1 port map( A1 => n671, A2 => N63, Z => n535);
   U1470 : NOR2D1 port map( A1 => n671, A2 => n697, Z => n536);
   U1471 : AOI22D1 port map( A1 => out_buf_80_port, A2 => n268, B1 => 
                           out_buf_16_port, B2 => n243, Z => n542);
   U1472 : NOR2D1 port map( A1 => N63, A2 => N64, Z => n537);
   U1473 : NOR2D1 port map( A1 => n697, A2 => N64, Z => n538);
   U1474 : AOI22D1 port map( A1 => out_buf_208_port, A2 => n269, B1 => 
                           out_buf_144_port, B2 => n244, Z => n541);
   U1475 : NOR2M1D1 port map( A1 => n535, A2 => N62, Z => n664);
   U1476 : NOR2M1D1 port map( A1 => n536, A2 => N62, Z => n663);
   U1477 : AOI22D1 port map( A1 => out_buf_112_port, A2 => n664, B1 => 
                           out_buf_48_port, B2 => n663, Z => n540);
   U1478 : NOR2M1D1 port map( A1 => n537, A2 => N62, Z => n666);
   U1479 : NOR2M1D1 port map( A1 => n538, A2 => N62, Z => n665);
   U1480 : AOI22D1 port map( A1 => out_buf_240_port, A2 => n666, B1 => 
                           out_buf_176_port, B2 => n665, Z => n539);
   U1481 : NAN4D1 port map( A1 => n542, A2 => n541, A3 => n540, A4 => n539, Z 
                           => N2882);
   U1482 : AOI22D1 port map( A1 => out_buf_81_port, A2 => n268, B1 => 
                           out_buf_17_port, B2 => n243, Z => n546);
   U1483 : AOI22D1 port map( A1 => out_buf_209_port, A2 => n269, B1 => 
                           out_buf_145_port, B2 => n244, Z => n545);
   U1484 : AOI22D1 port map( A1 => out_buf_113_port, A2 => n664, B1 => 
                           out_buf_49_port, B2 => n663, Z => n544);
   U1485 : AOI22D1 port map( A1 => out_buf_241_port, A2 => n666, B1 => 
                           out_buf_177_port, B2 => n665, Z => n543);
   U1486 : NAN4D1 port map( A1 => n546, A2 => n545, A3 => n544, A4 => n543, Z 
                           => N2881);
   U1487 : AOI22D1 port map( A1 => out_buf_82_port, A2 => n268, B1 => 
                           out_buf_18_port, B2 => n243, Z => n550);
   U1488 : AOI22D1 port map( A1 => out_buf_210_port, A2 => n269, B1 => 
                           out_buf_146_port, B2 => n244, Z => n549);
   U1489 : AOI22D1 port map( A1 => out_buf_114_port, A2 => n664, B1 => 
                           out_buf_50_port, B2 => n663, Z => n548);
   U1490 : AOI22D1 port map( A1 => out_buf_242_port, A2 => n666, B1 => 
                           out_buf_178_port, B2 => n665, Z => n547);
   U1491 : NAN4D1 port map( A1 => n550, A2 => n549, A3 => n548, A4 => n547, Z 
                           => N2880);
   U1492 : AOI22D1 port map( A1 => out_buf_83_port, A2 => n268, B1 => 
                           out_buf_19_port, B2 => n243, Z => n554);
   U1493 : AOI22D1 port map( A1 => out_buf_211_port, A2 => n269, B1 => 
                           out_buf_147_port, B2 => n244, Z => n553);
   U1494 : AOI22D1 port map( A1 => out_buf_115_port, A2 => n664, B1 => 
                           out_buf_51_port, B2 => n663, Z => n552);
   U1495 : AOI22D1 port map( A1 => out_buf_243_port, A2 => n666, B1 => 
                           out_buf_179_port, B2 => n665, Z => n551);
   U1496 : NAN4D1 port map( A1 => n554, A2 => n553, A3 => n552, A4 => n551, Z 
                           => N2879);
   U1497 : AOI22D1 port map( A1 => out_buf_84_port, A2 => n268, B1 => 
                           out_buf_20_port, B2 => n243, Z => n558);
   U1498 : AOI22D1 port map( A1 => out_buf_212_port, A2 => n269, B1 => 
                           out_buf_148_port, B2 => n244, Z => n557);
   U1499 : AOI22D1 port map( A1 => out_buf_116_port, A2 => n664, B1 => 
                           out_buf_52_port, B2 => n663, Z => n556);
   U1500 : AOI22D1 port map( A1 => out_buf_244_port, A2 => n666, B1 => 
                           out_buf_180_port, B2 => n665, Z => n555);
   U1501 : NAN4D1 port map( A1 => n558, A2 => n557, A3 => n556, A4 => n555, Z 
                           => N2878);
   U1502 : AOI22D1 port map( A1 => out_buf_85_port, A2 => n268, B1 => 
                           out_buf_21_port, B2 => n243, Z => n562);
   U1503 : AOI22D1 port map( A1 => out_buf_213_port, A2 => n269, B1 => 
                           out_buf_149_port, B2 => n244, Z => n561);
   U1504 : AOI22D1 port map( A1 => out_buf_117_port, A2 => n664, B1 => 
                           out_buf_53_port, B2 => n663, Z => n560);
   U1505 : AOI22D1 port map( A1 => out_buf_245_port, A2 => n666, B1 => 
                           out_buf_181_port, B2 => n665, Z => n559);
   U1506 : NAN4D1 port map( A1 => n562, A2 => n561, A3 => n560, A4 => n559, Z 
                           => N2877);
   U1507 : AOI22D1 port map( A1 => out_buf_86_port, A2 => n268, B1 => 
                           out_buf_22_port, B2 => n243, Z => n566);
   U1508 : AOI22D1 port map( A1 => out_buf_214_port, A2 => n269, B1 => 
                           out_buf_150_port, B2 => n244, Z => n565);
   U1509 : AOI22D1 port map( A1 => out_buf_118_port, A2 => n664, B1 => 
                           out_buf_54_port, B2 => n663, Z => n564);
   U1510 : AOI22D1 port map( A1 => out_buf_246_port, A2 => n666, B1 => 
                           out_buf_182_port, B2 => n665, Z => n563);
   U1511 : NAN4D1 port map( A1 => n566, A2 => n565, A3 => n564, A4 => n563, Z 
                           => N2876);
   U1512 : AOI22D1 port map( A1 => out_buf_87_port, A2 => n268, B1 => 
                           out_buf_23_port, B2 => n243, Z => n570);
   U1513 : AOI22D1 port map( A1 => out_buf_215_port, A2 => n269, B1 => 
                           out_buf_151_port, B2 => n244, Z => n569);
   U1514 : AOI22D1 port map( A1 => out_buf_119_port, A2 => n664, B1 => 
                           out_buf_55_port, B2 => n663, Z => n568);
   U1515 : AOI22D1 port map( A1 => out_buf_247_port, A2 => n666, B1 => 
                           out_buf_183_port, B2 => n665, Z => n567);
   U1516 : NAN4D1 port map( A1 => n570, A2 => n569, A3 => n568, A4 => n567, Z 
                           => N2875);
   U1517 : AOI22D1 port map( A1 => out_buf_88_port, A2 => n268, B1 => 
                           out_buf_24_port, B2 => n243, Z => n574);
   U1518 : AOI22D1 port map( A1 => out_buf_216_port, A2 => n269, B1 => 
                           out_buf_152_port, B2 => n244, Z => n573);
   U1519 : AOI22D1 port map( A1 => out_buf_120_port, A2 => n664, B1 => 
                           out_buf_56_port, B2 => n663, Z => n572);
   U1520 : AOI22D1 port map( A1 => out_buf_248_port, A2 => n666, B1 => 
                           out_buf_184_port, B2 => n665, Z => n571);
   U1521 : NAN4D1 port map( A1 => n574, A2 => n573, A3 => n572, A4 => n571, Z 
                           => N2874);
   U1522 : AOI22D1 port map( A1 => out_buf_89_port, A2 => n268, B1 => 
                           out_buf_25_port, B2 => n243, Z => n578);
   U1523 : AOI22D1 port map( A1 => out_buf_217_port, A2 => n269, B1 => 
                           out_buf_153_port, B2 => n244, Z => n577);
   U1524 : AOI22D1 port map( A1 => out_buf_121_port, A2 => n664, B1 => 
                           out_buf_57_port, B2 => n663, Z => n576);
   U1525 : AOI22D1 port map( A1 => out_buf_249_port, A2 => n666, B1 => 
                           out_buf_185_port, B2 => n665, Z => n575);
   U1526 : NAN4D1 port map( A1 => n578, A2 => n577, A3 => n576, A4 => n575, Z 
                           => N2873);
   U1527 : AOI22D1 port map( A1 => out_buf_90_port, A2 => n268, B1 => 
                           out_buf_26_port, B2 => n243, Z => n582);
   U1528 : AOI22D1 port map( A1 => out_buf_218_port, A2 => n269, B1 => 
                           out_buf_154_port, B2 => n244, Z => n581);
   U1529 : AOI22D1 port map( A1 => out_buf_122_port, A2 => n664, B1 => 
                           out_buf_58_port, B2 => n663, Z => n580);
   U1530 : AOI22D1 port map( A1 => out_buf_250_port, A2 => n666, B1 => 
                           out_buf_186_port, B2 => n665, Z => n579);
   U1531 : NAN4D1 port map( A1 => n582, A2 => n581, A3 => n580, A4 => n579, Z 
                           => N2872);
   U1532 : AOI22D1 port map( A1 => out_buf_91_port, A2 => n268, B1 => 
                           out_buf_27_port, B2 => n243, Z => n586);
   U1533 : AOI22D1 port map( A1 => out_buf_219_port, A2 => n269, B1 => 
                           out_buf_155_port, B2 => n244, Z => n585);
   U1534 : AOI22D1 port map( A1 => out_buf_123_port, A2 => n664, B1 => 
                           out_buf_59_port, B2 => n663, Z => n584);
   U1535 : AOI22D1 port map( A1 => out_buf_251_port, A2 => n666, B1 => 
                           out_buf_187_port, B2 => n665, Z => n583);
   U1536 : NAN4D1 port map( A1 => n586, A2 => n585, A3 => n584, A4 => n583, Z 
                           => N2871);
   U1537 : AOI22D1 port map( A1 => out_buf_92_port, A2 => n268, B1 => 
                           out_buf_28_port, B2 => n243, Z => n5901);
   U1538 : AOI22D1 port map( A1 => out_buf_220_port, A2 => n269, B1 => 
                           out_buf_156_port, B2 => n244, Z => n589);
   U1539 : AOI22D1 port map( A1 => out_buf_124_port, A2 => n664, B1 => 
                           out_buf_60_port, B2 => n663, Z => n588);
   U1540 : AOI22D1 port map( A1 => out_buf_252_port, A2 => n666, B1 => 
                           out_buf_188_port, B2 => n665, Z => n587);
   U1541 : NAN4D1 port map( A1 => n5901, A2 => n589, A3 => n588, A4 => n587, Z 
                           => N2870);
   U1542 : AOI22D1 port map( A1 => out_buf_93_port, A2 => n268, B1 => 
                           out_buf_29_port, B2 => n243, Z => n594);
   U1543 : AOI22D1 port map( A1 => out_buf_221_port, A2 => n269, B1 => 
                           out_buf_157_port, B2 => n244, Z => n593);
   U1544 : AOI22D1 port map( A1 => out_buf_125_port, A2 => n664, B1 => 
                           out_buf_61_port, B2 => n663, Z => n592);
   U1545 : AOI22D1 port map( A1 => out_buf_253_port, A2 => n666, B1 => 
                           out_buf_189_port, B2 => n665, Z => n591);
   U1546 : NAN4D1 port map( A1 => n594, A2 => n593, A3 => n592, A4 => n591, Z 
                           => N2869);
   U1547 : AOI22D1 port map( A1 => out_buf_94_port, A2 => n268, B1 => 
                           out_buf_30_port, B2 => n243, Z => n598);
   U1548 : AOI22D1 port map( A1 => out_buf_222_port, A2 => n269, B1 => 
                           out_buf_158_port, B2 => n244, Z => n597);
   U1549 : AOI22D1 port map( A1 => out_buf_126_port, A2 => n664, B1 => 
                           out_buf_62_port, B2 => n663, Z => n596);
   U1550 : AOI22D1 port map( A1 => out_buf_254_port, A2 => n666, B1 => 
                           out_buf_190_port, B2 => n665, Z => n595);
   U1551 : NAN4D1 port map( A1 => n598, A2 => n597, A3 => n596, A4 => n595, Z 
                           => N2868);
   U1552 : AOI22D1 port map( A1 => out_buf_95_port, A2 => n268, B1 => 
                           out_buf_31_port, B2 => n243, Z => n602);
   U1553 : AOI22D1 port map( A1 => out_buf_223_port, A2 => n269, B1 => 
                           out_buf_159_port, B2 => n244, Z => n601);
   U1554 : AOI22D1 port map( A1 => out_buf_127_port, A2 => n664, B1 => 
                           out_buf_63_port, B2 => n663, Z => n6001);
   U1555 : AOI22D1 port map( A1 => out_buf_255_port, A2 => n666, B1 => 
                           out_buf_191_port, B2 => n665, Z => n599);
   U1556 : NAN4D1 port map( A1 => n602, A2 => n601, A3 => n6001, A4 => n599, Z 
                           => N2867);
   U1557 : AOI22D1 port map( A1 => out_buf_64_port, A2 => n268, B1 => 
                           out_buf_0_port, B2 => n243, Z => n606);
   U1558 : AOI22D1 port map( A1 => out_buf_192_port, A2 => n269, B1 => 
                           out_buf_128_port, B2 => n244, Z => n605);
   U1559 : AOI22D1 port map( A1 => out_buf_96_port, A2 => n664, B1 => 
                           out_buf_32_port, B2 => n663, Z => n604);
   U1560 : AOI22D1 port map( A1 => out_buf_224_port, A2 => n666, B1 => 
                           out_buf_160_port, B2 => n665, Z => n603);
   U1561 : NAN4D1 port map( A1 => n606, A2 => n605, A3 => n604, A4 => n603, Z 
                           => N2865);
   U1562 : AOI22D1 port map( A1 => out_buf_65_port, A2 => n268, B1 => 
                           out_buf_1_port, B2 => n243, Z => n6101);
   U1563 : AOI22D1 port map( A1 => out_buf_193_port, A2 => n269, B1 => 
                           out_buf_129_port, B2 => n244, Z => n609);
   U1564 : AOI22D1 port map( A1 => out_buf_97_port, A2 => n664, B1 => 
                           out_buf_33_port, B2 => n663, Z => n608);
   U1565 : AOI22D1 port map( A1 => out_buf_225_port, A2 => n666, B1 => 
                           out_buf_161_port, B2 => n665, Z => n607);
   U1566 : NAN4D1 port map( A1 => n6101, A2 => n609, A3 => n608, A4 => n607, Z 
                           => N2864);
   U1567 : AOI22D1 port map( A1 => out_buf_66_port, A2 => n268, B1 => 
                           out_buf_2_port, B2 => n243, Z => n614);
   U1568 : AOI22D1 port map( A1 => out_buf_194_port, A2 => n269, B1 => 
                           out_buf_130_port, B2 => n244, Z => n613);
   U1569 : AOI22D1 port map( A1 => out_buf_98_port, A2 => n664, B1 => 
                           out_buf_34_port, B2 => n663, Z => n612);
   U1570 : AOI22D1 port map( A1 => out_buf_226_port, A2 => n666, B1 => 
                           out_buf_162_port, B2 => n665, Z => n611);
   U1571 : NAN4D1 port map( A1 => n614, A2 => n613, A3 => n612, A4 => n611, Z 
                           => N2863);
   U1572 : AOI22D1 port map( A1 => out_buf_67_port, A2 => n268, B1 => 
                           out_buf_3_port, B2 => n243, Z => n618);
   U1573 : AOI22D1 port map( A1 => out_buf_195_port, A2 => n269, B1 => 
                           out_buf_131_port, B2 => n244, Z => n617);
   U1574 : AOI22D1 port map( A1 => out_buf_99_port, A2 => n664, B1 => 
                           out_buf_35_port, B2 => n663, Z => n616);
   U1575 : AOI22D1 port map( A1 => out_buf_227_port, A2 => n666, B1 => 
                           out_buf_163_port, B2 => n665, Z => n615);
   U1576 : NAN4D1 port map( A1 => n618, A2 => n617, A3 => n616, A4 => n615, Z 
                           => N2862);
   U1577 : AOI22D1 port map( A1 => out_buf_68_port, A2 => n268, B1 => 
                           out_buf_4_port, B2 => n243, Z => n622);
   U1578 : AOI22D1 port map( A1 => out_buf_196_port, A2 => n269, B1 => 
                           out_buf_132_port, B2 => n244, Z => n621);
   U1579 : AOI22D1 port map( A1 => out_buf_100_port, A2 => n664, B1 => 
                           out_buf_36_port, B2 => n663, Z => n620);
   U1580 : AOI22D1 port map( A1 => out_buf_228_port, A2 => n666, B1 => 
                           out_buf_164_port, B2 => n665, Z => n619);
   U1581 : NAN4D1 port map( A1 => n622, A2 => n621, A3 => n620, A4 => n619, Z 
                           => N2861);
   U1582 : AOI22D1 port map( A1 => out_buf_69_port, A2 => n268, B1 => 
                           out_buf_5_port, B2 => n243, Z => n626);
   U1583 : AOI22D1 port map( A1 => out_buf_197_port, A2 => n269, B1 => 
                           out_buf_133_port, B2 => n244, Z => n625);
   U1584 : AOI22D1 port map( A1 => out_buf_101_port, A2 => n664, B1 => 
                           out_buf_37_port, B2 => n663, Z => n624);
   U1585 : AOI22D1 port map( A1 => out_buf_229_port, A2 => n666, B1 => 
                           out_buf_165_port, B2 => n665, Z => n623);
   U1586 : NAN4D1 port map( A1 => n626, A2 => n625, A3 => n624, A4 => n623, Z 
                           => N2860);
   U1587 : AOI22D1 port map( A1 => out_buf_70_port, A2 => n268, B1 => 
                           out_buf_6_port, B2 => n243, Z => n6301);
   U1588 : AOI22D1 port map( A1 => out_buf_198_port, A2 => n269, B1 => 
                           out_buf_134_port, B2 => n244, Z => n629);
   U1589 : AOI22D1 port map( A1 => out_buf_102_port, A2 => n664, B1 => 
                           out_buf_38_port, B2 => n663, Z => n628);
   U1590 : AOI22D1 port map( A1 => out_buf_230_port, A2 => n666, B1 => 
                           out_buf_166_port, B2 => n665, Z => n627);
   U1591 : NAN4D1 port map( A1 => n6301, A2 => n629, A3 => n628, A4 => n627, Z 
                           => N2859);
   U1592 : AOI22D1 port map( A1 => out_buf_71_port, A2 => n268, B1 => 
                           out_buf_7_port, B2 => n243, Z => n634);
   U1593 : AOI22D1 port map( A1 => out_buf_199_port, A2 => n269, B1 => 
                           out_buf_135_port, B2 => n244, Z => n633);
   U1594 : AOI22D1 port map( A1 => out_buf_103_port, A2 => n664, B1 => 
                           out_buf_39_port, B2 => n663, Z => n632);
   U1595 : AOI22D1 port map( A1 => out_buf_231_port, A2 => n666, B1 => 
                           out_buf_167_port, B2 => n665, Z => n631);
   U1596 : NAN4D1 port map( A1 => n634, A2 => n633, A3 => n632, A4 => n631, Z 
                           => N2858);
   U1597 : AOI22D1 port map( A1 => out_buf_72_port, A2 => n268, B1 => 
                           out_buf_8_port, B2 => n243, Z => n638);
   U1598 : AOI22D1 port map( A1 => out_buf_200_port, A2 => n269, B1 => 
                           out_buf_136_port, B2 => n244, Z => n637);
   U1599 : AOI22D1 port map( A1 => out_buf_104_port, A2 => n664, B1 => 
                           out_buf_40_port, B2 => n663, Z => n636);
   U1600 : AOI22D1 port map( A1 => out_buf_232_port, A2 => n666, B1 => 
                           out_buf_168_port, B2 => n665, Z => n635);
   U1601 : NAN4D1 port map( A1 => n638, A2 => n637, A3 => n636, A4 => n635, Z 
                           => N2857);
   U1602 : AOI22D1 port map( A1 => out_buf_73_port, A2 => n268, B1 => 
                           out_buf_9_port, B2 => n243, Z => n642);
   U1603 : AOI22D1 port map( A1 => out_buf_201_port, A2 => n269, B1 => 
                           out_buf_137_port, B2 => n244, Z => n641);
   U1604 : AOI22D1 port map( A1 => out_buf_105_port, A2 => n664, B1 => 
                           out_buf_41_port, B2 => n663, Z => n6401);
   U1605 : AOI22D1 port map( A1 => out_buf_233_port, A2 => n666, B1 => 
                           out_buf_169_port, B2 => n665, Z => n639);
   U1606 : NAN4D1 port map( A1 => n642, A2 => n641, A3 => n6401, A4 => n639, Z 
                           => N2856);
   U1607 : AOI22D1 port map( A1 => out_buf_74_port, A2 => n268, B1 => 
                           out_buf_10_port, B2 => n243, Z => n646);
   U1608 : AOI22D1 port map( A1 => out_buf_202_port, A2 => n269, B1 => 
                           out_buf_138_port, B2 => n244, Z => n645);
   U1609 : AOI22D1 port map( A1 => out_buf_106_port, A2 => n664, B1 => 
                           out_buf_42_port, B2 => n663, Z => n644);
   U1610 : AOI22D1 port map( A1 => out_buf_234_port, A2 => n666, B1 => 
                           out_buf_170_port, B2 => n665, Z => n643);
   U1611 : NAN4D1 port map( A1 => n646, A2 => n645, A3 => n644, A4 => n643, Z 
                           => N2855);
   U1612 : AOI22D1 port map( A1 => out_buf_75_port, A2 => n268, B1 => 
                           out_buf_11_port, B2 => n243, Z => n650);
   U1613 : AOI22D1 port map( A1 => out_buf_203_port, A2 => n269, B1 => 
                           out_buf_139_port, B2 => n244, Z => n649);
   U1614 : AOI22D1 port map( A1 => out_buf_107_port, A2 => n664, B1 => 
                           out_buf_43_port, B2 => n663, Z => n648);
   U1615 : AOI22D1 port map( A1 => out_buf_235_port, A2 => n666, B1 => 
                           out_buf_171_port, B2 => n665, Z => n647);
   U1616 : NAN4D1 port map( A1 => n650, A2 => n649, A3 => n648, A4 => n647, Z 
                           => N2854);
   U1617 : AOI22D1 port map( A1 => out_buf_76_port, A2 => n268, B1 => 
                           out_buf_12_port, B2 => n243, Z => n654);
   U1618 : AOI22D1 port map( A1 => out_buf_204_port, A2 => n269, B1 => 
                           out_buf_140_port, B2 => n244, Z => n653);
   U1619 : AOI22D1 port map( A1 => out_buf_108_port, A2 => n664, B1 => 
                           out_buf_44_port, B2 => n663, Z => n652);
   U1620 : AOI22D1 port map( A1 => out_buf_236_port, A2 => n666, B1 => 
                           out_buf_172_port, B2 => n665, Z => n651);
   U1621 : NAN4D1 port map( A1 => n654, A2 => n653, A3 => n652, A4 => n651, Z 
                           => N2853);
   U1622 : AOI22D1 port map( A1 => out_buf_77_port, A2 => n268, B1 => 
                           out_buf_13_port, B2 => n243, Z => n658);
   U1623 : AOI22D1 port map( A1 => out_buf_205_port, A2 => n269, B1 => 
                           out_buf_141_port, B2 => n244, Z => n657);
   U1624 : AOI22D1 port map( A1 => out_buf_109_port, A2 => n664, B1 => 
                           out_buf_45_port, B2 => n663, Z => n656);
   U1625 : AOI22D1 port map( A1 => out_buf_237_port, A2 => n666, B1 => 
                           out_buf_173_port, B2 => n665, Z => n655);
   U1626 : NAN4D1 port map( A1 => n658, A2 => n657, A3 => n656, A4 => n655, Z 
                           => N2852);
   U1627 : AOI22D1 port map( A1 => out_buf_78_port, A2 => n268, B1 => 
                           out_buf_14_port, B2 => n243, Z => n662);
   U1628 : AOI22D1 port map( A1 => out_buf_206_port, A2 => n269, B1 => 
                           out_buf_142_port, B2 => n244, Z => n661);
   U1629 : AOI22D1 port map( A1 => out_buf_110_port, A2 => n664, B1 => 
                           out_buf_46_port, B2 => n663, Z => n660);
   U1630 : AOI22D1 port map( A1 => out_buf_238_port, A2 => n666, B1 => 
                           out_buf_174_port, B2 => n665, Z => n659);
   U1631 : NAN4D1 port map( A1 => n662, A2 => n661, A3 => n660, A4 => n659, Z 
                           => N2851);
   U1632 : AOI22D1 port map( A1 => out_buf_79_port, A2 => n268, B1 => 
                           out_buf_15_port, B2 => n243, Z => n670);
   U1633 : AOI22D1 port map( A1 => out_buf_207_port, A2 => n269, B1 => 
                           out_buf_143_port, B2 => n244, Z => n669);
   U1634 : AOI22D1 port map( A1 => out_buf_111_port, A2 => n664, B1 => 
                           out_buf_47_port, B2 => n663, Z => n668);
   U1635 : AOI22D1 port map( A1 => out_buf_239_port, A2 => n666, B1 => 
                           out_buf_175_port, B2 => n665, Z => n667);
   U1636 : NAN4D1 port map( A1 => n670, A2 => n669, A3 => n668, A4 => n667, Z 
                           => N2850);
   U1637 : NOR3D1 port map( A1 => avs_addr(3), A2 => avs_addr(5), A3 => 
                           avs_addr(4), Z => N66);
   mult_21_C241_U1396 : AOI21D1 port map( A1 => N2940, A2 => N2941, B => 
                           mult_21_C241_n1421, Z => mult_21_C241_n940);
   mult_21_C241_U1395 : OAI21D1 port map( A1 => N2943, A2 => N2942, B => 
                           mult_21_C241_n1422, Z => mult_21_C241_n104);
   mult_21_C241_U1394 : AOI21D1 port map( A1 => N2942, A2 => N2943, B => 
                           mult_21_C241_n1422, Z => mult_21_C241_n939);
   mult_21_C241_U1393 : AOI21D1 port map( A1 => N2914, A2 => N2915, B => 
                           mult_21_C241_n1395, Z => mult_21_C241_n953);
   mult_21_C241_U1392 : AOI21D1 port map( A1 => N2916, A2 => N2917, B => 
                           mult_21_C241_n1397, Z => mult_21_C241_n952);
   mult_21_C241_U1391 : AOI21D1 port map( A1 => N2918, A2 => N2919, B => 
                           mult_21_C241_n1399, Z => mult_21_C241_n951);
   mult_21_C241_U1390 : AOI21D1 port map( A1 => N2920, A2 => N2921, B => 
                           mult_21_C241_n1401, Z => mult_21_C241_n950);
   mult_21_C241_U1389 : AOI21D1 port map( A1 => N2922, A2 => N2923, B => 
                           mult_21_C241_n1403, Z => mult_21_C241_n949);
   mult_21_C241_U1388 : AOI21D1 port map( A1 => N2924, A2 => N2925, B => 
                           mult_21_C241_n1405, Z => mult_21_C241_n948);
   mult_21_C241_U1387 : AOI21D1 port map( A1 => N2926, A2 => N2927, B => 
                           mult_21_C241_n1407, Z => mult_21_C241_n947);
   mult_21_C241_U1386 : EXOR2D1 port map( A1 => N2943, A2 => N2942, Z => 
                           mult_21_C241_n1451);
   mult_21_C241_U1385 : MUXB2DL port map( A0 => N3073, A1 => N3074, SL => 
                           mult_21_C241_n1451, Z => mult_21_C241_n652);
   mult_21_C241_U1384 : NAN2D1 port map( A1 => N3073, A2 => mult_21_C241_n1451,
                           Z => mult_21_C241_n653);
   mult_21_C241_U1383 : EXOR2D1 port map( A1 => N2941, A2 => N2940, Z => 
                           mult_21_C241_n1450);
   mult_21_C241_U1382 : MUXB2DL port map( A0 => N3075, A1 => N3076, SL => 
                           mult_21_C241_n1450, Z => mult_21_C241_n654);
   mult_21_C241_U1381 : MUXB2DL port map( A0 => mult_21_C241_n1388, A1 => N3075
                           , SL => mult_21_C241_n1450, Z => mult_21_C241_n655);
   mult_21_C241_U1380 : MUXB2DL port map( A0 => N3073, A1 => N3074, SL => 
                           mult_21_C241_n1450, Z => mult_21_C241_n656);
   mult_21_C241_U1379 : NAN2D1 port map( A1 => N3073, A2 => mult_21_C241_n1450,
                           Z => mult_21_C241_n657);
   mult_21_C241_U1378 : EXOR2D1 port map( A1 => N2939, A2 => N2938, Z => 
                           mult_21_C241_n1449);
   mult_21_C241_U1377 : MUXB2DL port map( A0 => N3077, A1 => N3078, SL => 
                           mult_21_C241_n1449, Z => mult_21_C241_n658);
   mult_21_C241_U1376 : MUXB2DL port map( A0 => mult_21_C241_n1386, A1 => N3077
                           , SL => mult_21_C241_n1449, Z => mult_21_C241_n659);
   mult_21_C241_U1375 : MUXB2DL port map( A0 => N3075, A1 => N3076, SL => 
                           mult_21_C241_n1449, Z => mult_21_C241_n660);
   mult_21_C241_U1374 : MUXB2DL port map( A0 => mult_21_C241_n1388, A1 => N3075
                           , SL => mult_21_C241_n1449, Z => mult_21_C241_n661);
   mult_21_C241_U1373 : MUXB2DL port map( A0 => N3073, A1 => N3074, SL => 
                           mult_21_C241_n1449, Z => mult_21_C241_n662);
   mult_21_C241_U1372 : NAN2D1 port map( A1 => N3073, A2 => mult_21_C241_n1449,
                           Z => mult_21_C241_n663);
   mult_21_C241_U1371 : EXOR2D1 port map( A1 => N2937, A2 => N2936, Z => 
                           mult_21_C241_n1448);
   mult_21_C241_U1370 : MUXB2DL port map( A0 => N3079, A1 => N3080, SL => 
                           mult_21_C241_n1448, Z => mult_21_C241_n664);
   mult_21_C241_U1369 : MUXB2DL port map( A0 => N3078, A1 => N3079, SL => 
                           mult_21_C241_n1448, Z => mult_21_C241_n665);
   mult_21_C241_U1368 : MUXB2DL port map( A0 => N3077, A1 => N3078, SL => 
                           mult_21_C241_n1448, Z => mult_21_C241_n666);
   mult_21_C241_U1367 : MUXB2DL port map( A0 => mult_21_C241_n1386, A1 => N3077
                           , SL => mult_21_C241_n1448, Z => mult_21_C241_n667);
   mult_21_C241_U1366 : MUXB2DL port map( A0 => N3075, A1 => N3076, SL => 
                           mult_21_C241_n1448, Z => mult_21_C241_n668);
   mult_21_C241_U1365 : MUXB2DL port map( A0 => mult_21_C241_n1388, A1 => N3075
                           , SL => mult_21_C241_n1448, Z => mult_21_C241_n669);
   mult_21_C241_U1364 : MUXB2DL port map( A0 => N3073, A1 => N3074, SL => 
                           mult_21_C241_n1448, Z => mult_21_C241_n670);
   mult_21_C241_U1363 : NAN2D1 port map( A1 => N3073, A2 => mult_21_C241_n1448,
                           Z => mult_21_C241_n671);
   mult_21_C241_U1362 : MUXB2DL port map( A0 => N3081, A1 => N3082, SL => 
                           mult_21_C241_n1447, Z => mult_21_C241_n672);
   mult_21_C241_U1361 : MUXB2DL port map( A0 => N3080, A1 => N3081, SL => 
                           mult_21_C241_n1447, Z => mult_21_C241_n673);
   mult_21_C241_U1360 : MUXB2DL port map( A0 => N3079, A1 => N3080, SL => 
                           mult_21_C241_n1447, Z => mult_21_C241_n674);
   mult_21_C241_U1359 : MUXB2DL port map( A0 => N3078, A1 => N3079, SL => 
                           mult_21_C241_n1447, Z => mult_21_C241_n675);
   mult_21_C241_U1358 : MUXB2DL port map( A0 => N3077, A1 => N3078, SL => 
                           mult_21_C241_n1447, Z => mult_21_C241_n676);
   mult_21_C241_U1357 : MUXB2DL port map( A0 => mult_21_C241_n1386, A1 => N3077
                           , SL => mult_21_C241_n1447, Z => mult_21_C241_n677);
   mult_21_C241_U1356 : MUXB2DL port map( A0 => N3075, A1 => N3076, SL => 
                           mult_21_C241_n1447, Z => mult_21_C241_n678);
   mult_21_C241_U1355 : MUXB2DL port map( A0 => mult_21_C241_n1388, A1 => N3075
                           , SL => mult_21_C241_n1447, Z => mult_21_C241_n679);
   mult_21_C241_U1354 : AOI21D1 port map( A1 => N2928, A2 => N2929, B => 
                           mult_21_C241_n1409, Z => mult_21_C241_n946);
   mult_21_C241_U1353 : MUXB2DL port map( A0 => N3073, A1 => N3074, SL => 
                           mult_21_C241_n1447, Z => mult_21_C241_n680);
   mult_21_C241_U1352 : NAN2D1 port map( A1 => N3073, A2 => mult_21_C241_n1447,
                           Z => mult_21_C241_n681);
   mult_21_C241_U1351 : MUXB2DL port map( A0 => N3083, A1 => N3084, SL => 
                           mult_21_C241_n1446, Z => mult_21_C241_n682);
   mult_21_C241_U1350 : MUXB2DL port map( A0 => N3082, A1 => N3083, SL => 
                           mult_21_C241_n1446, Z => mult_21_C241_n683);
   mult_21_C241_U1349 : MUXB2DL port map( A0 => N3081, A1 => N3082, SL => 
                           mult_21_C241_n1446, Z => mult_21_C241_n684);
   mult_21_C241_U1348 : MUXB2DL port map( A0 => N3080, A1 => N3081, SL => 
                           mult_21_C241_n1446, Z => mult_21_C241_n685);
   mult_21_C241_U1347 : MUXB2DL port map( A0 => N3079, A1 => N3080, SL => 
                           mult_21_C241_n1446, Z => mult_21_C241_n686);
   mult_21_C241_U1346 : MUXB2DL port map( A0 => N3078, A1 => N3079, SL => 
                           mult_21_C241_n1446, Z => mult_21_C241_n687);
   mult_21_C241_U1345 : MUXB2DL port map( A0 => N3077, A1 => N3078, SL => 
                           mult_21_C241_n1446, Z => mult_21_C241_n688);
   mult_21_C241_U1344 : MUXB2DL port map( A0 => mult_21_C241_n1386, A1 => N3077
                           , SL => mult_21_C241_n1446, Z => mult_21_C241_n689);
   mult_21_C241_U1343 : MUXB2DL port map( A0 => N3075, A1 => N3076, SL => 
                           mult_21_C241_n1446, Z => mult_21_C241_n690);
   mult_21_C241_U1342 : MUXB2DL port map( A0 => mult_21_C241_n1388, A1 => N3075
                           , SL => mult_21_C241_n1446, Z => mult_21_C241_n691);
   mult_21_C241_U1341 : MUXB2DL port map( A0 => N3073, A1 => N3074, SL => 
                           mult_21_C241_n1446, Z => mult_21_C241_n692);
   mult_21_C241_U1340 : NAN2D1 port map( A1 => N3073, A2 => mult_21_C241_n1446,
                           Z => mult_21_C241_n693);
   mult_21_C241_U1339 : MUXB2DL port map( A0 => N3085, A1 => N3086, SL => 
                           mult_21_C241_n1445, Z => mult_21_C241_n694);
   mult_21_C241_U1338 : MUXB2DL port map( A0 => N3084, A1 => N3085, SL => 
                           mult_21_C241_n1445, Z => mult_21_C241_n695);
   mult_21_C241_U1337 : MUXB2DL port map( A0 => N3083, A1 => N3084, SL => 
                           mult_21_C241_n1445, Z => mult_21_C241_n696);
   mult_21_C241_U1336 : MUXB2DL port map( A0 => N3082, A1 => N3083, SL => 
                           mult_21_C241_n1445, Z => mult_21_C241_n697);
   mult_21_C241_U1335 : MUXB2DL port map( A0 => N3081, A1 => N3082, SL => 
                           mult_21_C241_n1445, Z => mult_21_C241_n698);
   mult_21_C241_U1334 : MUXB2DL port map( A0 => N3080, A1 => N3081, SL => 
                           mult_21_C241_n1445, Z => mult_21_C241_n699);
   mult_21_C241_U1333 : MUXB2DL port map( A0 => N3079, A1 => N3080, SL => 
                           mult_21_C241_n1445, Z => mult_21_C241_n700);
   mult_21_C241_U1332 : MUXB2DL port map( A0 => N3078, A1 => N3079, SL => 
                           mult_21_C241_n1445, Z => mult_21_C241_n701);
   mult_21_C241_U1331 : MUXB2DL port map( A0 => N3077, A1 => N3078, SL => 
                           mult_21_C241_n1445, Z => mult_21_C241_n702);
   mult_21_C241_U1330 : MUXB2DL port map( A0 => mult_21_C241_n1386, A1 => N3077
                           , SL => mult_21_C241_n1445, Z => mult_21_C241_n703);
   mult_21_C241_U1329 : MUXB2DL port map( A0 => N3075, A1 => N3076, SL => 
                           mult_21_C241_n1445, Z => mult_21_C241_n704);
   mult_21_C241_U1328 : MUXB2DL port map( A0 => mult_21_C241_n1388, A1 => N3075
                           , SL => mult_21_C241_n1445, Z => mult_21_C241_n705);
   mult_21_C241_U1327 : MUXB2DL port map( A0 => N3073, A1 => N3074, SL => 
                           mult_21_C241_n1445, Z => mult_21_C241_n706);
   mult_21_C241_U1326 : NAN2D1 port map( A1 => N3073, A2 => mult_21_C241_n1445,
                           Z => mult_21_C241_n707);
   mult_21_C241_U1325 : MUXB2DL port map( A0 => N3087, A1 => N3088, SL => 
                           mult_21_C241_n1444, Z => mult_21_C241_n708);
   mult_21_C241_U1324 : MUXB2DL port map( A0 => N3086, A1 => N3087, SL => 
                           mult_21_C241_n1444, Z => mult_21_C241_n709);
   mult_21_C241_U1323 : MUXB2DL port map( A0 => N3085, A1 => N3086, SL => 
                           mult_21_C241_n1444, Z => mult_21_C241_n710);
   mult_21_C241_U1322 : MUXB2DL port map( A0 => N3084, A1 => N3085, SL => 
                           mult_21_C241_n1444, Z => mult_21_C241_n711);
   mult_21_C241_U1321 : MUXB2DL port map( A0 => N3083, A1 => N3084, SL => 
                           mult_21_C241_n1444, Z => mult_21_C241_n712);
   mult_21_C241_U1320 : MUXB2DL port map( A0 => N3082, A1 => N3083, SL => 
                           mult_21_C241_n1444, Z => mult_21_C241_n713);
   mult_21_C241_U1319 : MUXB2DL port map( A0 => N3081, A1 => N3082, SL => 
                           mult_21_C241_n1444, Z => mult_21_C241_n714);
   mult_21_C241_U1318 : MUXB2DL port map( A0 => N3080, A1 => N3081, SL => 
                           mult_21_C241_n1444, Z => mult_21_C241_n715);
   mult_21_C241_U1317 : MUXB2DL port map( A0 => N3079, A1 => N3080, SL => 
                           mult_21_C241_n1444, Z => mult_21_C241_n716);
   mult_21_C241_U1316 : MUXB2DL port map( A0 => N3078, A1 => N3079, SL => 
                           mult_21_C241_n1444, Z => mult_21_C241_n717);
   mult_21_C241_U1315 : MUXB2DL port map( A0 => N3077, A1 => N3078, SL => 
                           mult_21_C241_n1444, Z => mult_21_C241_n718);
   mult_21_C241_U1314 : MUXB2DL port map( A0 => mult_21_C241_n1386, A1 => N3077
                           , SL => mult_21_C241_n1444, Z => mult_21_C241_n719);
   mult_21_C241_U1313 : MUXB2DL port map( A0 => N3075, A1 => N3076, SL => 
                           mult_21_C241_n1444, Z => mult_21_C241_n720);
   mult_21_C241_U1312 : MUXB2DL port map( A0 => mult_21_C241_n1388, A1 => N3075
                           , SL => mult_21_C241_n1444, Z => mult_21_C241_n721);
   mult_21_C241_U1311 : MUXB2DL port map( A0 => N3073, A1 => N3074, SL => 
                           mult_21_C241_n1444, Z => mult_21_C241_n722);
   mult_21_C241_U1310 : NAN2D1 port map( A1 => N3073, A2 => mult_21_C241_n1444,
                           Z => mult_21_C241_n723);
   mult_21_C241_U1309 : MUXB2DL port map( A0 => N3089, A1 => N3090, SL => 
                           mult_21_C241_n1443, Z => mult_21_C241_n724);
   mult_21_C241_U1308 : MUXB2DL port map( A0 => N3088, A1 => N3089, SL => 
                           mult_21_C241_n1443, Z => mult_21_C241_n725);
   mult_21_C241_U1307 : MUXB2DL port map( A0 => N3087, A1 => N3088, SL => 
                           mult_21_C241_n1443, Z => mult_21_C241_n726);
   mult_21_C241_U1306 : MUXB2DL port map( A0 => N3086, A1 => N3087, SL => 
                           mult_21_C241_n1443, Z => mult_21_C241_n727);
   mult_21_C241_U1305 : MUXB2DL port map( A0 => N3085, A1 => N3086, SL => 
                           mult_21_C241_n1443, Z => mult_21_C241_n728);
   mult_21_C241_U1304 : MUXB2DL port map( A0 => N3084, A1 => N3085, SL => 
                           mult_21_C241_n1443, Z => mult_21_C241_n729);
   mult_21_C241_U1303 : MUXB2DL port map( A0 => N3083, A1 => N3084, SL => 
                           mult_21_C241_n1443, Z => mult_21_C241_n730);
   mult_21_C241_U1302 : MUXB2DL port map( A0 => N3082, A1 => N3083, SL => 
                           mult_21_C241_n1443, Z => mult_21_C241_n731);
   mult_21_C241_U1301 : MUXB2DL port map( A0 => N3081, A1 => N3082, SL => 
                           mult_21_C241_n1443, Z => mult_21_C241_n732);
   mult_21_C241_U1300 : MUXB2DL port map( A0 => N3080, A1 => N3081, SL => 
                           mult_21_C241_n1443, Z => mult_21_C241_n733);
   mult_21_C241_U1299 : MUXB2DL port map( A0 => N3079, A1 => N3080, SL => 
                           mult_21_C241_n1443, Z => mult_21_C241_n734);
   mult_21_C241_U1298 : MUXB2DL port map( A0 => N3078, A1 => N3079, SL => 
                           mult_21_C241_n1443, Z => mult_21_C241_n735);
   mult_21_C241_U1297 : MUXB2DL port map( A0 => N3077, A1 => N3078, SL => 
                           mult_21_C241_n1443, Z => mult_21_C241_n736);
   mult_21_C241_U1296 : MUXB2DL port map( A0 => mult_21_C241_n1386, A1 => N3077
                           , SL => mult_21_C241_n1443, Z => mult_21_C241_n737);
   mult_21_C241_U1295 : MUXB2DL port map( A0 => N3075, A1 => N3076, SL => 
                           mult_21_C241_n1443, Z => mult_21_C241_n738);
   mult_21_C241_U1294 : MUXB2DL port map( A0 => mult_21_C241_n1388, A1 => N3075
                           , SL => mult_21_C241_n1443, Z => mult_21_C241_n739);
   mult_21_C241_U1293 : MUXB2DL port map( A0 => N3073, A1 => N3074, SL => 
                           mult_21_C241_n1443, Z => mult_21_C241_n740);
   mult_21_C241_U1292 : NAN2D1 port map( A1 => N3073, A2 => mult_21_C241_n1443,
                           Z => mult_21_C241_n741);
   mult_21_C241_U1291 : MUXB2DL port map( A0 => N3091, A1 => N3092, SL => 
                           mult_21_C241_n1442, Z => mult_21_C241_n742);
   mult_21_C241_U1290 : MUXB2DL port map( A0 => N3090, A1 => N3091, SL => 
                           mult_21_C241_n1442, Z => mult_21_C241_n743);
   mult_21_C241_U1289 : MUXB2DL port map( A0 => N3089, A1 => N3090, SL => 
                           mult_21_C241_n1442, Z => mult_21_C241_n744);
   mult_21_C241_U1288 : MUXB2DL port map( A0 => N3088, A1 => N3089, SL => 
                           mult_21_C241_n1442, Z => mult_21_C241_n745);
   mult_21_C241_U1287 : MUXB2DL port map( A0 => N3087, A1 => N3088, SL => 
                           mult_21_C241_n1442, Z => mult_21_C241_n746);
   mult_21_C241_U1286 : MUXB2DL port map( A0 => N3086, A1 => N3087, SL => 
                           mult_21_C241_n1442, Z => mult_21_C241_n747);
   mult_21_C241_U1285 : MUXB2DL port map( A0 => N3085, A1 => N3086, SL => 
                           mult_21_C241_n1442, Z => mult_21_C241_n748);
   mult_21_C241_U1284 : MUXB2DL port map( A0 => N3084, A1 => N3085, SL => 
                           mult_21_C241_n1442, Z => mult_21_C241_n749);
   mult_21_C241_U1283 : AOI21D1 port map( A1 => N2930, A2 => N2931, B => 
                           mult_21_C241_n1411, Z => mult_21_C241_n945);
   mult_21_C241_U1282 : MUXB2DL port map( A0 => N3083, A1 => N3084, SL => 
                           mult_21_C241_n1442, Z => mult_21_C241_n750);
   mult_21_C241_U1281 : MUXB2DL port map( A0 => N3082, A1 => N3083, SL => 
                           mult_21_C241_n1442, Z => mult_21_C241_n751);
   mult_21_C241_U1280 : MUXB2DL port map( A0 => N3081, A1 => N3082, SL => 
                           mult_21_C241_n1442, Z => mult_21_C241_n752);
   mult_21_C241_U1279 : MUXB2DL port map( A0 => N3080, A1 => N3081, SL => 
                           mult_21_C241_n1442, Z => mult_21_C241_n753);
   mult_21_C241_U1278 : MUXB2DL port map( A0 => N3079, A1 => N3080, SL => 
                           mult_21_C241_n1442, Z => mult_21_C241_n754);
   mult_21_C241_U1277 : MUXB2DL port map( A0 => N3078, A1 => N3079, SL => 
                           mult_21_C241_n1442, Z => mult_21_C241_n755);
   mult_21_C241_U1276 : MUXB2DL port map( A0 => N3077, A1 => N3078, SL => 
                           mult_21_C241_n1442, Z => mult_21_C241_n756);
   mult_21_C241_U1275 : MUXB2DL port map( A0 => mult_21_C241_n1386, A1 => N3077
                           , SL => mult_21_C241_n1442, Z => mult_21_C241_n757);
   mult_21_C241_U1274 : MUXB2DL port map( A0 => N3075, A1 => N3076, SL => 
                           mult_21_C241_n1442, Z => mult_21_C241_n758);
   mult_21_C241_U1273 : MUXB2DL port map( A0 => N3074, A1 => N3075, SL => 
                           mult_21_C241_n1442, Z => mult_21_C241_n759);
   mult_21_C241_U1272 : MUXB2DL port map( A0 => N3073, A1 => N3074, SL => 
                           mult_21_C241_n1442, Z => mult_21_C241_n760);
   mult_21_C241_U1271 : NAN2D1 port map( A1 => N3073, A2 => mult_21_C241_n1442,
                           Z => mult_21_C241_n761);
   mult_21_C241_U1270 : MUXB2DL port map( A0 => N3093, A1 => N3094, SL => 
                           mult_21_C241_n1441, Z => mult_21_C241_n762);
   mult_21_C241_U1269 : MUXB2DL port map( A0 => N3092, A1 => N3093, SL => 
                           mult_21_C241_n1441, Z => mult_21_C241_n763);
   mult_21_C241_U1268 : MUXB2DL port map( A0 => N3091, A1 => N3092, SL => 
                           mult_21_C241_n1441, Z => mult_21_C241_n764);
   mult_21_C241_U1267 : MUXB2DL port map( A0 => N3090, A1 => N3091, SL => 
                           mult_21_C241_n1441, Z => mult_21_C241_n765);
   mult_21_C241_U1266 : MUXB2DL port map( A0 => N3089, A1 => N3090, SL => 
                           mult_21_C241_n1441, Z => mult_21_C241_n766);
   mult_21_C241_U1265 : MUXB2DL port map( A0 => N3088, A1 => N3089, SL => 
                           mult_21_C241_n1441, Z => mult_21_C241_n767);
   mult_21_C241_U1264 : MUXB2DL port map( A0 => N3087, A1 => N3088, SL => 
                           mult_21_C241_n1441, Z => mult_21_C241_n768);
   mult_21_C241_U1263 : MUXB2DL port map( A0 => N3086, A1 => N3087, SL => 
                           mult_21_C241_n1441, Z => mult_21_C241_n769);
   mult_21_C241_U1262 : MUXB2DL port map( A0 => N3085, A1 => N3086, SL => 
                           mult_21_C241_n1441, Z => mult_21_C241_n770);
   mult_21_C241_U1261 : MUXB2DL port map( A0 => N3084, A1 => N3085, SL => 
                           mult_21_C241_n1441, Z => mult_21_C241_n771);
   mult_21_C241_U1260 : MUXB2DL port map( A0 => N3083, A1 => N3084, SL => 
                           mult_21_C241_n1441, Z => mult_21_C241_n772);
   mult_21_C241_U1259 : MUXB2DL port map( A0 => N3082, A1 => N3083, SL => 
                           mult_21_C241_n1441, Z => mult_21_C241_n773);
   mult_21_C241_U1258 : MUXB2DL port map( A0 => N3081, A1 => N3082, SL => 
                           mult_21_C241_n1441, Z => mult_21_C241_n774);
   mult_21_C241_U1257 : MUXB2DL port map( A0 => N3080, A1 => N3081, SL => 
                           mult_21_C241_n1441, Z => mult_21_C241_n775);
   mult_21_C241_U1256 : MUXB2DL port map( A0 => N3079, A1 => N3080, SL => 
                           mult_21_C241_n1441, Z => mult_21_C241_n776);
   mult_21_C241_U1255 : MUXB2DL port map( A0 => N3078, A1 => N3079, SL => 
                           mult_21_C241_n1441, Z => mult_21_C241_n777);
   mult_21_C241_U1254 : MUXB2DL port map( A0 => N3077, A1 => N3078, SL => 
                           mult_21_C241_n1441, Z => mult_21_C241_n778);
   mult_21_C241_U1253 : MUXB2DL port map( A0 => N3076, A1 => N3077, SL => 
                           mult_21_C241_n1441, Z => mult_21_C241_n779);
   mult_21_C241_U1252 : MUXB2DL port map( A0 => N3075, A1 => N3076, SL => 
                           mult_21_C241_n1441, Z => mult_21_C241_n780);
   mult_21_C241_U1251 : MUXB2DL port map( A0 => mult_21_C241_n1388, A1 => N3075
                           , SL => mult_21_C241_n1441, Z => mult_21_C241_n781);
   mult_21_C241_U1250 : MUXB2DL port map( A0 => N3073, A1 => N3074, SL => 
                           mult_21_C241_n1441, Z => mult_21_C241_n782);
   mult_21_C241_U1249 : NAN2D1 port map( A1 => N3073, A2 => mult_21_C241_n1441,
                           Z => mult_21_C241_n783);
   mult_21_C241_U1248 : MUXB2DL port map( A0 => N3095, A1 => N3096, SL => 
                           mult_21_C241_n1379, Z => mult_21_C241_n784);
   mult_21_C241_U1247 : MUXB2DL port map( A0 => N3094, A1 => N3095, SL => 
                           mult_21_C241_n1379, Z => mult_21_C241_n785);
   mult_21_C241_U1246 : MUXB2DL port map( A0 => N3093, A1 => N3094, SL => 
                           mult_21_C241_n1379, Z => mult_21_C241_n786);
   mult_21_C241_U1245 : MUXB2DL port map( A0 => N3092, A1 => N3093, SL => 
                           mult_21_C241_n1379, Z => mult_21_C241_n787);
   mult_21_C241_U1244 : MUXB2DL port map( A0 => N3091, A1 => N3092, SL => 
                           mult_21_C241_n1379, Z => mult_21_C241_n788);
   mult_21_C241_U1243 : MUXB2DL port map( A0 => N3090, A1 => N3091, SL => 
                           mult_21_C241_n1379, Z => mult_21_C241_n789);
   mult_21_C241_U1242 : MUXB2DL port map( A0 => N3089, A1 => N3090, SL => 
                           mult_21_C241_n1379, Z => mult_21_C241_n790);
   mult_21_C241_U1241 : MUXB2DL port map( A0 => N3088, A1 => N3089, SL => 
                           mult_21_C241_n1379, Z => mult_21_C241_n791);
   mult_21_C241_U1240 : MUXB2DL port map( A0 => N3087, A1 => N3088, SL => 
                           mult_21_C241_n1379, Z => mult_21_C241_n792);
   mult_21_C241_U1239 : MUXB2DL port map( A0 => N3086, A1 => N3087, SL => 
                           mult_21_C241_n1379, Z => mult_21_C241_n793);
   mult_21_C241_U1238 : MUXB2DL port map( A0 => N3085, A1 => N3086, SL => 
                           mult_21_C241_n1379, Z => mult_21_C241_n794);
   mult_21_C241_U1237 : MUXB2DL port map( A0 => N3084, A1 => N3085, SL => 
                           mult_21_C241_n1379, Z => mult_21_C241_n795);
   mult_21_C241_U1236 : MUXB2DL port map( A0 => N3083, A1 => N3084, SL => 
                           mult_21_C241_n1379, Z => mult_21_C241_n796);
   mult_21_C241_U1235 : MUXB2DL port map( A0 => N3082, A1 => N3083, SL => 
                           mult_21_C241_n1379, Z => mult_21_C241_n797);
   mult_21_C241_U1234 : MUXB2DL port map( A0 => N3081, A1 => N3082, SL => 
                           mult_21_C241_n1379, Z => mult_21_C241_n798);
   mult_21_C241_U1233 : MUXB2DL port map( A0 => N3080, A1 => N3081, SL => 
                           mult_21_C241_n1379, Z => mult_21_C241_n799);
   mult_21_C241_U1232 : MUXB2DL port map( A0 => N3079, A1 => N3080, SL => 
                           mult_21_C241_n1379, Z => mult_21_C241_n800);
   mult_21_C241_U1231 : MUXB2DL port map( A0 => N3078, A1 => N3079, SL => 
                           mult_21_C241_n1379, Z => mult_21_C241_n801);
   mult_21_C241_U1230 : MUXB2DL port map( A0 => N3077, A1 => N3078, SL => 
                           mult_21_C241_n1379, Z => mult_21_C241_n802);
   mult_21_C241_U1229 : MUXB2DL port map( A0 => mult_21_C241_n1386, A1 => N3077
                           , SL => mult_21_C241_n1379, Z => mult_21_C241_n803);
   mult_21_C241_U1228 : MUXB2DL port map( A0 => N3075, A1 => N3076, SL => 
                           mult_21_C241_n1379, Z => mult_21_C241_n804);
   mult_21_C241_U1227 : MUXB2DL port map( A0 => N3074, A1 => N3075, SL => 
                           mult_21_C241_n1379, Z => mult_21_C241_n805);
   mult_21_C241_U1226 : MUXB2DL port map( A0 => N3073, A1 => N3074, SL => 
                           mult_21_C241_n1379, Z => mult_21_C241_n806);
   mult_21_C241_U1225 : NAN2D1 port map( A1 => N3073, A2 => mult_21_C241_n1379,
                           Z => mult_21_C241_n807);
   mult_21_C241_U1224 : MUXB2DL port map( A0 => N3097, A1 => N3098, SL => 
                           mult_21_C241_n1378, Z => mult_21_C241_n808);
   mult_21_C241_U1223 : MUXB2DL port map( A0 => N3096, A1 => N3097, SL => 
                           mult_21_C241_n1378, Z => mult_21_C241_n809);
   mult_21_C241_U1222 : AOI21D1 port map( A1 => N2932, A2 => N2933, B => 
                           mult_21_C241_n1413, Z => mult_21_C241_n944);
   mult_21_C241_U1221 : MUXB2DL port map( A0 => N3095, A1 => N3096, SL => 
                           mult_21_C241_n1378, Z => mult_21_C241_n810);
   mult_21_C241_U1220 : MUXB2DL port map( A0 => N3094, A1 => N3095, SL => 
                           mult_21_C241_n1378, Z => mult_21_C241_n811);
   mult_21_C241_U1219 : MUXB2DL port map( A0 => N3093, A1 => N3094, SL => 
                           mult_21_C241_n1378, Z => mult_21_C241_n812);
   mult_21_C241_U1218 : MUXB2DL port map( A0 => N3092, A1 => N3093, SL => 
                           mult_21_C241_n1378, Z => mult_21_C241_n813);
   mult_21_C241_U1217 : MUXB2DL port map( A0 => N3091, A1 => N3092, SL => 
                           mult_21_C241_n1378, Z => mult_21_C241_n814);
   mult_21_C241_U1216 : MUXB2DL port map( A0 => N3090, A1 => N3091, SL => 
                           mult_21_C241_n1378, Z => mult_21_C241_n815);
   mult_21_C241_U1215 : MUXB2DL port map( A0 => N3089, A1 => N3090, SL => 
                           mult_21_C241_n1378, Z => mult_21_C241_n816);
   mult_21_C241_U1214 : MUXB2DL port map( A0 => N3088, A1 => N3089, SL => 
                           mult_21_C241_n1378, Z => mult_21_C241_n817);
   mult_21_C241_U1213 : MUXB2DL port map( A0 => N3087, A1 => N3088, SL => 
                           mult_21_C241_n1378, Z => mult_21_C241_n818);
   mult_21_C241_U1212 : MUXB2DL port map( A0 => N3086, A1 => N3087, SL => 
                           mult_21_C241_n1378, Z => mult_21_C241_n819);
   mult_21_C241_U1211 : MUXB2DL port map( A0 => N3085, A1 => N3086, SL => 
                           mult_21_C241_n1378, Z => mult_21_C241_n820);
   mult_21_C241_U1210 : MUXB2DL port map( A0 => N3084, A1 => N3085, SL => 
                           mult_21_C241_n1378, Z => mult_21_C241_n821);
   mult_21_C241_U1209 : MUXB2DL port map( A0 => N3083, A1 => N3084, SL => 
                           mult_21_C241_n1378, Z => mult_21_C241_n822);
   mult_21_C241_U1208 : MUXB2DL port map( A0 => N3082, A1 => N3083, SL => 
                           mult_21_C241_n1378, Z => mult_21_C241_n823);
   mult_21_C241_U1207 : MUXB2DL port map( A0 => N3081, A1 => N3082, SL => 
                           mult_21_C241_n1378, Z => mult_21_C241_n824);
   mult_21_C241_U1206 : MUXB2DL port map( A0 => N3080, A1 => N3081, SL => 
                           mult_21_C241_n1378, Z => mult_21_C241_n825);
   mult_21_C241_U1205 : MUXB2DL port map( A0 => N3079, A1 => N3080, SL => 
                           mult_21_C241_n1378, Z => mult_21_C241_n826);
   mult_21_C241_U1204 : MUXB2DL port map( A0 => N3078, A1 => N3079, SL => 
                           mult_21_C241_n1378, Z => mult_21_C241_n827);
   mult_21_C241_U1203 : MUXB2DL port map( A0 => N3077, A1 => N3078, SL => 
                           mult_21_C241_n1378, Z => mult_21_C241_n828);
   mult_21_C241_U1202 : MUXB2DL port map( A0 => mult_21_C241_n1386, A1 => N3077
                           , SL => mult_21_C241_n1378, Z => mult_21_C241_n829);
   mult_21_C241_U1201 : MUXB2DL port map( A0 => N3075, A1 => N3076, SL => 
                           mult_21_C241_n1378, Z => mult_21_C241_n830);
   mult_21_C241_U1200 : MUXB2DL port map( A0 => mult_21_C241_n1388, A1 => N3075
                           , SL => mult_21_C241_n1378, Z => mult_21_C241_n831);
   mult_21_C241_U1199 : MUXB2DL port map( A0 => N3073, A1 => N3074, SL => 
                           mult_21_C241_n1378, Z => mult_21_C241_n832);
   mult_21_C241_U1198 : NAN2D1 port map( A1 => N3073, A2 => mult_21_C241_n1378,
                           Z => mult_21_C241_n833);
   mult_21_C241_U1197 : MUXB2DL port map( A0 => N3099, A1 => N3100, SL => 
                           mult_21_C241_n1385, Z => mult_21_C241_n834);
   mult_21_C241_U1196 : MUXB2DL port map( A0 => N3098, A1 => N3099, SL => 
                           mult_21_C241_n1385, Z => mult_21_C241_n835);
   mult_21_C241_U1195 : MUXB2DL port map( A0 => N3097, A1 => N3098, SL => 
                           mult_21_C241_n1385, Z => mult_21_C241_n836);
   mult_21_C241_U1194 : MUXB2DL port map( A0 => N3096, A1 => N3097, SL => 
                           mult_21_C241_n1385, Z => mult_21_C241_n837);
   mult_21_C241_U1193 : MUXB2DL port map( A0 => N3095, A1 => N3096, SL => 
                           mult_21_C241_n1385, Z => mult_21_C241_n838);
   mult_21_C241_U1192 : MUXB2DL port map( A0 => N3094, A1 => N3095, SL => 
                           mult_21_C241_n1385, Z => mult_21_C241_n839);
   mult_21_C241_U1191 : MUXB2DL port map( A0 => N3093, A1 => N3094, SL => 
                           mult_21_C241_n1385, Z => mult_21_C241_n840);
   mult_21_C241_U1190 : MUXB2DL port map( A0 => N3092, A1 => N3093, SL => 
                           mult_21_C241_n1385, Z => mult_21_C241_n841);
   mult_21_C241_U1189 : MUXB2DL port map( A0 => N3091, A1 => N3092, SL => 
                           mult_21_C241_n1385, Z => mult_21_C241_n842);
   mult_21_C241_U1188 : MUXB2DL port map( A0 => N3090, A1 => N3091, SL => 
                           mult_21_C241_n1385, Z => mult_21_C241_n843);
   mult_21_C241_U1187 : MUXB2DL port map( A0 => N3089, A1 => N3090, SL => 
                           mult_21_C241_n1385, Z => mult_21_C241_n844);
   mult_21_C241_U1186 : MUXB2DL port map( A0 => N3088, A1 => N3089, SL => 
                           mult_21_C241_n1385, Z => mult_21_C241_n845);
   mult_21_C241_U1185 : MUXB2DL port map( A0 => N3087, A1 => N3088, SL => 
                           mult_21_C241_n1385, Z => mult_21_C241_n846);
   mult_21_C241_U1184 : MUXB2DL port map( A0 => N3086, A1 => N3087, SL => 
                           mult_21_C241_n1385, Z => mult_21_C241_n847);
   mult_21_C241_U1183 : MUXB2DL port map( A0 => N3085, A1 => N3086, SL => 
                           mult_21_C241_n1385, Z => mult_21_C241_n848);
   mult_21_C241_U1182 : MUXB2DL port map( A0 => N3084, A1 => N3085, SL => 
                           mult_21_C241_n1385, Z => mult_21_C241_n849);
   mult_21_C241_U1181 : MUXB2DL port map( A0 => N3083, A1 => N3084, SL => 
                           mult_21_C241_n1385, Z => mult_21_C241_n850);
   mult_21_C241_U1180 : MUXB2DL port map( A0 => N3082, A1 => N3083, SL => 
                           mult_21_C241_n1385, Z => mult_21_C241_n851);
   mult_21_C241_U1179 : MUXB2DL port map( A0 => N3081, A1 => N3082, SL => 
                           mult_21_C241_n1385, Z => mult_21_C241_n852);
   mult_21_C241_U1178 : MUXB2DL port map( A0 => N3080, A1 => N3081, SL => 
                           mult_21_C241_n1385, Z => mult_21_C241_n853);
   mult_21_C241_U1177 : MUXB2DL port map( A0 => N3079, A1 => N3080, SL => 
                           mult_21_C241_n1385, Z => mult_21_C241_n854);
   mult_21_C241_U1176 : MUXB2DL port map( A0 => N3078, A1 => N3079, SL => 
                           mult_21_C241_n1385, Z => mult_21_C241_n855);
   mult_21_C241_U1175 : MUXB2DL port map( A0 => N3077, A1 => N3078, SL => 
                           mult_21_C241_n1385, Z => mult_21_C241_n856);
   mult_21_C241_U1174 : MUXB2DL port map( A0 => mult_21_C241_n1386, A1 => N3077
                           , SL => mult_21_C241_n1385, Z => mult_21_C241_n857);
   mult_21_C241_U1173 : MUXB2DL port map( A0 => N3075, A1 => N3076, SL => 
                           mult_21_C241_n1385, Z => mult_21_C241_n858);
   mult_21_C241_U1172 : MUXB2DL port map( A0 => mult_21_C241_n1388, A1 => N3075
                           , SL => mult_21_C241_n1385, Z => mult_21_C241_n859);
   mult_21_C241_U1171 : AOI21D1 port map( A1 => N2934, A2 => N2935, B => 
                           mult_21_C241_n1415, Z => mult_21_C241_n943);
   mult_21_C241_U1170 : MUXB2DL port map( A0 => N3073, A1 => N3074, SL => 
                           mult_21_C241_n1385, Z => mult_21_C241_n860);
   mult_21_C241_U1169 : NAN2D1 port map( A1 => N3073, A2 => mult_21_C241_n1385,
                           Z => mult_21_C241_n861);
   mult_21_C241_U1168 : MUXB2DL port map( A0 => N3100, A1 => N3101, SL => 
                           mult_21_C241_n1384, Z => mult_21_C241_n863);
   mult_21_C241_U1167 : MUXB2DL port map( A0 => N3099, A1 => N3100, SL => 
                           mult_21_C241_n1384, Z => mult_21_C241_n864);
   mult_21_C241_U1166 : MUXB2DL port map( A0 => N3098, A1 => N3099, SL => 
                           mult_21_C241_n1384, Z => mult_21_C241_n865);
   mult_21_C241_U1165 : MUXB2DL port map( A0 => N3097, A1 => N3098, SL => 
                           mult_21_C241_n1384, Z => mult_21_C241_n866);
   mult_21_C241_U1164 : MUXB2DL port map( A0 => N3096, A1 => N3097, SL => 
                           mult_21_C241_n1384, Z => mult_21_C241_n867);
   mult_21_C241_U1163 : MUXB2DL port map( A0 => N3095, A1 => N3096, SL => 
                           mult_21_C241_n1384, Z => mult_21_C241_n868);
   mult_21_C241_U1162 : MUXB2DL port map( A0 => N3094, A1 => N3095, SL => 
                           mult_21_C241_n1384, Z => mult_21_C241_n869);
   mult_21_C241_U1161 : MUXB2DL port map( A0 => N3093, A1 => N3094, SL => 
                           mult_21_C241_n1384, Z => mult_21_C241_n870);
   mult_21_C241_U1160 : MUXB2DL port map( A0 => N3092, A1 => N3093, SL => 
                           mult_21_C241_n1384, Z => mult_21_C241_n871);
   mult_21_C241_U1159 : MUXB2DL port map( A0 => N3091, A1 => N3092, SL => 
                           mult_21_C241_n1384, Z => mult_21_C241_n872);
   mult_21_C241_U1158 : MUXB2DL port map( A0 => N3090, A1 => N3091, SL => 
                           mult_21_C241_n1384, Z => mult_21_C241_n873);
   mult_21_C241_U1157 : MUXB2DL port map( A0 => N3089, A1 => N3090, SL => 
                           mult_21_C241_n1384, Z => mult_21_C241_n874);
   mult_21_C241_U1156 : MUXB2DL port map( A0 => N3088, A1 => N3089, SL => 
                           mult_21_C241_n1384, Z => mult_21_C241_n875);
   mult_21_C241_U1155 : MUXB2DL port map( A0 => N3087, A1 => N3088, SL => 
                           mult_21_C241_n1384, Z => mult_21_C241_n876);
   mult_21_C241_U1154 : MUXB2DL port map( A0 => N3086, A1 => N3087, SL => 
                           mult_21_C241_n1384, Z => mult_21_C241_n877);
   mult_21_C241_U1153 : MUXB2DL port map( A0 => N3085, A1 => N3086, SL => 
                           mult_21_C241_n1384, Z => mult_21_C241_n878);
   mult_21_C241_U1152 : MUXB2DL port map( A0 => N3084, A1 => N3085, SL => 
                           mult_21_C241_n1384, Z => mult_21_C241_n879);
   mult_21_C241_U1151 : MUXB2DL port map( A0 => N3083, A1 => N3084, SL => 
                           mult_21_C241_n1384, Z => mult_21_C241_n880);
   mult_21_C241_U1150 : MUXB2DL port map( A0 => N3082, A1 => N3083, SL => 
                           mult_21_C241_n1384, Z => mult_21_C241_n881);
   mult_21_C241_U1149 : MUXB2DL port map( A0 => N3081, A1 => N3082, SL => 
                           mult_21_C241_n1384, Z => mult_21_C241_n882);
   mult_21_C241_U1148 : MUXB2DL port map( A0 => N3080, A1 => N3081, SL => 
                           mult_21_C241_n1384, Z => mult_21_C241_n883);
   mult_21_C241_U1147 : MUXB2DL port map( A0 => N3079, A1 => N3080, SL => 
                           mult_21_C241_n1384, Z => mult_21_C241_n884);
   mult_21_C241_U1146 : MUXB2DL port map( A0 => N3078, A1 => N3079, SL => 
                           mult_21_C241_n1384, Z => mult_21_C241_n885);
   mult_21_C241_U1145 : MUXB2DL port map( A0 => N3077, A1 => N3078, SL => 
                           mult_21_C241_n1384, Z => mult_21_C241_n886);
   mult_21_C241_U1144 : MUXB2DL port map( A0 => mult_21_C241_n1386, A1 => N3077
                           , SL => mult_21_C241_n1384, Z => mult_21_C241_n887);
   mult_21_C241_U1143 : MUXB2DL port map( A0 => N3075, A1 => N3076, SL => 
                           mult_21_C241_n1384, Z => mult_21_C241_n888);
   mult_21_C241_U1142 : MUXB2DL port map( A0 => mult_21_C241_n1388, A1 => N3075
                           , SL => mult_21_C241_n1384, Z => mult_21_C241_n889);
   mult_21_C241_U1141 : OAI21D1 port map( A1 => N2937, A2 => N2936, B => 
                           mult_21_C241_n1417, Z => mult_21_C241_n89);
   mult_21_C241_U1140 : MUXB2DL port map( A0 => N3073, A1 => N3074, SL => 
                           mult_21_C241_n1384, Z => mult_21_C241_n890);
   mult_21_C241_U1139 : NAN2D1 port map( A1 => N3073, A2 => mult_21_C241_n1384,
                           Z => mult_21_C241_n891);
   mult_21_C241_U1138 : MUXB2DL port map( A0 => N3103, A1 => N3104, SL => 
                           mult_21_C241_n1390, Z => mult_21_C241_n892);
   mult_21_C241_U1137 : MUXB2DL port map( A0 => N3102, A1 => N3103, SL => N2913
                           , Z => mult_21_C241_n893);
   mult_21_C241_U1136 : MUXB2DL port map( A0 => N3101, A1 => N3102, SL => N2913
                           , Z => mult_21_C241_n894);
   mult_21_C241_U1135 : MUXB2DL port map( A0 => N3100, A1 => N3101, SL => N2913
                           , Z => mult_21_C241_n895);
   mult_21_C241_U1134 : MUXB2DL port map( A0 => N3099, A1 => N3100, SL => N2913
                           , Z => mult_21_C241_n896);
   mult_21_C241_U1133 : MUXB2DL port map( A0 => N3098, A1 => N3099, SL => N2913
                           , Z => mult_21_C241_n897);
   mult_21_C241_U1132 : MUXB2DL port map( A0 => N3097, A1 => N3098, SL => N2913
                           , Z => mult_21_C241_n898);
   mult_21_C241_U1131 : MUXB2DL port map( A0 => N3096, A1 => N3097, SL => N2913
                           , Z => mult_21_C241_n899);
   mult_21_C241_U1130 : MUXB2DL port map( A0 => N3095, A1 => N3096, SL => N2913
                           , Z => mult_21_C241_n900);
   mult_21_C241_U1129 : MUXB2DL port map( A0 => N3094, A1 => N3095, SL => N2913
                           , Z => mult_21_C241_n901);
   mult_21_C241_U1128 : MUXB2DL port map( A0 => N3093, A1 => N3094, SL => N2913
                           , Z => mult_21_C241_n902);
   mult_21_C241_U1127 : MUXB2DL port map( A0 => N3092, A1 => N3093, SL => N2913
                           , Z => mult_21_C241_n903);
   mult_21_C241_U1126 : MUXB2DL port map( A0 => N3091, A1 => N3092, SL => N2913
                           , Z => mult_21_C241_n904);
   mult_21_C241_U1125 : MUXB2DL port map( A0 => N3090, A1 => N3091, SL => N2913
                           , Z => mult_21_C241_n905);
   mult_21_C241_U1124 : MUXB2DL port map( A0 => N3089, A1 => N3090, SL => N2913
                           , Z => mult_21_C241_n906);
   mult_21_C241_U1123 : MUXB2DL port map( A0 => N3088, A1 => N3089, SL => N2913
                           , Z => mult_21_C241_n907);
   mult_21_C241_U1122 : MUXB2DL port map( A0 => N3087, A1 => N3088, SL => N2913
                           , Z => mult_21_C241_n908);
   mult_21_C241_U1121 : MUXB2DL port map( A0 => N3086, A1 => N3087, SL => N2913
                           , Z => mult_21_C241_n909);
   mult_21_C241_U1120 : AOI21D1 port map( A1 => N2936, A2 => N2937, B => 
                           mult_21_C241_n1417, Z => mult_21_C241_n942);
   mult_21_C241_U1119 : MUXB2DL port map( A0 => N3085, A1 => N3086, SL => 
                           mult_21_C241_n1390, Z => mult_21_C241_n910);
   mult_21_C241_U1118 : MUXB2DL port map( A0 => N3084, A1 => N3085, SL => 
                           mult_21_C241_n1390, Z => mult_21_C241_n911);
   mult_21_C241_U1117 : MUXB2DL port map( A0 => N3083, A1 => N3084, SL => 
                           mult_21_C241_n1390, Z => mult_21_C241_n912);
   mult_21_C241_U1116 : MUXB2DL port map( A0 => N3082, A1 => N3083, SL => 
                           mult_21_C241_n1390, Z => mult_21_C241_n913);
   mult_21_C241_U1115 : MUXB2DL port map( A0 => N3081, A1 => N3082, SL => 
                           mult_21_C241_n1390, Z => mult_21_C241_n914);
   mult_21_C241_U1114 : MUXB2DL port map( A0 => N3080, A1 => N3081, SL => 
                           mult_21_C241_n1390, Z => mult_21_C241_n915);
   mult_21_C241_U1113 : MUXB2DL port map( A0 => N3079, A1 => N3080, SL => 
                           mult_21_C241_n1390, Z => mult_21_C241_n916);
   mult_21_C241_U1112 : MUXB2DL port map( A0 => N3078, A1 => N3079, SL => 
                           mult_21_C241_n1390, Z => mult_21_C241_n917);
   mult_21_C241_U1111 : MUXB2DL port map( A0 => N3077, A1 => N3078, SL => 
                           mult_21_C241_n1390, Z => mult_21_C241_n918);
   mult_21_C241_U1110 : MUXB2DL port map( A0 => mult_21_C241_n1386, A1 => N3077
                           , SL => mult_21_C241_n1390, Z => mult_21_C241_n919);
   mult_21_C241_U1109 : MUXB2DL port map( A0 => N3075, A1 => mult_21_C241_n1386
                           , SL => mult_21_C241_n1390, Z => mult_21_C241_n920);
   mult_21_C241_U1108 : MUXB2DL port map( A0 => mult_21_C241_n1388, A1 => N3075
                           , SL => mult_21_C241_n1390, Z => mult_21_C241_n921);
   mult_21_C241_U1107 : MUXB2DL port map( A0 => N3073, A1 => mult_21_C241_n1388
                           , SL => mult_21_C241_n1390, Z => mult_21_C241_n922);
   mult_21_C241_U1106 : NAN2D1 port map( A1 => N3073, A2 => mult_21_C241_n1390,
                           Z => mult_21_C241_n923);
   mult_21_C241_U1105 : OAI21D1 port map( A1 => N2939, A2 => N2938, B => 
                           mult_21_C241_n1418, Z => mult_21_C241_n94);
   mult_21_C241_U1104 : AOI21D1 port map( A1 => N2938, A2 => N2939, B => 
                           mult_21_C241_n1418, Z => mult_21_C241_n941);
   mult_21_C241_U1103 : OAI21D1 port map( A1 => N2941, A2 => N2940, B => 
                           mult_21_C241_n1421, Z => mult_21_C241_n99);
   mult_21_C241_U1102 : EXOR2D1 port map( A1 => mult_21_C241_n230, A2 => 
                           mult_21_C241_n228, Z => mult_21_C241_n1440);
   mult_21_C241_U1101 : EXOR3D1 port map( A1 => mult_21_C241_n226, A2 => 
                           mult_21_C241_n224, A3 => mult_21_C241_n1440, Z => 
                           mult_21_C241_n1435);
   mult_21_C241_U1100 : EXOR2D1 port map( A1 => mult_21_C241_n222, A2 => 
                           mult_21_C241_n220, Z => mult_21_C241_n1439);
   mult_21_C241_U1099 : EXOR3D1 port map( A1 => mult_21_C241_n216, A2 => 
                           mult_21_C241_n1195, A3 => mult_21_C241_n1439, Z => 
                           mult_21_C241_n1436);
   mult_21_C241_U1098 : EXOR3D1 port map( A1 => mult_21_C241_n1165, A2 => 
                           mult_21_C241_n1137, A3 => mult_21_C241_n1045, Z => 
                           mult_21_C241_n1438);
   mult_21_C241_U1097 : EXOR3D1 port map( A1 => mult_21_C241_n1027, A2 => 
                           mult_21_C241_n1011, A3 => mult_21_C241_n1438, Z => 
                           mult_21_C241_n1437);
   mult_21_C241_U1096 : EXOR3D1 port map( A1 => mult_21_C241_n1435, A2 => 
                           mult_21_C241_n1436, A3 => mult_21_C241_n1437, Z => 
                           mult_21_C241_n1427);
   mult_21_C241_U1095 : EXOR2D1 port map( A1 => mult_21_C241_n985, A2 => 
                           mult_21_C241_n967, Z => mult_21_C241_n1434);
   mult_21_C241_U1094 : EXOR3D1 port map( A1 => mult_21_C241_n961, A2 => 
                           mult_21_C241_n218, A3 => mult_21_C241_n1434, Z => 
                           mult_21_C241_n1431);
   mult_21_C241_U1093 : EXNOR2D1 port map( A1 => mult_21_C241_n210, A2 => 
                           mult_21_C241_n1111, Z => mult_21_C241_n1433);
   mult_21_C241_U1092 : EXOR3D1 port map( A1 => mult_21_C241_n1087, A2 => 
                           mult_21_C241_n1065, A3 => mult_21_C241_n1433, Z => 
                           mult_21_C241_n1432);
   mult_21_C241_U1091 : EXOR3D1 port map( A1 => mult_21_C241_n1431, A2 => 
                           mult_21_C241_n204, A3 => mult_21_C241_n1432, Z => 
                           mult_21_C241_n1428);
   mult_21_C241_U1090 : EXNOR2D1 port map( A1 => mult_21_C241_n997, A2 => 
                           mult_21_C241_n975, Z => mult_21_C241_n1430);
   mult_21_C241_U1089 : EXOR3D1 port map( A1 => mult_21_C241_n957, A2 => 
                           mult_21_C241_n955, A3 => mult_21_C241_n1430, Z => 
                           mult_21_C241_n1429);
   mult_21_C241_U1088 : EXOR3D1 port map( A1 => mult_21_C241_n1427, A2 => 
                           mult_21_C241_n1428, A3 => mult_21_C241_n1429, Z => 
                           mult_21_C241_n1423);
   mult_21_C241_U1087 : EXOR2D1 port map( A1 => mult_21_C241_n202, A2 => 
                           mult_21_C241_n156, Z => mult_21_C241_n1424);
   mult_21_C241_U1086 : EXOR2D1 port map( A1 => mult_21_C241_n214, A2 => 
                           mult_21_C241_n212, Z => mult_21_C241_n1426);
   mult_21_C241_U1085 : EXOR3D1 port map( A1 => mult_21_C241_n208, A2 => 
                           mult_21_C241_n206, A3 => mult_21_C241_n1426, Z => 
                           mult_21_C241_n1425);
   mult_21_C241_U1084 : EXOR3D1 port map( A1 => mult_21_C241_n1423, A2 => 
                           mult_21_C241_n1424, A3 => mult_21_C241_n1425, Z => 
                           N3264);
   mult_21_C241_U1083 : INVD1 port map( A => N2944, Z => mult_21_C241_n1422);
   mult_21_C241_U1082 : INVD1 port map( A => N3076, Z => mult_21_C241_n1387);
   mult_21_C241_U1081 : INVD1 port map( A => N3074, Z => mult_21_C241_n1389);
   mult_21_C241_U1080 : INVD1 port map( A => N2913, Z => mult_21_C241_n1391);
   mult_21_C241_U1079 : MUXB2DL port map( A0 => N3102, A1 => N3101, SL => 
                           mult_21_C241_n1382, Z => mult_21_C241_n862);
   mult_21_C241_U1078 : INVD1 port map( A => N2942, Z => mult_21_C241_n1421);
   mult_21_C241_U1077 : INVD1 port map( A => N2940, Z => mult_21_C241_n1418);
   mult_21_C241_U1076 : INVD1 port map( A => N2938, Z => mult_21_C241_n1417);
   mult_21_C241_U1075 : OAI21D1 port map( A1 => N2935, A2 => N2934, B => 
                           mult_21_C241_n1415, Z => mult_21_C241_n84);
   mult_21_C241_U1074 : INVD1 port map( A => N2936, Z => mult_21_C241_n1415);
   mult_21_C241_U1073 : EXOR2D1 port map( A1 => N2935, A2 => N2934, Z => 
                           mult_21_C241_n1447);
   mult_21_C241_U1072 : OAI21D1 port map( A1 => N2933, A2 => N2932, B => 
                           mult_21_C241_n1413, Z => mult_21_C241_n80);
   mult_21_C241_U1071 : INVD1 port map( A => N2934, Z => mult_21_C241_n1413);
   mult_21_C241_U1070 : EXOR2D1 port map( A1 => N2933, A2 => N2932, Z => 
                           mult_21_C241_n1446);
   mult_21_C241_U1069 : OAI21D1 port map( A1 => N2931, A2 => N2930, B => 
                           mult_21_C241_n1411, Z => mult_21_C241_n73);
   mult_21_C241_U1068 : INVD1 port map( A => N2932, Z => mult_21_C241_n1411);
   mult_21_C241_U1067 : EXOR2D1 port map( A1 => N2931, A2 => N2930, Z => 
                           mult_21_C241_n1445);
   mult_21_C241_U1066 : OAI21D1 port map( A1 => N2929, A2 => N2928, B => 
                           mult_21_C241_n1409, Z => mult_21_C241_n66);
   mult_21_C241_U1065 : INVD1 port map( A => N2930, Z => mult_21_C241_n1409);
   mult_21_C241_U1064 : EXOR2D1 port map( A1 => N2929, A2 => N2928, Z => 
                           mult_21_C241_n1444);
   mult_21_C241_U1063 : OAI21D1 port map( A1 => N2927, A2 => N2926, B => 
                           mult_21_C241_n1407, Z => mult_21_C241_n58);
   mult_21_C241_U1062 : INVD1 port map( A => N2928, Z => mult_21_C241_n1407);
   mult_21_C241_U1061 : EXOR2D1 port map( A1 => N2927, A2 => N2926, Z => 
                           mult_21_C241_n1443);
   mult_21_C241_U1060 : OAI21D1 port map( A1 => N2925, A2 => N2924, B => 
                           mult_21_C241_n1405, Z => mult_21_C241_n50);
   mult_21_C241_U1059 : INVD1 port map( A => N2926, Z => mult_21_C241_n1405);
   mult_21_C241_U1058 : EXOR2D1 port map( A1 => N2925, A2 => N2924, Z => 
                           mult_21_C241_n1442);
   mult_21_C241_U1057 : OAI21D1 port map( A1 => N2922, A2 => N2923, B => 
                           mult_21_C241_n1403, Z => mult_21_C241_n42);
   mult_21_C241_U1056 : INVD1 port map( A => N2924, Z => mult_21_C241_n1403);
   mult_21_C241_U1055 : EXOR2D1 port map( A1 => N2923, A2 => N2922, Z => 
                           mult_21_C241_n1441);
   mult_21_C241_U1054 : INVD1 port map( A => N2922, Z => mult_21_C241_n1401);
   mult_21_C241_U1053 : INVD1 port map( A => N2920, Z => mult_21_C241_n1399);
   mult_21_C241_U1052 : INVD1 port map( A => N2918, Z => mult_21_C241_n1397);
   mult_21_C241_U1051 : INVD1 port map( A => N2916, Z => mult_21_C241_n1395);
   mult_21_C241_U1050 : INVD1 port map( A => mult_21_C241_n1387, Z => 
                           mult_21_C241_n1386);
   mult_21_C241_U1049 : EXNOR2D1 port map( A1 => N2917, A2 => N2916, Z => 
                           mult_21_C241_n1383);
   mult_21_C241_U1048 : INVD1 port map( A => mult_21_C241_n1389, Z => 
                           mult_21_C241_n1388);
   mult_21_C241_U1047 : EXNOR2D1 port map( A1 => N2915, A2 => N2914, Z => 
                           mult_21_C241_n1382);
   mult_21_C241_U1046 : INVD1 port map( A => N2914, Z => mult_21_C241_n1392);
   mult_21_C241_U1045 : INVD1 port map( A => mult_21_C241_n1391, Z => 
                           mult_21_C241_n1390);
   mult_21_C241_U1044 : INVD1 port map( A => mult_21_C241_n939, Z => 
                           mult_21_C241_n1420);
   mult_21_C241_U1043 : INVD1 port map( A => mult_21_C241_n940, Z => 
                           mult_21_C241_n1419);
   mult_21_C241_U1042 : INVD1 port map( A => mult_21_C241_n941, Z => 
                           mult_21_C241_n1416);
   mult_21_C241_U1041 : INVD1 port map( A => mult_21_C241_n942, Z => 
                           mult_21_C241_n1414);
   mult_21_C241_U1040 : INVD1 port map( A => mult_21_C241_n943, Z => 
                           mult_21_C241_n1412);
   mult_21_C241_U1039 : INVD1 port map( A => mult_21_C241_n944, Z => 
                           mult_21_C241_n1410);
   mult_21_C241_U1038 : INVD1 port map( A => mult_21_C241_n945, Z => 
                           mult_21_C241_n1408);
   mult_21_C241_U1037 : INVD1 port map( A => mult_21_C241_n946, Z => 
                           mult_21_C241_n1406);
   mult_21_C241_U1036 : INVD1 port map( A => mult_21_C241_n947, Z => 
                           mult_21_C241_n1404);
   mult_21_C241_U1035 : INVD1 port map( A => mult_21_C241_n948, Z => 
                           mult_21_C241_n1402);
   mult_21_C241_U1034 : INVD1 port map( A => mult_21_C241_n949, Z => 
                           mult_21_C241_n1400);
   mult_21_C241_U1033 : INVD1 port map( A => mult_21_C241_n950, Z => 
                           mult_21_C241_n1398);
   mult_21_C241_U1032 : INVD1 port map( A => mult_21_C241_n951, Z => 
                           mult_21_C241_n1396);
   mult_21_C241_U1031 : INVD1 port map( A => mult_21_C241_n952, Z => 
                           mult_21_C241_n1394);
   mult_21_C241_U1030 : INVD1 port map( A => mult_21_C241_n953, Z => 
                           mult_21_C241_n1393);
   mult_21_C241_U1029 : INVD1 port map( A => mult_21_C241_n1383, Z => 
                           mult_21_C241_n1385);
   mult_21_C241_U1028 : INVD1 port map( A => mult_21_C241_n1382, Z => 
                           mult_21_C241_n1384);
   mult_21_C241_U1027 : OAI21D1 port map( A1 => N2921, A2 => N2920, B => 
                           mult_21_C241_n1401, Z => mult_21_C241_n1381);
   mult_21_C241_U1026 : OAI21D1 port map( A1 => N2919, A2 => N2918, B => 
                           mult_21_C241_n1399, Z => mult_21_C241_n1380);
   mult_21_C241_U1025 : EXOR2D1 port map( A1 => N2921, A2 => N2920, Z => 
                           mult_21_C241_n1379);
   mult_21_C241_U1024 : EXOR2D1 port map( A1 => N2919, A2 => N2918, Z => 
                           mult_21_C241_n1378);
   mult_21_C241_U1023 : OAI21D1 port map( A1 => N2917, A2 => N2916, B => 
                           mult_21_C241_n1397, Z => mult_21_C241_n1377);
   mult_21_C241_U1022 : OAI21D1 port map( A1 => N2915, A2 => N2914, B => 
                           mult_21_C241_n1395, Z => mult_21_C241_n1376);
   mult_21_C241_U1021 : NAN2D1 port map( A1 => mult_21_C241_n1390, A2 => 
                           mult_21_C241_n1392, Z => mult_21_C241_n1375);
   mult_21_C241_U954 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n923, Z => 
                           mult_21_C241_n1226);
   mult_21_C241_U952 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n922, Z => 
                           mult_21_C241_n1225);
   mult_21_C241_U950 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n921, Z => 
                           mult_21_C241_n1224);
   mult_21_C241_U948 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n920, Z => 
                           mult_21_C241_n1223);
   mult_21_C241_U946 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n919, Z => 
                           mult_21_C241_n1222);
   mult_21_C241_U944 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n918, Z => 
                           mult_21_C241_n1221);
   mult_21_C241_U942 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n917, Z => 
                           mult_21_C241_n1220);
   mult_21_C241_U940 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n916, Z => 
                           mult_21_C241_n1219);
   mult_21_C241_U938 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n915, Z => 
                           mult_21_C241_n1218);
   mult_21_C241_U936 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n914, Z => 
                           mult_21_C241_n1217);
   mult_21_C241_U934 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n913, Z => 
                           mult_21_C241_n1216);
   mult_21_C241_U932 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n912, Z => 
                           mult_21_C241_n1215);
   mult_21_C241_U930 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n911, Z => 
                           mult_21_C241_n1214);
   mult_21_C241_U928 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n910, Z => 
                           mult_21_C241_n1213);
   mult_21_C241_U926 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n909, Z => 
                           mult_21_C241_n1212);
   mult_21_C241_U924 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n908, Z => 
                           mult_21_C241_n1211);
   mult_21_C241_U922 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n907, Z => 
                           mult_21_C241_n1210);
   mult_21_C241_U920 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n906, Z => 
                           mult_21_C241_n1209);
   mult_21_C241_U918 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n905, Z => 
                           mult_21_C241_n1208);
   mult_21_C241_U916 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n904, Z => 
                           mult_21_C241_n1207);
   mult_21_C241_U914 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n903, Z => 
                           mult_21_C241_n1206);
   mult_21_C241_U912 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n902, Z => 
                           mult_21_C241_n1205);
   mult_21_C241_U910 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n901, Z => 
                           mult_21_C241_n1204);
   mult_21_C241_U908 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n900, Z => 
                           mult_21_C241_n1203);
   mult_21_C241_U906 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n899, Z => 
                           mult_21_C241_n1202);
   mult_21_C241_U904 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n898, Z => 
                           mult_21_C241_n1201);
   mult_21_C241_U902 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n897, Z => 
                           mult_21_C241_n1200);
   mult_21_C241_U900 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n896, Z => 
                           mult_21_C241_n1199);
   mult_21_C241_U898 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n895, Z => 
                           mult_21_C241_n1198);
   mult_21_C241_U896 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n894, Z => 
                           mult_21_C241_n1197);
   mult_21_C241_U894 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n893, Z => 
                           mult_21_C241_n1196);
   mult_21_C241_U892 : MUXB2DL port map( A0 => mult_21_C241_n1375, A1 => 
                           mult_21_C241_n1392, SL => mult_21_C241_n892, Z => 
                           mult_21_C241_n1195);
   mult_21_C241_U889 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n891, Z => 
                           mult_21_C241_n1194);
   mult_21_C241_U887 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n890, Z => 
                           mult_21_C241_n1193);
   mult_21_C241_U885 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n889, Z => 
                           mult_21_C241_n1192);
   mult_21_C241_U883 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n888, Z => 
                           mult_21_C241_n1191);
   mult_21_C241_U881 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n887, Z => 
                           mult_21_C241_n1190);
   mult_21_C241_U879 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n886, Z => 
                           mult_21_C241_n1189);
   mult_21_C241_U877 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n885, Z => 
                           mult_21_C241_n1188);
   mult_21_C241_U875 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n884, Z => 
                           mult_21_C241_n1187);
   mult_21_C241_U873 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n883, Z => 
                           mult_21_C241_n1186);
   mult_21_C241_U871 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n882, Z => 
                           mult_21_C241_n1185);
   mult_21_C241_U869 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n881, Z => 
                           mult_21_C241_n1184);
   mult_21_C241_U867 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n880, Z => 
                           mult_21_C241_n1183);
   mult_21_C241_U865 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n879, Z => 
                           mult_21_C241_n1182);
   mult_21_C241_U863 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n878, Z => 
                           mult_21_C241_n1181);
   mult_21_C241_U861 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n877, Z => 
                           mult_21_C241_n1180);
   mult_21_C241_U859 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n876, Z => 
                           mult_21_C241_n1179);
   mult_21_C241_U857 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n875, Z => 
                           mult_21_C241_n1178);
   mult_21_C241_U855 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n874, Z => 
                           mult_21_C241_n1177);
   mult_21_C241_U853 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n873, Z => 
                           mult_21_C241_n1176);
   mult_21_C241_U851 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n872, Z => 
                           mult_21_C241_n1175);
   mult_21_C241_U849 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n871, Z => 
                           mult_21_C241_n1174);
   mult_21_C241_U847 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n870, Z => 
                           mult_21_C241_n1173);
   mult_21_C241_U845 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n869, Z => 
                           mult_21_C241_n1172);
   mult_21_C241_U843 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n868, Z => 
                           mult_21_C241_n1171);
   mult_21_C241_U841 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n867, Z => 
                           mult_21_C241_n1170);
   mult_21_C241_U839 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n866, Z => 
                           mult_21_C241_n1169);
   mult_21_C241_U837 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n865, Z => 
                           mult_21_C241_n1168);
   mult_21_C241_U835 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n864, Z => 
                           mult_21_C241_n1167);
   mult_21_C241_U833 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n863, Z => 
                           mult_21_C241_n1166);
   mult_21_C241_U831 : MUXB2DL port map( A0 => mult_21_C241_n1376, A1 => 
                           mult_21_C241_n1393, SL => mult_21_C241_n862, Z => 
                           mult_21_C241_n1165);
   mult_21_C241_U828 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n861, Z => 
                           mult_21_C241_n1164);
   mult_21_C241_U826 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n860, Z => 
                           mult_21_C241_n1163);
   mult_21_C241_U824 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n859, Z => 
                           mult_21_C241_n1162);
   mult_21_C241_U822 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n858, Z => 
                           mult_21_C241_n1161);
   mult_21_C241_U820 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n857, Z => 
                           mult_21_C241_n1160);
   mult_21_C241_U818 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n856, Z => 
                           mult_21_C241_n1159);
   mult_21_C241_U816 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n855, Z => 
                           mult_21_C241_n1158);
   mult_21_C241_U814 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n854, Z => 
                           mult_21_C241_n1157);
   mult_21_C241_U812 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n853, Z => 
                           mult_21_C241_n1156);
   mult_21_C241_U810 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n852, Z => 
                           mult_21_C241_n1155);
   mult_21_C241_U808 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n851, Z => 
                           mult_21_C241_n1154);
   mult_21_C241_U806 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n850, Z => 
                           mult_21_C241_n1153);
   mult_21_C241_U804 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n849, Z => 
                           mult_21_C241_n1152);
   mult_21_C241_U802 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n848, Z => 
                           mult_21_C241_n1151);
   mult_21_C241_U800 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n847, Z => 
                           mult_21_C241_n1150);
   mult_21_C241_U798 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n846, Z => 
                           mult_21_C241_n1149);
   mult_21_C241_U796 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n845, Z => 
                           mult_21_C241_n1148);
   mult_21_C241_U794 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n844, Z => 
                           mult_21_C241_n1147);
   mult_21_C241_U792 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n843, Z => 
                           mult_21_C241_n1146);
   mult_21_C241_U790 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n842, Z => 
                           mult_21_C241_n1145);
   mult_21_C241_U788 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n841, Z => 
                           mult_21_C241_n1144);
   mult_21_C241_U786 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n840, Z => 
                           mult_21_C241_n1143);
   mult_21_C241_U784 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n839, Z => 
                           mult_21_C241_n1142);
   mult_21_C241_U782 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n838, Z => 
                           mult_21_C241_n1141);
   mult_21_C241_U780 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n837, Z => 
                           mult_21_C241_n1140);
   mult_21_C241_U778 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n836, Z => 
                           mult_21_C241_n1139);
   mult_21_C241_U776 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n835, Z => 
                           mult_21_C241_n1138);
   mult_21_C241_U774 : MUXB2DL port map( A0 => mult_21_C241_n1377, A1 => 
                           mult_21_C241_n1394, SL => mult_21_C241_n834, Z => 
                           mult_21_C241_n1137);
   mult_21_C241_U771 : MUXB2DL port map( A0 => mult_21_C241_n1380, A1 => 
                           mult_21_C241_n1396, SL => mult_21_C241_n833, Z => 
                           mult_21_C241_n1136);
   mult_21_C241_U769 : MUXB2DL port map( A0 => mult_21_C241_n1380, A1 => 
                           mult_21_C241_n1396, SL => mult_21_C241_n832, Z => 
                           mult_21_C241_n1135);
   mult_21_C241_U767 : MUXB2DL port map( A0 => mult_21_C241_n1380, A1 => 
                           mult_21_C241_n1396, SL => mult_21_C241_n831, Z => 
                           mult_21_C241_n1134);
   mult_21_C241_U765 : MUXB2DL port map( A0 => mult_21_C241_n1380, A1 => 
                           mult_21_C241_n1396, SL => mult_21_C241_n830, Z => 
                           mult_21_C241_n1133);
   mult_21_C241_U763 : MUXB2DL port map( A0 => mult_21_C241_n1380, A1 => 
                           mult_21_C241_n1396, SL => mult_21_C241_n829, Z => 
                           mult_21_C241_n1132);
   mult_21_C241_U761 : MUXB2DL port map( A0 => mult_21_C241_n1380, A1 => 
                           mult_21_C241_n1396, SL => mult_21_C241_n828, Z => 
                           mult_21_C241_n1131);
   mult_21_C241_U759 : MUXB2DL port map( A0 => mult_21_C241_n1380, A1 => 
                           mult_21_C241_n1396, SL => mult_21_C241_n827, Z => 
                           mult_21_C241_n1130);
   mult_21_C241_U757 : MUXB2DL port map( A0 => mult_21_C241_n1380, A1 => 
                           mult_21_C241_n1396, SL => mult_21_C241_n826, Z => 
                           mult_21_C241_n1129);
   mult_21_C241_U755 : MUXB2DL port map( A0 => mult_21_C241_n1380, A1 => 
                           mult_21_C241_n1396, SL => mult_21_C241_n825, Z => 
                           mult_21_C241_n1128);
   mult_21_C241_U753 : MUXB2DL port map( A0 => mult_21_C241_n1380, A1 => 
                           mult_21_C241_n1396, SL => mult_21_C241_n824, Z => 
                           mult_21_C241_n1127);
   mult_21_C241_U751 : MUXB2DL port map( A0 => mult_21_C241_n1380, A1 => 
                           mult_21_C241_n1396, SL => mult_21_C241_n823, Z => 
                           mult_21_C241_n1126);
   mult_21_C241_U749 : MUXB2DL port map( A0 => mult_21_C241_n1380, A1 => 
                           mult_21_C241_n1396, SL => mult_21_C241_n822, Z => 
                           mult_21_C241_n1125);
   mult_21_C241_U747 : MUXB2DL port map( A0 => mult_21_C241_n1380, A1 => 
                           mult_21_C241_n1396, SL => mult_21_C241_n821, Z => 
                           mult_21_C241_n1124);
   mult_21_C241_U745 : MUXB2DL port map( A0 => mult_21_C241_n1380, A1 => 
                           mult_21_C241_n1396, SL => mult_21_C241_n820, Z => 
                           mult_21_C241_n1123);
   mult_21_C241_U743 : MUXB2DL port map( A0 => mult_21_C241_n1380, A1 => 
                           mult_21_C241_n1396, SL => mult_21_C241_n819, Z => 
                           mult_21_C241_n1122);
   mult_21_C241_U741 : MUXB2DL port map( A0 => mult_21_C241_n1380, A1 => 
                           mult_21_C241_n1396, SL => mult_21_C241_n818, Z => 
                           mult_21_C241_n1121);
   mult_21_C241_U739 : MUXB2DL port map( A0 => mult_21_C241_n1380, A1 => 
                           mult_21_C241_n1396, SL => mult_21_C241_n817, Z => 
                           mult_21_C241_n1120);
   mult_21_C241_U737 : MUXB2DL port map( A0 => mult_21_C241_n1380, A1 => 
                           mult_21_C241_n1396, SL => mult_21_C241_n816, Z => 
                           mult_21_C241_n1119);
   mult_21_C241_U735 : MUXB2DL port map( A0 => mult_21_C241_n1380, A1 => 
                           mult_21_C241_n1396, SL => mult_21_C241_n815, Z => 
                           mult_21_C241_n1118);
   mult_21_C241_U733 : MUXB2DL port map( A0 => mult_21_C241_n1380, A1 => 
                           mult_21_C241_n1396, SL => mult_21_C241_n814, Z => 
                           mult_21_C241_n1117);
   mult_21_C241_U731 : MUXB2DL port map( A0 => mult_21_C241_n1380, A1 => 
                           mult_21_C241_n1396, SL => mult_21_C241_n813, Z => 
                           mult_21_C241_n1116);
   mult_21_C241_U729 : MUXB2DL port map( A0 => mult_21_C241_n1380, A1 => 
                           mult_21_C241_n1396, SL => mult_21_C241_n812, Z => 
                           mult_21_C241_n1115);
   mult_21_C241_U727 : MUXB2DL port map( A0 => mult_21_C241_n1380, A1 => 
                           mult_21_C241_n1396, SL => mult_21_C241_n811, Z => 
                           mult_21_C241_n1114);
   mult_21_C241_U725 : MUXB2DL port map( A0 => mult_21_C241_n1380, A1 => 
                           mult_21_C241_n1396, SL => mult_21_C241_n810, Z => 
                           mult_21_C241_n1113);
   mult_21_C241_U723 : MUXB2DL port map( A0 => mult_21_C241_n1380, A1 => 
                           mult_21_C241_n1396, SL => mult_21_C241_n809, Z => 
                           mult_21_C241_n1112);
   mult_21_C241_U721 : MUXB2DL port map( A0 => mult_21_C241_n1380, A1 => 
                           mult_21_C241_n1396, SL => mult_21_C241_n808, Z => 
                           mult_21_C241_n1111);
   mult_21_C241_U718 : MUXB2DL port map( A0 => mult_21_C241_n1381, A1 => 
                           mult_21_C241_n1398, SL => mult_21_C241_n807, Z => 
                           mult_21_C241_n1110);
   mult_21_C241_U716 : MUXB2DL port map( A0 => mult_21_C241_n1381, A1 => 
                           mult_21_C241_n1398, SL => mult_21_C241_n806, Z => 
                           mult_21_C241_n1109);
   mult_21_C241_U714 : MUXB2DL port map( A0 => mult_21_C241_n1381, A1 => 
                           mult_21_C241_n1398, SL => mult_21_C241_n805, Z => 
                           mult_21_C241_n1108);
   mult_21_C241_U712 : MUXB2DL port map( A0 => mult_21_C241_n1381, A1 => 
                           mult_21_C241_n1398, SL => mult_21_C241_n804, Z => 
                           mult_21_C241_n1107);
   mult_21_C241_U710 : MUXB2DL port map( A0 => mult_21_C241_n1381, A1 => 
                           mult_21_C241_n1398, SL => mult_21_C241_n803, Z => 
                           mult_21_C241_n1106);
   mult_21_C241_U708 : MUXB2DL port map( A0 => mult_21_C241_n1381, A1 => 
                           mult_21_C241_n1398, SL => mult_21_C241_n802, Z => 
                           mult_21_C241_n1105);
   mult_21_C241_U706 : MUXB2DL port map( A0 => mult_21_C241_n1381, A1 => 
                           mult_21_C241_n1398, SL => mult_21_C241_n801, Z => 
                           mult_21_C241_n1104);
   mult_21_C241_U704 : MUXB2DL port map( A0 => mult_21_C241_n1381, A1 => 
                           mult_21_C241_n1398, SL => mult_21_C241_n800, Z => 
                           mult_21_C241_n1103);
   mult_21_C241_U702 : MUXB2DL port map( A0 => mult_21_C241_n1381, A1 => 
                           mult_21_C241_n1398, SL => mult_21_C241_n799, Z => 
                           mult_21_C241_n1102);
   mult_21_C241_U700 : MUXB2DL port map( A0 => mult_21_C241_n1381, A1 => 
                           mult_21_C241_n1398, SL => mult_21_C241_n798, Z => 
                           mult_21_C241_n1101);
   mult_21_C241_U698 : MUXB2DL port map( A0 => mult_21_C241_n1381, A1 => 
                           mult_21_C241_n1398, SL => mult_21_C241_n797, Z => 
                           mult_21_C241_n1100);
   mult_21_C241_U696 : MUXB2DL port map( A0 => mult_21_C241_n1381, A1 => 
                           mult_21_C241_n1398, SL => mult_21_C241_n796, Z => 
                           mult_21_C241_n1099);
   mult_21_C241_U694 : MUXB2DL port map( A0 => mult_21_C241_n1381, A1 => 
                           mult_21_C241_n1398, SL => mult_21_C241_n795, Z => 
                           mult_21_C241_n1098);
   mult_21_C241_U692 : MUXB2DL port map( A0 => mult_21_C241_n1381, A1 => 
                           mult_21_C241_n1398, SL => mult_21_C241_n794, Z => 
                           mult_21_C241_n1097);
   mult_21_C241_U690 : MUXB2DL port map( A0 => mult_21_C241_n1381, A1 => 
                           mult_21_C241_n1398, SL => mult_21_C241_n793, Z => 
                           mult_21_C241_n1096);
   mult_21_C241_U688 : MUXB2DL port map( A0 => mult_21_C241_n1381, A1 => 
                           mult_21_C241_n1398, SL => mult_21_C241_n792, Z => 
                           mult_21_C241_n1095);
   mult_21_C241_U686 : MUXB2DL port map( A0 => mult_21_C241_n1381, A1 => 
                           mult_21_C241_n1398, SL => mult_21_C241_n791, Z => 
                           mult_21_C241_n1094);
   mult_21_C241_U684 : MUXB2DL port map( A0 => mult_21_C241_n1381, A1 => 
                           mult_21_C241_n1398, SL => mult_21_C241_n790, Z => 
                           mult_21_C241_n1093);
   mult_21_C241_U682 : MUXB2DL port map( A0 => mult_21_C241_n1381, A1 => 
                           mult_21_C241_n1398, SL => mult_21_C241_n789, Z => 
                           mult_21_C241_n1092);
   mult_21_C241_U680 : MUXB2DL port map( A0 => mult_21_C241_n1381, A1 => 
                           mult_21_C241_n1398, SL => mult_21_C241_n788, Z => 
                           mult_21_C241_n1091);
   mult_21_C241_U678 : MUXB2DL port map( A0 => mult_21_C241_n1381, A1 => 
                           mult_21_C241_n1398, SL => mult_21_C241_n787, Z => 
                           mult_21_C241_n1090);
   mult_21_C241_U676 : MUXB2DL port map( A0 => mult_21_C241_n1381, A1 => 
                           mult_21_C241_n1398, SL => mult_21_C241_n786, Z => 
                           mult_21_C241_n1089);
   mult_21_C241_U674 : MUXB2DL port map( A0 => mult_21_C241_n1381, A1 => 
                           mult_21_C241_n1398, SL => mult_21_C241_n785, Z => 
                           mult_21_C241_n1088);
   mult_21_C241_U672 : MUXB2DL port map( A0 => mult_21_C241_n1381, A1 => 
                           mult_21_C241_n1398, SL => mult_21_C241_n784, Z => 
                           mult_21_C241_n1087);
   mult_21_C241_U669 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n1400, SL => mult_21_C241_n783, Z => 
                           mult_21_C241_n1086);
   mult_21_C241_U667 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n1400, SL => mult_21_C241_n782, Z => 
                           mult_21_C241_n1085);
   mult_21_C241_U665 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n1400, SL => mult_21_C241_n781, Z => 
                           mult_21_C241_n1084);
   mult_21_C241_U663 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n1400, SL => mult_21_C241_n780, Z => 
                           mult_21_C241_n1083);
   mult_21_C241_U661 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n1400, SL => mult_21_C241_n779, Z => 
                           mult_21_C241_n1082);
   mult_21_C241_U659 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n1400, SL => mult_21_C241_n778, Z => 
                           mult_21_C241_n1081);
   mult_21_C241_U657 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n1400, SL => mult_21_C241_n777, Z => 
                           mult_21_C241_n1080);
   mult_21_C241_U655 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n1400, SL => mult_21_C241_n776, Z => 
                           mult_21_C241_n1079);
   mult_21_C241_U653 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n1400, SL => mult_21_C241_n775, Z => 
                           mult_21_C241_n1078);
   mult_21_C241_U651 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n1400, SL => mult_21_C241_n774, Z => 
                           mult_21_C241_n1077);
   mult_21_C241_U649 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n1400, SL => mult_21_C241_n773, Z => 
                           mult_21_C241_n1076);
   mult_21_C241_U647 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n1400, SL => mult_21_C241_n772, Z => 
                           mult_21_C241_n1075);
   mult_21_C241_U645 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n1400, SL => mult_21_C241_n771, Z => 
                           mult_21_C241_n1074);
   mult_21_C241_U643 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n1400, SL => mult_21_C241_n770, Z => 
                           mult_21_C241_n1073);
   mult_21_C241_U641 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n1400, SL => mult_21_C241_n769, Z => 
                           mult_21_C241_n1072);
   mult_21_C241_U639 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n1400, SL => mult_21_C241_n768, Z => 
                           mult_21_C241_n1071);
   mult_21_C241_U637 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n1400, SL => mult_21_C241_n767, Z => 
                           mult_21_C241_n1070);
   mult_21_C241_U635 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n1400, SL => mult_21_C241_n766, Z => 
                           mult_21_C241_n1069);
   mult_21_C241_U633 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n1400, SL => mult_21_C241_n765, Z => 
                           mult_21_C241_n1068);
   mult_21_C241_U631 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n1400, SL => mult_21_C241_n764, Z => 
                           mult_21_C241_n1067);
   mult_21_C241_U629 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n1400, SL => mult_21_C241_n763, Z => 
                           mult_21_C241_n1066);
   mult_21_C241_U627 : MUXB2DL port map( A0 => mult_21_C241_n42, A1 => 
                           mult_21_C241_n1400, SL => mult_21_C241_n762, Z => 
                           mult_21_C241_n1065);
   mult_21_C241_U624 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n1402, SL => mult_21_C241_n761, Z => 
                           mult_21_C241_n1064);
   mult_21_C241_U622 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n1402, SL => mult_21_C241_n760, Z => 
                           mult_21_C241_n1063);
   mult_21_C241_U620 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n1402, SL => mult_21_C241_n759, Z => 
                           mult_21_C241_n1062);
   mult_21_C241_U618 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n1402, SL => mult_21_C241_n758, Z => 
                           mult_21_C241_n1061);
   mult_21_C241_U616 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n1402, SL => mult_21_C241_n757, Z => 
                           mult_21_C241_n1060);
   mult_21_C241_U614 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n1402, SL => mult_21_C241_n756, Z => 
                           mult_21_C241_n1059);
   mult_21_C241_U612 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n1402, SL => mult_21_C241_n755, Z => 
                           mult_21_C241_n1058);
   mult_21_C241_U610 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n1402, SL => mult_21_C241_n754, Z => 
                           mult_21_C241_n1057);
   mult_21_C241_U608 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n1402, SL => mult_21_C241_n753, Z => 
                           mult_21_C241_n1056);
   mult_21_C241_U606 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n1402, SL => mult_21_C241_n752, Z => 
                           mult_21_C241_n1055);
   mult_21_C241_U604 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n1402, SL => mult_21_C241_n751, Z => 
                           mult_21_C241_n1054);
   mult_21_C241_U602 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n1402, SL => mult_21_C241_n750, Z => 
                           mult_21_C241_n1053);
   mult_21_C241_U600 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n1402, SL => mult_21_C241_n749, Z => 
                           mult_21_C241_n1052);
   mult_21_C241_U598 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n1402, SL => mult_21_C241_n748, Z => 
                           mult_21_C241_n1051);
   mult_21_C241_U596 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n1402, SL => mult_21_C241_n747, Z => 
                           mult_21_C241_n1050);
   mult_21_C241_U594 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n1402, SL => mult_21_C241_n746, Z => 
                           mult_21_C241_n1049);
   mult_21_C241_U592 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n1402, SL => mult_21_C241_n745, Z => 
                           mult_21_C241_n1048);
   mult_21_C241_U590 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n1402, SL => mult_21_C241_n744, Z => 
                           mult_21_C241_n1047);
   mult_21_C241_U588 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n1402, SL => mult_21_C241_n743, Z => 
                           mult_21_C241_n1046);
   mult_21_C241_U586 : MUXB2DL port map( A0 => mult_21_C241_n50, A1 => 
                           mult_21_C241_n1402, SL => mult_21_C241_n742, Z => 
                           mult_21_C241_n1045);
   mult_21_C241_U583 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n1404, SL => mult_21_C241_n741, Z => 
                           mult_21_C241_n1044);
   mult_21_C241_U581 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n1404, SL => mult_21_C241_n740, Z => 
                           mult_21_C241_n1043);
   mult_21_C241_U579 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n1404, SL => mult_21_C241_n739, Z => 
                           mult_21_C241_n1042);
   mult_21_C241_U577 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n1404, SL => mult_21_C241_n738, Z => 
                           mult_21_C241_n1041);
   mult_21_C241_U575 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n1404, SL => mult_21_C241_n737, Z => 
                           mult_21_C241_n1040);
   mult_21_C241_U573 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n1404, SL => mult_21_C241_n736, Z => 
                           mult_21_C241_n1039);
   mult_21_C241_U571 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n1404, SL => mult_21_C241_n735, Z => 
                           mult_21_C241_n1038);
   mult_21_C241_U569 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n1404, SL => mult_21_C241_n734, Z => 
                           mult_21_C241_n1037);
   mult_21_C241_U567 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n1404, SL => mult_21_C241_n733, Z => 
                           mult_21_C241_n1036);
   mult_21_C241_U565 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n1404, SL => mult_21_C241_n732, Z => 
                           mult_21_C241_n1035);
   mult_21_C241_U563 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n1404, SL => mult_21_C241_n731, Z => 
                           mult_21_C241_n1034);
   mult_21_C241_U561 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n1404, SL => mult_21_C241_n730, Z => 
                           mult_21_C241_n1033);
   mult_21_C241_U559 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n1404, SL => mult_21_C241_n729, Z => 
                           mult_21_C241_n1032);
   mult_21_C241_U557 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n1404, SL => mult_21_C241_n728, Z => 
                           mult_21_C241_n1031);
   mult_21_C241_U555 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n1404, SL => mult_21_C241_n727, Z => 
                           mult_21_C241_n1030);
   mult_21_C241_U553 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n1404, SL => mult_21_C241_n726, Z => 
                           mult_21_C241_n1029);
   mult_21_C241_U551 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n1404, SL => mult_21_C241_n725, Z => 
                           mult_21_C241_n1028);
   mult_21_C241_U549 : MUXB2DL port map( A0 => mult_21_C241_n58, A1 => 
                           mult_21_C241_n1404, SL => mult_21_C241_n724, Z => 
                           mult_21_C241_n1027);
   mult_21_C241_U546 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n1406, SL => mult_21_C241_n723, Z => 
                           mult_21_C241_n1026);
   mult_21_C241_U544 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n1406, SL => mult_21_C241_n722, Z => 
                           mult_21_C241_n1025);
   mult_21_C241_U542 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n1406, SL => mult_21_C241_n721, Z => 
                           mult_21_C241_n1024);
   mult_21_C241_U540 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n1406, SL => mult_21_C241_n720, Z => 
                           mult_21_C241_n1023);
   mult_21_C241_U538 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n1406, SL => mult_21_C241_n719, Z => 
                           mult_21_C241_n1022);
   mult_21_C241_U536 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n1406, SL => mult_21_C241_n718, Z => 
                           mult_21_C241_n1021);
   mult_21_C241_U534 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n1406, SL => mult_21_C241_n717, Z => 
                           mult_21_C241_n1020);
   mult_21_C241_U532 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n1406, SL => mult_21_C241_n716, Z => 
                           mult_21_C241_n1019);
   mult_21_C241_U530 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n1406, SL => mult_21_C241_n715, Z => 
                           mult_21_C241_n1018);
   mult_21_C241_U528 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n1406, SL => mult_21_C241_n714, Z => 
                           mult_21_C241_n1017);
   mult_21_C241_U526 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n1406, SL => mult_21_C241_n713, Z => 
                           mult_21_C241_n1016);
   mult_21_C241_U524 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n1406, SL => mult_21_C241_n712, Z => 
                           mult_21_C241_n1015);
   mult_21_C241_U522 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n1406, SL => mult_21_C241_n711, Z => 
                           mult_21_C241_n1014);
   mult_21_C241_U520 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n1406, SL => mult_21_C241_n710, Z => 
                           mult_21_C241_n1013);
   mult_21_C241_U518 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n1406, SL => mult_21_C241_n709, Z => 
                           mult_21_C241_n1012);
   mult_21_C241_U516 : MUXB2DL port map( A0 => mult_21_C241_n66, A1 => 
                           mult_21_C241_n1406, SL => mult_21_C241_n708, Z => 
                           mult_21_C241_n1011);
   mult_21_C241_U513 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n1408, SL => mult_21_C241_n707, Z => 
                           mult_21_C241_n1010);
   mult_21_C241_U511 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n1408, SL => mult_21_C241_n706, Z => 
                           mult_21_C241_n1009);
   mult_21_C241_U509 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n1408, SL => mult_21_C241_n705, Z => 
                           mult_21_C241_n1008);
   mult_21_C241_U507 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n1408, SL => mult_21_C241_n704, Z => 
                           mult_21_C241_n1007);
   mult_21_C241_U505 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n1408, SL => mult_21_C241_n703, Z => 
                           mult_21_C241_n1006);
   mult_21_C241_U503 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n1408, SL => mult_21_C241_n702, Z => 
                           mult_21_C241_n1005);
   mult_21_C241_U501 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n1408, SL => mult_21_C241_n701, Z => 
                           mult_21_C241_n1004);
   mult_21_C241_U499 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n1408, SL => mult_21_C241_n700, Z => 
                           mult_21_C241_n1003);
   mult_21_C241_U497 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n1408, SL => mult_21_C241_n699, Z => 
                           mult_21_C241_n1002);
   mult_21_C241_U495 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n1408, SL => mult_21_C241_n698, Z => 
                           mult_21_C241_n1001);
   mult_21_C241_U493 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n1408, SL => mult_21_C241_n697, Z => 
                           mult_21_C241_n1000);
   mult_21_C241_U491 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n1408, SL => mult_21_C241_n696, Z => 
                           mult_21_C241_n999);
   mult_21_C241_U489 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n1408, SL => mult_21_C241_n695, Z => 
                           mult_21_C241_n998);
   mult_21_C241_U487 : MUXB2DL port map( A0 => mult_21_C241_n73, A1 => 
                           mult_21_C241_n1408, SL => mult_21_C241_n694, Z => 
                           mult_21_C241_n997);
   mult_21_C241_U484 : MUXB2DL port map( A0 => mult_21_C241_n80, A1 => 
                           mult_21_C241_n1410, SL => mult_21_C241_n693, Z => 
                           mult_21_C241_n996);
   mult_21_C241_U482 : MUXB2DL port map( A0 => mult_21_C241_n80, A1 => 
                           mult_21_C241_n1410, SL => mult_21_C241_n692, Z => 
                           mult_21_C241_n995);
   mult_21_C241_U480 : MUXB2DL port map( A0 => mult_21_C241_n80, A1 => 
                           mult_21_C241_n1410, SL => mult_21_C241_n691, Z => 
                           mult_21_C241_n994);
   mult_21_C241_U478 : MUXB2DL port map( A0 => mult_21_C241_n80, A1 => 
                           mult_21_C241_n1410, SL => mult_21_C241_n690, Z => 
                           mult_21_C241_n993);
   mult_21_C241_U476 : MUXB2DL port map( A0 => mult_21_C241_n80, A1 => 
                           mult_21_C241_n1410, SL => mult_21_C241_n689, Z => 
                           mult_21_C241_n992);
   mult_21_C241_U474 : MUXB2DL port map( A0 => mult_21_C241_n80, A1 => 
                           mult_21_C241_n1410, SL => mult_21_C241_n688, Z => 
                           mult_21_C241_n991);
   mult_21_C241_U472 : MUXB2DL port map( A0 => mult_21_C241_n80, A1 => 
                           mult_21_C241_n1410, SL => mult_21_C241_n687, Z => 
                           mult_21_C241_n990);
   mult_21_C241_U470 : MUXB2DL port map( A0 => mult_21_C241_n80, A1 => 
                           mult_21_C241_n1410, SL => mult_21_C241_n686, Z => 
                           mult_21_C241_n989);
   mult_21_C241_U468 : MUXB2DL port map( A0 => mult_21_C241_n80, A1 => 
                           mult_21_C241_n1410, SL => mult_21_C241_n685, Z => 
                           mult_21_C241_n988);
   mult_21_C241_U466 : MUXB2DL port map( A0 => mult_21_C241_n80, A1 => 
                           mult_21_C241_n1410, SL => mult_21_C241_n684, Z => 
                           mult_21_C241_n987);
   mult_21_C241_U464 : MUXB2DL port map( A0 => mult_21_C241_n80, A1 => 
                           mult_21_C241_n1410, SL => mult_21_C241_n683, Z => 
                           mult_21_C241_n986);
   mult_21_C241_U462 : MUXB2DL port map( A0 => mult_21_C241_n80, A1 => 
                           mult_21_C241_n1410, SL => mult_21_C241_n682, Z => 
                           mult_21_C241_n985);
   mult_21_C241_U459 : MUXB2DL port map( A0 => mult_21_C241_n84, A1 => 
                           mult_21_C241_n1412, SL => mult_21_C241_n681, Z => 
                           mult_21_C241_n984);
   mult_21_C241_U457 : MUXB2DL port map( A0 => mult_21_C241_n84, A1 => 
                           mult_21_C241_n1412, SL => mult_21_C241_n680, Z => 
                           mult_21_C241_n983);
   mult_21_C241_U455 : MUXB2DL port map( A0 => mult_21_C241_n84, A1 => 
                           mult_21_C241_n1412, SL => mult_21_C241_n679, Z => 
                           mult_21_C241_n982);
   mult_21_C241_U453 : MUXB2DL port map( A0 => mult_21_C241_n84, A1 => 
                           mult_21_C241_n1412, SL => mult_21_C241_n678, Z => 
                           mult_21_C241_n981);
   mult_21_C241_U451 : MUXB2DL port map( A0 => mult_21_C241_n84, A1 => 
                           mult_21_C241_n1412, SL => mult_21_C241_n677, Z => 
                           mult_21_C241_n980);
   mult_21_C241_U449 : MUXB2DL port map( A0 => mult_21_C241_n84, A1 => 
                           mult_21_C241_n1412, SL => mult_21_C241_n676, Z => 
                           mult_21_C241_n979);
   mult_21_C241_U447 : MUXB2DL port map( A0 => mult_21_C241_n84, A1 => 
                           mult_21_C241_n1412, SL => mult_21_C241_n675, Z => 
                           mult_21_C241_n978);
   mult_21_C241_U445 : MUXB2DL port map( A0 => mult_21_C241_n84, A1 => 
                           mult_21_C241_n1412, SL => mult_21_C241_n674, Z => 
                           mult_21_C241_n977);
   mult_21_C241_U443 : MUXB2DL port map( A0 => mult_21_C241_n84, A1 => 
                           mult_21_C241_n1412, SL => mult_21_C241_n673, Z => 
                           mult_21_C241_n976);
   mult_21_C241_U441 : MUXB2DL port map( A0 => mult_21_C241_n84, A1 => 
                           mult_21_C241_n1412, SL => mult_21_C241_n672, Z => 
                           mult_21_C241_n975);
   mult_21_C241_U438 : MUXB2DL port map( A0 => mult_21_C241_n89, A1 => 
                           mult_21_C241_n1414, SL => mult_21_C241_n671, Z => 
                           mult_21_C241_n974);
   mult_21_C241_U436 : MUXB2DL port map( A0 => mult_21_C241_n89, A1 => 
                           mult_21_C241_n1414, SL => mult_21_C241_n670, Z => 
                           mult_21_C241_n973);
   mult_21_C241_U434 : MUXB2DL port map( A0 => mult_21_C241_n89, A1 => 
                           mult_21_C241_n1414, SL => mult_21_C241_n669, Z => 
                           mult_21_C241_n972);
   mult_21_C241_U432 : MUXB2DL port map( A0 => mult_21_C241_n89, A1 => 
                           mult_21_C241_n1414, SL => mult_21_C241_n668, Z => 
                           mult_21_C241_n971);
   mult_21_C241_U430 : MUXB2DL port map( A0 => mult_21_C241_n89, A1 => 
                           mult_21_C241_n1414, SL => mult_21_C241_n667, Z => 
                           mult_21_C241_n970);
   mult_21_C241_U428 : MUXB2DL port map( A0 => mult_21_C241_n89, A1 => 
                           mult_21_C241_n1414, SL => mult_21_C241_n666, Z => 
                           mult_21_C241_n969);
   mult_21_C241_U426 : MUXB2DL port map( A0 => mult_21_C241_n89, A1 => 
                           mult_21_C241_n1414, SL => mult_21_C241_n665, Z => 
                           mult_21_C241_n968);
   mult_21_C241_U424 : MUXB2DL port map( A0 => mult_21_C241_n89, A1 => 
                           mult_21_C241_n1414, SL => mult_21_C241_n664, Z => 
                           mult_21_C241_n967);
   mult_21_C241_U421 : MUXB2DL port map( A0 => mult_21_C241_n94, A1 => 
                           mult_21_C241_n1416, SL => mult_21_C241_n663, Z => 
                           mult_21_C241_n966);
   mult_21_C241_U419 : MUXB2DL port map( A0 => mult_21_C241_n94, A1 => 
                           mult_21_C241_n1416, SL => mult_21_C241_n662, Z => 
                           mult_21_C241_n965);
   mult_21_C241_U417 : MUXB2DL port map( A0 => mult_21_C241_n94, A1 => 
                           mult_21_C241_n1416, SL => mult_21_C241_n661, Z => 
                           mult_21_C241_n964);
   mult_21_C241_U415 : MUXB2DL port map( A0 => mult_21_C241_n94, A1 => 
                           mult_21_C241_n1416, SL => mult_21_C241_n660, Z => 
                           mult_21_C241_n963);
   mult_21_C241_U413 : MUXB2DL port map( A0 => mult_21_C241_n94, A1 => 
                           mult_21_C241_n1416, SL => mult_21_C241_n659, Z => 
                           mult_21_C241_n962);
   mult_21_C241_U411 : MUXB2DL port map( A0 => mult_21_C241_n94, A1 => 
                           mult_21_C241_n1416, SL => mult_21_C241_n658, Z => 
                           mult_21_C241_n961);
   mult_21_C241_U408 : MUXB2DL port map( A0 => mult_21_C241_n99, A1 => 
                           mult_21_C241_n1419, SL => mult_21_C241_n657, Z => 
                           mult_21_C241_n960);
   mult_21_C241_U406 : MUXB2DL port map( A0 => mult_21_C241_n99, A1 => 
                           mult_21_C241_n1419, SL => mult_21_C241_n656, Z => 
                           mult_21_C241_n959);
   mult_21_C241_U404 : MUXB2DL port map( A0 => mult_21_C241_n99, A1 => 
                           mult_21_C241_n1419, SL => mult_21_C241_n655, Z => 
                           mult_21_C241_n958);
   mult_21_C241_U402 : MUXB2DL port map( A0 => mult_21_C241_n99, A1 => 
                           mult_21_C241_n1419, SL => mult_21_C241_n654, Z => 
                           mult_21_C241_n957);
   mult_21_C241_U399 : MUXB2DL port map( A0 => mult_21_C241_n104, A1 => 
                           mult_21_C241_n1420, SL => mult_21_C241_n653, Z => 
                           mult_21_C241_n956);
   mult_21_C241_U397 : MUXB2DL port map( A0 => mult_21_C241_n104, A1 => 
                           mult_21_C241_n1420, SL => mult_21_C241_n652, Z => 
                           mult_21_C241_n955);
   mult_21_C241_U395 : ADHALFDL port map( A => mult_21_C241_n1224, B => 
                           mult_21_C241_n953, CO => mult_21_C241_n650, S => 
                           mult_21_C241_n651);
   mult_21_C241_U394 : ADHALFDL port map( A => mult_21_C241_n650, B => 
                           mult_21_C241_n1223, CO => mult_21_C241_n648, S => 
                           mult_21_C241_n649);
   mult_21_C241_U393 : ADHALFDL port map( A => mult_21_C241_n1222, B => 
                           mult_21_C241_n952, CO => mult_21_C241_n646, S => 
                           mult_21_C241_n647);
   mult_21_C241_U392 : ADFULD1 port map( A => mult_21_C241_n1192, B => 
                           mult_21_C241_n1164, CI => mult_21_C241_n647, CO => 
                           mult_21_C241_n644, S => mult_21_C241_n645);
   mult_21_C241_U391 : ADHALFDL port map( A => mult_21_C241_n646, B => 
                           mult_21_C241_n1221, CO => mult_21_C241_n642, S => 
                           mult_21_C241_n643);
   mult_21_C241_U390 : ADFULD1 port map( A => mult_21_C241_n1163, B => 
                           mult_21_C241_n1191, CI => mult_21_C241_n643, CO => 
                           mult_21_C241_n640, S => mult_21_C241_n641);
   mult_21_C241_U389 : ADHALFDL port map( A => mult_21_C241_n1220, B => 
                           mult_21_C241_n951, CO => mult_21_C241_n638, S => 
                           mult_21_C241_n639);
   mult_21_C241_U388 : ADFULD1 port map( A => mult_21_C241_n1190, B => 
                           mult_21_C241_n1136, CI => mult_21_C241_n1162, CO => 
                           mult_21_C241_n636, S => mult_21_C241_n637);
   mult_21_C241_U387 : ADFULD1 port map( A => mult_21_C241_n642, B => 
                           mult_21_C241_n639, CI => mult_21_C241_n637, CO => 
                           mult_21_C241_n634, S => mult_21_C241_n635);
   mult_21_C241_U386 : ADHALFDL port map( A => mult_21_C241_n638, B => 
                           mult_21_C241_n1219, CO => mult_21_C241_n632, S => 
                           mult_21_C241_n633);
   mult_21_C241_U385 : ADFULD1 port map( A => mult_21_C241_n1135, B => 
                           mult_21_C241_n1189, CI => mult_21_C241_n1161, CO => 
                           mult_21_C241_n630, S => mult_21_C241_n631);
   mult_21_C241_U384 : ADFULD1 port map( A => mult_21_C241_n636, B => 
                           mult_21_C241_n633, CI => mult_21_C241_n631, CO => 
                           mult_21_C241_n628, S => mult_21_C241_n629);
   mult_21_C241_U383 : ADHALFDL port map( A => mult_21_C241_n1218, B => 
                           mult_21_C241_n950, CO => mult_21_C241_n626, S => 
                           mult_21_C241_n627);
   mult_21_C241_U382 : ADFULD1 port map( A => mult_21_C241_n1188, B => 
                           mult_21_C241_n1110, CI => mult_21_C241_n1134, CO => 
                           mult_21_C241_n624, S => mult_21_C241_n625);
   mult_21_C241_U381 : ADFULD1 port map( A => mult_21_C241_n627, B => 
                           mult_21_C241_n1160, CI => mult_21_C241_n632, CO => 
                           mult_21_C241_n622, S => mult_21_C241_n623);
   mult_21_C241_U380 : ADFULD1 port map( A => mult_21_C241_n625, B => 
                           mult_21_C241_n630, CI => mult_21_C241_n623, CO => 
                           mult_21_C241_n620, S => mult_21_C241_n621);
   mult_21_C241_U379 : ADHALFDL port map( A => mult_21_C241_n626, B => 
                           mult_21_C241_n1217, CO => mult_21_C241_n618, S => 
                           mult_21_C241_n619);
   mult_21_C241_U378 : ADFULD1 port map( A => mult_21_C241_n1109, B => 
                           mult_21_C241_n1133, CI => mult_21_C241_n1159, CO => 
                           mult_21_C241_n616, S => mult_21_C241_n617);
   mult_21_C241_U377 : ADFULD1 port map( A => mult_21_C241_n619, B => 
                           mult_21_C241_n1187, CI => mult_21_C241_n624, CO => 
                           mult_21_C241_n614, S => mult_21_C241_n615);
   mult_21_C241_U376 : ADFULD1 port map( A => mult_21_C241_n617, B => 
                           mult_21_C241_n622, CI => mult_21_C241_n615, CO => 
                           mult_21_C241_n612, S => mult_21_C241_n613);
   mult_21_C241_U375 : ADHALFDL port map( A => mult_21_C241_n1216, B => 
                           mult_21_C241_n949, CO => mult_21_C241_n610, S => 
                           mult_21_C241_n611);
   mult_21_C241_U374 : ADFULD1 port map( A => mult_21_C241_n1132, B => 
                           mult_21_C241_n1086, CI => mult_21_C241_n1186, CO => 
                           mult_21_C241_n608, S => mult_21_C241_n609);
   mult_21_C241_U373 : ADFULD1 port map( A => mult_21_C241_n1108, B => 
                           mult_21_C241_n1158, CI => mult_21_C241_n611, CO => 
                           mult_21_C241_n606, S => mult_21_C241_n607);
   mult_21_C241_U372 : ADFULD1 port map( A => mult_21_C241_n616, B => 
                           mult_21_C241_n618, CI => mult_21_C241_n609, CO => 
                           mult_21_C241_n604, S => mult_21_C241_n605);
   mult_21_C241_U371 : ADFULD1 port map( A => mult_21_C241_n614, B => 
                           mult_21_C241_n607, CI => mult_21_C241_n605, CO => 
                           mult_21_C241_n602, S => mult_21_C241_n603);
   mult_21_C241_U370 : ADHALFDL port map( A => mult_21_C241_n610, B => 
                           mult_21_C241_n1215, CO => mult_21_C241_n600, S => 
                           mult_21_C241_n601);
   mult_21_C241_U369 : ADFULD1 port map( A => mult_21_C241_n1085, B => 
                           mult_21_C241_n1131, CI => mult_21_C241_n1185, CO => 
                           mult_21_C241_n598, S => mult_21_C241_n599);
   mult_21_C241_U368 : ADFULD1 port map( A => mult_21_C241_n1107, B => 
                           mult_21_C241_n1157, CI => mult_21_C241_n601, CO => 
                           mult_21_C241_n596, S => mult_21_C241_n597);
   mult_21_C241_U367 : ADFULD1 port map( A => mult_21_C241_n606, B => 
                           mult_21_C241_n608, CI => mult_21_C241_n599, CO => 
                           mult_21_C241_n594, S => mult_21_C241_n595);
   mult_21_C241_U366 : ADFULD1 port map( A => mult_21_C241_n604, B => 
                           mult_21_C241_n597, CI => mult_21_C241_n595, CO => 
                           mult_21_C241_n592, S => mult_21_C241_n593);
   mult_21_C241_U365 : ADHALFDL port map( A => mult_21_C241_n1214, B => 
                           mult_21_C241_n948, CO => mult_21_C241_n590, S => 
                           mult_21_C241_n591);
   mult_21_C241_U364 : ADFULD1 port map( A => mult_21_C241_n1130, B => 
                           mult_21_C241_n1064, CI => mult_21_C241_n1184, CO => 
                           mult_21_C241_n588, S => mult_21_C241_n589);
   mult_21_C241_U363 : ADFULD1 port map( A => mult_21_C241_n1084, B => 
                           mult_21_C241_n1156, CI => mult_21_C241_n591, CO => 
                           mult_21_C241_n586, S => mult_21_C241_n587);
   mult_21_C241_U362 : ADFULD1 port map( A => mult_21_C241_n600, B => 
                           mult_21_C241_n1106, CI => mult_21_C241_n598, CO => 
                           mult_21_C241_n584, S => mult_21_C241_n585);
   mult_21_C241_U361 : ADFULD1 port map( A => mult_21_C241_n587, B => 
                           mult_21_C241_n589, CI => mult_21_C241_n596, CO => 
                           mult_21_C241_n582, S => mult_21_C241_n583);
   mult_21_C241_U360 : ADFULD1 port map( A => mult_21_C241_n585, B => 
                           mult_21_C241_n594, CI => mult_21_C241_n583, CO => 
                           mult_21_C241_n580, S => mult_21_C241_n581);
   mult_21_C241_U359 : ADHALFDL port map( A => mult_21_C241_n590, B => 
                           mult_21_C241_n1213, CO => mult_21_C241_n578, S => 
                           mult_21_C241_n579);
   mult_21_C241_U358 : ADFULD1 port map( A => mult_21_C241_n1183, B => 
                           mult_21_C241_n1105, CI => mult_21_C241_n1155, CO => 
                           mult_21_C241_n576, S => mult_21_C241_n577);
   mult_21_C241_U357 : ADFULD1 port map( A => mult_21_C241_n1063, B => 
                           mult_21_C241_n1129, CI => mult_21_C241_n1083, CO => 
                           mult_21_C241_n574, S => mult_21_C241_n575);
   mult_21_C241_U356 : ADFULD1 port map( A => mult_21_C241_n588, B => 
                           mult_21_C241_n579, CI => mult_21_C241_n586, CO => 
                           mult_21_C241_n572, S => mult_21_C241_n573);
   mult_21_C241_U355 : ADFULD1 port map( A => mult_21_C241_n577, B => 
                           mult_21_C241_n575, CI => mult_21_C241_n584, CO => 
                           mult_21_C241_n570, S => mult_21_C241_n571);
   mult_21_C241_U354 : ADFULD1 port map( A => mult_21_C241_n582, B => 
                           mult_21_C241_n573, CI => mult_21_C241_n571, CO => 
                           mult_21_C241_n568, S => mult_21_C241_n569);
   mult_21_C241_U353 : ADHALFDL port map( A => mult_21_C241_n1212, B => 
                           mult_21_C241_n947, CO => mult_21_C241_n566, S => 
                           mult_21_C241_n567);
   mult_21_C241_U352 : ADFULD1 port map( A => mult_21_C241_n1104, B => 
                           mult_21_C241_n1044, CI => mult_21_C241_n1182, CO => 
                           mult_21_C241_n564, S => mult_21_C241_n565);
   mult_21_C241_U351 : ADFULD1 port map( A => mult_21_C241_n1154, B => 
                           mult_21_C241_n1082, CI => mult_21_C241_n567, CO => 
                           mult_21_C241_n562, S => mult_21_C241_n563);
   mult_21_C241_U350 : ADFULD1 port map( A => mult_21_C241_n1062, B => 
                           mult_21_C241_n1128, CI => mult_21_C241_n578, CO => 
                           mult_21_C241_n560, S => mult_21_C241_n561);
   mult_21_C241_U349 : ADFULD1 port map( A => mult_21_C241_n574, B => 
                           mult_21_C241_n576, CI => mult_21_C241_n565, CO => 
                           mult_21_C241_n558, S => mult_21_C241_n559);
   mult_21_C241_U348 : ADFULD1 port map( A => mult_21_C241_n561, B => 
                           mult_21_C241_n563, CI => mult_21_C241_n572, CO => 
                           mult_21_C241_n556, S => mult_21_C241_n557);
   mult_21_C241_U347 : ADFULD1 port map( A => mult_21_C241_n570, B => 
                           mult_21_C241_n559, CI => mult_21_C241_n557, CO => 
                           mult_21_C241_n554, S => mult_21_C241_n555);
   mult_21_C241_U346 : ADHALFDL port map( A => mult_21_C241_n566, B => 
                           mult_21_C241_n1211, CO => mult_21_C241_n552, S => 
                           mult_21_C241_n553);
   mult_21_C241_U345 : ADFULD1 port map( A => mult_21_C241_n1043, B => 
                           mult_21_C241_n1103, CI => mult_21_C241_n1061, CO => 
                           mult_21_C241_n550, S => mult_21_C241_n551);
   mult_21_C241_U344 : ADFULD1 port map( A => mult_21_C241_n1181, B => 
                           mult_21_C241_n1081, CI => mult_21_C241_n1127, CO => 
                           mult_21_C241_n548, S => mult_21_C241_n549);
   mult_21_C241_U343 : ADFULD1 port map( A => mult_21_C241_n553, B => 
                           mult_21_C241_n1153, CI => mult_21_C241_n564, CO => 
                           mult_21_C241_n546, S => mult_21_C241_n547);
   mult_21_C241_U342 : ADFULD1 port map( A => mult_21_C241_n560, B => 
                           mult_21_C241_n562, CI => mult_21_C241_n549, CO => 
                           mult_21_C241_n544, S => mult_21_C241_n545);
   mult_21_C241_U341 : ADFULD1 port map( A => mult_21_C241_n547, B => 
                           mult_21_C241_n551, CI => mult_21_C241_n558, CO => 
                           mult_21_C241_n542, S => mult_21_C241_n543);
   mult_21_C241_U340 : ADFULD1 port map( A => mult_21_C241_n556, B => 
                           mult_21_C241_n545, CI => mult_21_C241_n543, CO => 
                           mult_21_C241_n540, S => mult_21_C241_n541);
   mult_21_C241_U339 : ADHALFDL port map( A => mult_21_C241_n1210, B => 
                           mult_21_C241_n946, CO => mult_21_C241_n538, S => 
                           mult_21_C241_n539);
   mult_21_C241_U338 : ADFULD1 port map( A => mult_21_C241_n1102, B => 
                           mult_21_C241_n1026, CI => mult_21_C241_n1180, CO => 
                           mult_21_C241_n536, S => mult_21_C241_n537);
   mult_21_C241_U337 : ADFULD1 port map( A => mult_21_C241_n1042, B => 
                           mult_21_C241_n1060, CI => mult_21_C241_n539, CO => 
                           mult_21_C241_n534, S => mult_21_C241_n535);
   mult_21_C241_U336 : ADFULD1 port map( A => mult_21_C241_n1080, B => 
                           mult_21_C241_n1152, CI => mult_21_C241_n1126, CO => 
                           mult_21_C241_n532, S => mult_21_C241_n533);
   mult_21_C241_U335 : ADFULD1 port map( A => mult_21_C241_n550, B => 
                           mult_21_C241_n552, CI => mult_21_C241_n548, CO => 
                           mult_21_C241_n530, S => mult_21_C241_n531);
   mult_21_C241_U334 : ADFULD1 port map( A => mult_21_C241_n533, B => 
                           mult_21_C241_n537, CI => mult_21_C241_n535, CO => 
                           mult_21_C241_n528, S => mult_21_C241_n529);
   mult_21_C241_U333 : ADFULD1 port map( A => mult_21_C241_n544, B => 
                           mult_21_C241_n546, CI => mult_21_C241_n531, CO => 
                           mult_21_C241_n526, S => mult_21_C241_n527);
   mult_21_C241_U332 : ADFULD1 port map( A => mult_21_C241_n542, B => 
                           mult_21_C241_n529, CI => mult_21_C241_n527, CO => 
                           mult_21_C241_n524, S => mult_21_C241_n525);
   mult_21_C241_U331 : ADHALFDL port map( A => mult_21_C241_n538, B => 
                           mult_21_C241_n1209, CO => mult_21_C241_n522, S => 
                           mult_21_C241_n523);
   mult_21_C241_U330 : ADFULD1 port map( A => mult_21_C241_n1179, B => 
                           mult_21_C241_n1079, CI => mult_21_C241_n1151, CO => 
                           mult_21_C241_n520, S => mult_21_C241_n521);
   mult_21_C241_U329 : ADFULD1 port map( A => mult_21_C241_n1025, B => 
                           mult_21_C241_n1041, CI => mult_21_C241_n1059, CO => 
                           mult_21_C241_n518, S => mult_21_C241_n519);
   mult_21_C241_U328 : ADFULD1 port map( A => mult_21_C241_n1101, B => 
                           mult_21_C241_n1125, CI => mult_21_C241_n523, CO => 
                           mult_21_C241_n516, S => mult_21_C241_n517);
   mult_21_C241_U327 : ADFULD1 port map( A => mult_21_C241_n534, B => 
                           mult_21_C241_n536, CI => mult_21_C241_n532, CO => 
                           mult_21_C241_n514, S => mult_21_C241_n515);
   mult_21_C241_U326 : ADFULD1 port map( A => mult_21_C241_n521, B => 
                           mult_21_C241_n519, CI => mult_21_C241_n517, CO => 
                           mult_21_C241_n512, S => mult_21_C241_n513);
   mult_21_C241_U325 : ADFULD1 port map( A => mult_21_C241_n528, B => 
                           mult_21_C241_n530, CI => mult_21_C241_n515, CO => 
                           mult_21_C241_n510, S => mult_21_C241_n511);
   mult_21_C241_U324 : ADFULD1 port map( A => mult_21_C241_n526, B => 
                           mult_21_C241_n513, CI => mult_21_C241_n511, CO => 
                           mult_21_C241_n508, S => mult_21_C241_n509);
   mult_21_C241_U323 : ADHALFDL port map( A => mult_21_C241_n1208, B => 
                           mult_21_C241_n945, CO => mult_21_C241_n506, S => 
                           mult_21_C241_n507);
   mult_21_C241_U322 : ADFULD1 port map( A => mult_21_C241_n1078, B => 
                           mult_21_C241_n1010, CI => mult_21_C241_n1024, CO => 
                           mult_21_C241_n504, S => mult_21_C241_n505);
   mult_21_C241_U321 : ADFULD1 port map( A => mult_21_C241_n1178, B => 
                           mult_21_C241_n1100, CI => mult_21_C241_n507, CO => 
                           mult_21_C241_n502, S => mult_21_C241_n503);
   mult_21_C241_U320 : ADFULD1 port map( A => mult_21_C241_n1040, B => 
                           mult_21_C241_n1150, CI => mult_21_C241_n1058, CO => 
                           mult_21_C241_n500, S => mult_21_C241_n501);
   mult_21_C241_U319 : ADFULD1 port map( A => mult_21_C241_n522, B => 
                           mult_21_C241_n1124, CI => mult_21_C241_n520, CO => 
                           mult_21_C241_n498, S => mult_21_C241_n499);
   mult_21_C241_U318 : ADFULD1 port map( A => mult_21_C241_n505, B => 
                           mult_21_C241_n518, CI => mult_21_C241_n501, CO => 
                           mult_21_C241_n496, S => mult_21_C241_n497);
   mult_21_C241_U317 : ADFULD1 port map( A => mult_21_C241_n516, B => 
                           mult_21_C241_n503, CI => mult_21_C241_n514, CO => 
                           mult_21_C241_n494, S => mult_21_C241_n495);
   mult_21_C241_U316 : ADFULD1 port map( A => mult_21_C241_n497, B => 
                           mult_21_C241_n499, CI => mult_21_C241_n512, CO => 
                           mult_21_C241_n492, S => mult_21_C241_n493);
   mult_21_C241_U315 : ADFULD1 port map( A => mult_21_C241_n510, B => 
                           mult_21_C241_n495, CI => mult_21_C241_n493, CO => 
                           mult_21_C241_n490, S => mult_21_C241_n491);
   mult_21_C241_U314 : ADHALFDL port map( A => mult_21_C241_n506, B => 
                           mult_21_C241_n1207, CO => mult_21_C241_n488, S => 
                           mult_21_C241_n489);
   mult_21_C241_U313 : ADFULD1 port map( A => mult_21_C241_n1009, B => 
                           mult_21_C241_n1077, CI => mult_21_C241_n1023, CO => 
                           mult_21_C241_n486, S => mult_21_C241_n487);
   mult_21_C241_U312 : ADFULD1 port map( A => mult_21_C241_n1177, B => 
                           mult_21_C241_n1099, CI => mult_21_C241_n1039, CO => 
                           mult_21_C241_n484, S => mult_21_C241_n485);
   mult_21_C241_U311 : ADFULD1 port map( A => mult_21_C241_n1057, B => 
                           mult_21_C241_n1149, CI => mult_21_C241_n1123, CO => 
                           mult_21_C241_n482, S => mult_21_C241_n483);
   mult_21_C241_U310 : ADFULD1 port map( A => mult_21_C241_n504, B => 
                           mult_21_C241_n489, CI => mult_21_C241_n502, CO => 
                           mult_21_C241_n480, S => mult_21_C241_n481);
   mult_21_C241_U309 : ADFULD1 port map( A => mult_21_C241_n483, B => 
                           mult_21_C241_n500, CI => mult_21_C241_n485, CO => 
                           mult_21_C241_n478, S => mult_21_C241_n479);
   mult_21_C241_U308 : ADFULD1 port map( A => mult_21_C241_n498, B => 
                           mult_21_C241_n487, CI => mult_21_C241_n496, CO => 
                           mult_21_C241_n476, S => mult_21_C241_n477);
   mult_21_C241_U307 : ADFULD1 port map( A => mult_21_C241_n479, B => 
                           mult_21_C241_n481, CI => mult_21_C241_n494, CO => 
                           mult_21_C241_n474, S => mult_21_C241_n475);
   mult_21_C241_U306 : ADFULD1 port map( A => mult_21_C241_n492, B => 
                           mult_21_C241_n477, CI => mult_21_C241_n475, CO => 
                           mult_21_C241_n472, S => mult_21_C241_n473);
   mult_21_C241_U305 : ADHALFDL port map( A => mult_21_C241_n1206, B => 
                           mult_21_C241_n944, CO => mult_21_C241_n470, S => 
                           mult_21_C241_n471);
   mult_21_C241_U304 : ADFULD1 port map( A => mult_21_C241_n1076, B => 
                           mult_21_C241_n996, CI => mult_21_C241_n1176, CO => 
                           mult_21_C241_n468, S => mult_21_C241_n469);
   mult_21_C241_U303 : ADFULD1 port map( A => mult_21_C241_n1008, B => 
                           mult_21_C241_n1038, CI => mult_21_C241_n471, CO => 
                           mult_21_C241_n466, S => mult_21_C241_n467);
   mult_21_C241_U302 : ADFULD1 port map( A => mult_21_C241_n1022, B => 
                           mult_21_C241_n1148, CI => mult_21_C241_n1056, CO => 
                           mult_21_C241_n464, S => mult_21_C241_n465);
   mult_21_C241_U301 : ADFULD1 port map( A => mult_21_C241_n1098, B => 
                           mult_21_C241_n1122, CI => mult_21_C241_n488, CO => 
                           mult_21_C241_n462, S => mult_21_C241_n463);
   mult_21_C241_U300 : ADFULD1 port map( A => mult_21_C241_n482, B => 
                           mult_21_C241_n486, CI => mult_21_C241_n484, CO => 
                           mult_21_C241_n460, S => mult_21_C241_n461);
   mult_21_C241_U299 : ADFULD1 port map( A => mult_21_C241_n465, B => 
                           mult_21_C241_n469, CI => mult_21_C241_n467, CO => 
                           mult_21_C241_n458, S => mult_21_C241_n459);
   mult_21_C241_U298 : ADFULD1 port map( A => mult_21_C241_n480, B => 
                           mult_21_C241_n463, CI => mult_21_C241_n478, CO => 
                           mult_21_C241_n456, S => mult_21_C241_n457);
   mult_21_C241_U297 : ADFULD1 port map( A => mult_21_C241_n459, B => 
                           mult_21_C241_n461, CI => mult_21_C241_n476, CO => 
                           mult_21_C241_n454, S => mult_21_C241_n455);
   mult_21_C241_U296 : ADFULD1 port map( A => mult_21_C241_n474, B => 
                           mult_21_C241_n457, CI => mult_21_C241_n455, CO => 
                           mult_21_C241_n452, S => mult_21_C241_n453);
   mult_21_C241_U295 : ADHALFDL port map( A => mult_21_C241_n470, B => 
                           mult_21_C241_n1205, CO => mult_21_C241_n450, S => 
                           mult_21_C241_n451);
   mult_21_C241_U294 : ADFULD1 port map( A => mult_21_C241_n1175, B => 
                           mult_21_C241_n1055, CI => mult_21_C241_n1147, CO => 
                           mult_21_C241_n448, S => mult_21_C241_n449);
   mult_21_C241_U293 : ADFULD1 port map( A => mult_21_C241_n1121, B => 
                           mult_21_C241_n1021, CI => mult_21_C241_n1097, CO => 
                           mult_21_C241_n446, S => mult_21_C241_n447);
   mult_21_C241_U292 : ADFULD1 port map( A => mult_21_C241_n995, B => 
                           mult_21_C241_n1075, CI => mult_21_C241_n1007, CO => 
                           mult_21_C241_n444, S => mult_21_C241_n445);
   mult_21_C241_U291 : ADFULD1 port map( A => mult_21_C241_n451, B => 
                           mult_21_C241_n1037, CI => mult_21_C241_n468, CO => 
                           mult_21_C241_n442, S => mult_21_C241_n443);
   mult_21_C241_U290 : ADFULD1 port map( A => mult_21_C241_n464, B => 
                           mult_21_C241_n466, CI => mult_21_C241_n462, CO => 
                           mult_21_C241_n440, S => mult_21_C241_n441);
   mult_21_C241_U289 : ADFULD1 port map( A => mult_21_C241_n449, B => 
                           mult_21_C241_n445, CI => mult_21_C241_n447, CO => 
                           mult_21_C241_n438, S => mult_21_C241_n439);
   mult_21_C241_U288 : ADFULD1 port map( A => mult_21_C241_n443, B => 
                           mult_21_C241_n460, CI => mult_21_C241_n458, CO => 
                           mult_21_C241_n436, S => mult_21_C241_n437);
   mult_21_C241_U287 : ADFULD1 port map( A => mult_21_C241_n439, B => 
                           mult_21_C241_n441, CI => mult_21_C241_n456, CO => 
                           mult_21_C241_n434, S => mult_21_C241_n435);
   mult_21_C241_U286 : ADFULD1 port map( A => mult_21_C241_n454, B => 
                           mult_21_C241_n437, CI => mult_21_C241_n435, CO => 
                           mult_21_C241_n432, S => mult_21_C241_n433);
   mult_21_C241_U285 : ADHALFDL port map( A => mult_21_C241_n1204, B => 
                           mult_21_C241_n943, CO => mult_21_C241_n430, S => 
                           mult_21_C241_n431);
   mult_21_C241_U284 : ADFULD1 port map( A => mult_21_C241_n1054, B => 
                           mult_21_C241_n984, CI => mult_21_C241_n994, CO => 
                           mult_21_C241_n428, S => mult_21_C241_n429);
   mult_21_C241_U283 : ADFULD1 port map( A => mult_21_C241_n1174, B => 
                           mult_21_C241_n1036, CI => mult_21_C241_n431, CO => 
                           mult_21_C241_n426, S => mult_21_C241_n427);
   mult_21_C241_U282 : ADFULD1 port map( A => mult_21_C241_n1006, B => 
                           mult_21_C241_n1146, CI => mult_21_C241_n1020, CO => 
                           mult_21_C241_n424, S => mult_21_C241_n425);
   mult_21_C241_U281 : ADFULD1 port map( A => mult_21_C241_n1074, B => 
                           mult_21_C241_n1120, CI => mult_21_C241_n1096, CO => 
                           mult_21_C241_n422, S => mult_21_C241_n423);
   mult_21_C241_U280 : ADFULD1 port map( A => mult_21_C241_n448, B => 
                           mult_21_C241_n450, CI => mult_21_C241_n446, CO => 
                           mult_21_C241_n420, S => mult_21_C241_n421);
   mult_21_C241_U279 : ADFULD1 port map( A => mult_21_C241_n429, B => 
                           mult_21_C241_n444, CI => mult_21_C241_n423, CO => 
                           mult_21_C241_n418, S => mult_21_C241_n419);
   mult_21_C241_U278 : ADFULD1 port map( A => mult_21_C241_n427, B => 
                           mult_21_C241_n425, CI => mult_21_C241_n442, CO => 
                           mult_21_C241_n416, S => mult_21_C241_n417);
   mult_21_C241_U277 : ADFULD1 port map( A => mult_21_C241_n421, B => 
                           mult_21_C241_n440, CI => mult_21_C241_n438, CO => 
                           mult_21_C241_n414, S => mult_21_C241_n415);
   mult_21_C241_U276 : ADFULD1 port map( A => mult_21_C241_n417, B => 
                           mult_21_C241_n419, CI => mult_21_C241_n436, CO => 
                           mult_21_C241_n412, S => mult_21_C241_n413);
   mult_21_C241_U275 : ADFULD1 port map( A => mult_21_C241_n434, B => 
                           mult_21_C241_n415, CI => mult_21_C241_n413, CO => 
                           mult_21_C241_n410, S => mult_21_C241_n411);
   mult_21_C241_U274 : ADHALFDL port map( A => mult_21_C241_n430, B => 
                           mult_21_C241_n1203, CO => mult_21_C241_n408, S => 
                           mult_21_C241_n409);
   mult_21_C241_U273 : ADFULD1 port map( A => mult_21_C241_n983, B => 
                           mult_21_C241_n1053, CI => mult_21_C241_n993, CO => 
                           mult_21_C241_n406, S => mult_21_C241_n407);
   mult_21_C241_U272 : ADFULD1 port map( A => mult_21_C241_n1173, B => 
                           mult_21_C241_n1035, CI => mult_21_C241_n1145, CO => 
                           mult_21_C241_n404, S => mult_21_C241_n405);
   mult_21_C241_U271 : ADFULD1 port map( A => mult_21_C241_n1005, B => 
                           mult_21_C241_n1119, CI => mult_21_C241_n1019, CO => 
                           mult_21_C241_n402, S => mult_21_C241_n403);
   mult_21_C241_U270 : ADFULD1 port map( A => mult_21_C241_n1073, B => 
                           mult_21_C241_n1095, CI => mult_21_C241_n409, CO => 
                           mult_21_C241_n400, S => mult_21_C241_n401);
   mult_21_C241_U269 : ADFULD1 port map( A => mult_21_C241_n426, B => 
                           mult_21_C241_n428, CI => mult_21_C241_n422, CO => 
                           mult_21_C241_n398, S => mult_21_C241_n399);
   mult_21_C241_U268 : ADFULD1 port map( A => mult_21_C241_n403, B => 
                           mult_21_C241_n424, CI => mult_21_C241_n405, CO => 
                           mult_21_C241_n396, S => mult_21_C241_n397);
   mult_21_C241_U267 : ADFULD1 port map( A => mult_21_C241_n401, B => 
                           mult_21_C241_n407, CI => mult_21_C241_n420, CO => 
                           mult_21_C241_n394, S => mult_21_C241_n395);
   mult_21_C241_U266 : ADFULD1 port map( A => mult_21_C241_n399, B => 
                           mult_21_C241_n418, CI => mult_21_C241_n416, CO => 
                           mult_21_C241_n392, S => mult_21_C241_n393);
   mult_21_C241_U265 : ADFULD1 port map( A => mult_21_C241_n395, B => 
                           mult_21_C241_n397, CI => mult_21_C241_n414, CO => 
                           mult_21_C241_n390, S => mult_21_C241_n391);
   mult_21_C241_U264 : ADFULD1 port map( A => mult_21_C241_n412, B => 
                           mult_21_C241_n393, CI => mult_21_C241_n391, CO => 
                           mult_21_C241_n388, S => mult_21_C241_n389);
   mult_21_C241_U263 : ADHALFDL port map( A => mult_21_C241_n1202, B => 
                           mult_21_C241_n942, CO => mult_21_C241_n386, S => 
                           mult_21_C241_n387);
   mult_21_C241_U262 : ADFULD1 port map( A => mult_21_C241_n1052, B => 
                           mult_21_C241_n974, CI => mult_21_C241_n1172, CO => 
                           mult_21_C241_n384, S => mult_21_C241_n385);
   mult_21_C241_U261 : ADFULD1 port map( A => mult_21_C241_n982, B => 
                           mult_21_C241_n1018, CI => mult_21_C241_n387, CO => 
                           mult_21_C241_n382, S => mult_21_C241_n383);
   mult_21_C241_U260 : ADFULD1 port map( A => mult_21_C241_n992, B => 
                           mult_21_C241_n1144, CI => mult_21_C241_n1118, CO => 
                           mult_21_C241_n380, S => mult_21_C241_n381);
   mult_21_C241_U259 : ADFULD1 port map( A => mult_21_C241_n1004, B => 
                           mult_21_C241_n1094, CI => mult_21_C241_n1034, CO => 
                           mult_21_C241_n378, S => mult_21_C241_n379);
   mult_21_C241_U258 : ADFULD1 port map( A => mult_21_C241_n408, B => 
                           mult_21_C241_n1072, CI => mult_21_C241_n406, CO => 
                           mult_21_C241_n376, S => mult_21_C241_n377);
   mult_21_C241_U257 : ADFULD1 port map( A => mult_21_C241_n402, B => 
                           mult_21_C241_n404, CI => mult_21_C241_n385, CO => 
                           mult_21_C241_n374, S => mult_21_C241_n375);
   mult_21_C241_U256 : ADFULD1 port map( A => mult_21_C241_n383, B => 
                           mult_21_C241_n379, CI => mult_21_C241_n381, CO => 
                           mult_21_C241_n372, S => mult_21_C241_n373);
   mult_21_C241_U255 : ADFULD1 port map( A => mult_21_C241_n398, B => 
                           mult_21_C241_n400, CI => mult_21_C241_n377, CO => 
                           mult_21_C241_n370, S => mult_21_C241_n371);
   mult_21_C241_U254 : ADFULD1 port map( A => mult_21_C241_n375, B => 
                           mult_21_C241_n396, CI => mult_21_C241_n373, CO => 
                           mult_21_C241_n368, S => mult_21_C241_n369);
   mult_21_C241_U253 : ADFULD1 port map( A => mult_21_C241_n371, B => 
                           mult_21_C241_n394, CI => mult_21_C241_n392, CO => 
                           mult_21_C241_n366, S => mult_21_C241_n367);
   mult_21_C241_U252 : ADFULD1 port map( A => mult_21_C241_n390, B => 
                           mult_21_C241_n369, CI => mult_21_C241_n367, CO => 
                           mult_21_C241_n364, S => mult_21_C241_n365);
   mult_21_C241_U251 : ADHALFDL port map( A => mult_21_C241_n386, B => 
                           mult_21_C241_n1201, CO => mult_21_C241_n362, S => 
                           mult_21_C241_n363);
   mult_21_C241_U250 : ADFULD1 port map( A => mult_21_C241_n1171, B => 
                           mult_21_C241_n1051, CI => mult_21_C241_n1143, CO => 
                           mult_21_C241_n360, S => mult_21_C241_n361);
   mult_21_C241_U249 : ADFULD1 port map( A => mult_21_C241_n973, B => 
                           mult_21_C241_n1003, CI => mult_21_C241_n981, CO => 
                           mult_21_C241_n358, S => mult_21_C241_n359);
   mult_21_C241_U248 : ADFULD1 port map( A => mult_21_C241_n991, B => 
                           mult_21_C241_n1117, CI => mult_21_C241_n1017, CO => 
                           mult_21_C241_n356, S => mult_21_C241_n357);
   mult_21_C241_U247 : ADFULD1 port map( A => mult_21_C241_n1033, B => 
                           mult_21_C241_n1093, CI => mult_21_C241_n1071, CO => 
                           mult_21_C241_n354, S => mult_21_C241_n355);
   mult_21_C241_U246 : ADFULD1 port map( A => mult_21_C241_n384, B => 
                           mult_21_C241_n363, CI => mult_21_C241_n382, CO => 
                           mult_21_C241_n352, S => mult_21_C241_n353);
   mult_21_C241_U245 : ADFULD1 port map( A => mult_21_C241_n378, B => 
                           mult_21_C241_n380, CI => mult_21_C241_n355, CO => 
                           mult_21_C241_n350, S => mult_21_C241_n351);
   mult_21_C241_U244 : ADFULD1 port map( A => mult_21_C241_n361, B => 
                           mult_21_C241_n357, CI => mult_21_C241_n359, CO => 
                           mult_21_C241_n348, S => mult_21_C241_n349);
   mult_21_C241_U243 : ADFULD1 port map( A => mult_21_C241_n374, B => 
                           mult_21_C241_n376, CI => mult_21_C241_n353, CO => 
                           mult_21_C241_n346, S => mult_21_C241_n347);
   mult_21_C241_U242 : ADFULD1 port map( A => mult_21_C241_n351, B => 
                           mult_21_C241_n372, CI => mult_21_C241_n349, CO => 
                           mult_21_C241_n344, S => mult_21_C241_n345);
   mult_21_C241_U241 : ADFULD1 port map( A => mult_21_C241_n347, B => 
                           mult_21_C241_n370, CI => mult_21_C241_n368, CO => 
                           mult_21_C241_n342, S => mult_21_C241_n343);
   mult_21_C241_U240 : ADFULD1 port map( A => mult_21_C241_n366, B => 
                           mult_21_C241_n345, CI => mult_21_C241_n343, CO => 
                           mult_21_C241_n340, S => mult_21_C241_n341);
   mult_21_C241_U239 : ADHALFDL port map( A => mult_21_C241_n1200, B => 
                           mult_21_C241_n941, CO => mult_21_C241_n338, S => 
                           mult_21_C241_n339);
   mult_21_C241_U238 : ADFULD1 port map( A => mult_21_C241_n1050, B => 
                           mult_21_C241_n966, CI => mult_21_C241_n972, CO => 
                           mult_21_C241_n336, S => mult_21_C241_n337);
   mult_21_C241_U237 : ADFULD1 port map( A => mult_21_C241_n980, B => 
                           mult_21_C241_n1032, CI => mult_21_C241_n339, CO => 
                           mult_21_C241_n334, S => mult_21_C241_n335);
   mult_21_C241_U236 : ADFULD1 port map( A => mult_21_C241_n990, B => 
                           mult_21_C241_n1170, CI => mult_21_C241_n1002, CO => 
                           mult_21_C241_n332, S => mult_21_C241_n333);
   mult_21_C241_U235 : ADFULD1 port map( A => mult_21_C241_n1016, B => 
                           mult_21_C241_n1142, CI => mult_21_C241_n1070, CO => 
                           mult_21_C241_n330, S => mult_21_C241_n331);
   mult_21_C241_U234 : ADFULD1 port map( A => mult_21_C241_n1092, B => 
                           mult_21_C241_n1116, CI => mult_21_C241_n362, CO => 
                           mult_21_C241_n328, S => mult_21_C241_n329);
   mult_21_C241_U233 : ADFULD1 port map( A => mult_21_C241_n354, B => 
                           mult_21_C241_n360, CI => mult_21_C241_n356, CO => 
                           mult_21_C241_n326, S => mult_21_C241_n327);
   mult_21_C241_U232 : ADFULD1 port map( A => mult_21_C241_n337, B => 
                           mult_21_C241_n358, CI => mult_21_C241_n331, CO => 
                           mult_21_C241_n324, S => mult_21_C241_n325);
   mult_21_C241_U231 : ADFULD1 port map( A => mult_21_C241_n333, B => 
                           mult_21_C241_n335, CI => mult_21_C241_n329, CO => 
                           mult_21_C241_n322, S => mult_21_C241_n323);
   mult_21_C241_U230 : ADFULD1 port map( A => mult_21_C241_n350, B => 
                           mult_21_C241_n352, CI => mult_21_C241_n348, CO => 
                           mult_21_C241_n320, S => mult_21_C241_n321);
   mult_21_C241_U229 : ADFULD1 port map( A => mult_21_C241_n325, B => 
                           mult_21_C241_n327, CI => mult_21_C241_n323, CO => 
                           mult_21_C241_n318, S => mult_21_C241_n319);
   mult_21_C241_U228 : ADFULD1 port map( A => mult_21_C241_n344, B => 
                           mult_21_C241_n346, CI => mult_21_C241_n321, CO => 
                           mult_21_C241_n316, S => mult_21_C241_n317);
   mult_21_C241_U227 : ADFULD1 port map( A => mult_21_C241_n342, B => 
                           mult_21_C241_n319, CI => mult_21_C241_n317, CO => 
                           mult_21_C241_n314, S => mult_21_C241_n315);
   mult_21_C241_U226 : ADHALFDL port map( A => mult_21_C241_n338, B => 
                           mult_21_C241_n1199, CO => mult_21_C241_n312, S => 
                           mult_21_C241_n313);
   mult_21_C241_U225 : ADFULD1 port map( A => mult_21_C241_n965, B => 
                           mult_21_C241_n1031, CI => mult_21_C241_n971, CO => 
                           mult_21_C241_n310, S => mult_21_C241_n311);
   mult_21_C241_U224 : ADFULD1 port map( A => mult_21_C241_n979, B => 
                           mult_21_C241_n1049, CI => mult_21_C241_n1169, CO => 
                           mult_21_C241_n308, S => mult_21_C241_n309);
   mult_21_C241_U223 : ADFULD1 port map( A => mult_21_C241_n1141, B => 
                           mult_21_C241_n1001, CI => mult_21_C241_n989, CO => 
                           mult_21_C241_n306, S => mult_21_C241_n307);
   mult_21_C241_U222 : ADFULD1 port map( A => mult_21_C241_n1015, B => 
                           mult_21_C241_n1115, CI => mult_21_C241_n1069, CO => 
                           mult_21_C241_n304, S => mult_21_C241_n305);
   mult_21_C241_U221 : ADFULD1 port map( A => mult_21_C241_n313, B => 
                           mult_21_C241_n1091, CI => mult_21_C241_n336, CO => 
                           mult_21_C241_n302, S => mult_21_C241_n303);
   mult_21_C241_U220 : ADFULD1 port map( A => mult_21_C241_n332, B => 
                           mult_21_C241_n330, CI => mult_21_C241_n334, CO => 
                           mult_21_C241_n300, S => mult_21_C241_n301);
   mult_21_C241_U219 : ADFULD1 port map( A => mult_21_C241_n305, B => 
                           mult_21_C241_n328, CI => mult_21_C241_n311, CO => 
                           mult_21_C241_n298, S => mult_21_C241_n299);
   mult_21_C241_U218 : ADFULD1 port map( A => mult_21_C241_n307, B => 
                           mult_21_C241_n309, CI => mult_21_C241_n326, CO => 
                           mult_21_C241_n296, S => mult_21_C241_n297);
   mult_21_C241_U217 : ADFULD1 port map( A => mult_21_C241_n324, B => 
                           mult_21_C241_n303, CI => mult_21_C241_n301, CO => 
                           mult_21_C241_n294, S => mult_21_C241_n295);
   mult_21_C241_U216 : ADFULD1 port map( A => mult_21_C241_n299, B => 
                           mult_21_C241_n322, CI => mult_21_C241_n320, CO => 
                           mult_21_C241_n292, S => mult_21_C241_n293);
   mult_21_C241_U215 : ADFULD1 port map( A => mult_21_C241_n318, B => 
                           mult_21_C241_n297, CI => mult_21_C241_n295, CO => 
                           mult_21_C241_n290, S => mult_21_C241_n291);
   mult_21_C241_U214 : ADFULD1 port map( A => mult_21_C241_n316, B => 
                           mult_21_C241_n293, CI => mult_21_C241_n291, CO => 
                           mult_21_C241_n288, S => mult_21_C241_n289);
   mult_21_C241_U213 : ADHALFDL port map( A => mult_21_C241_n1198, B => 
                           mult_21_C241_n940, CO => mult_21_C241_n286, S => 
                           mult_21_C241_n287);
   mult_21_C241_U212 : ADFULD1 port map( A => mult_21_C241_n1030, B => 
                           mult_21_C241_n960, CI => mult_21_C241_n1168, CO => 
                           mult_21_C241_n284, S => mult_21_C241_n285);
   mult_21_C241_U211 : ADFULD1 port map( A => mult_21_C241_n1140, B => 
                           mult_21_C241_n1000, CI => mult_21_C241_n287, CO => 
                           mult_21_C241_n282, S => mult_21_C241_n283);
   mult_21_C241_U210 : ADFULD1 port map( A => mult_21_C241_n964, B => 
                           mult_21_C241_n1114, CI => mult_21_C241_n970, CO => 
                           mult_21_C241_n280, S => mult_21_C241_n281);
   mult_21_C241_U209 : ADFULD1 port map( A => mult_21_C241_n978, B => 
                           mult_21_C241_n1090, CI => mult_21_C241_n988, CO => 
                           mult_21_C241_n278, S => mult_21_C241_n279);
   mult_21_C241_U208 : ADFULD1 port map( A => mult_21_C241_n1014, B => 
                           mult_21_C241_n1068, CI => mult_21_C241_n1048, CO => 
                           mult_21_C241_n276, S => mult_21_C241_n277);
   mult_21_C241_U207 : ADFULD1 port map( A => mult_21_C241_n304, B => 
                           mult_21_C241_n312, CI => mult_21_C241_n306, CO => 
                           mult_21_C241_n274, S => mult_21_C241_n275);
   mult_21_C241_U206 : ADFULD1 port map( A => mult_21_C241_n310, B => 
                           mult_21_C241_n308, CI => mult_21_C241_n285, CO => 
                           mult_21_C241_n272, S => mult_21_C241_n273);
   mult_21_C241_U205 : ADFULD1 port map( A => mult_21_C241_n283, B => 
                           mult_21_C241_n277, CI => mult_21_C241_n279, CO => 
                           mult_21_C241_n270, S => mult_21_C241_n271);
   mult_21_C241_U204 : ADFULD1 port map( A => mult_21_C241_n302, B => 
                           mult_21_C241_n281, CI => mult_21_C241_n300, CO => 
                           mult_21_C241_n268, S => mult_21_C241_n269);
   mult_21_C241_U203 : ADFULD1 port map( A => mult_21_C241_n275, B => 
                           mult_21_C241_n298, CI => mult_21_C241_n273, CO => 
                           mult_21_C241_n266, S => mult_21_C241_n267);
   mult_21_C241_U202 : ADFULD1 port map( A => mult_21_C241_n296, B => 
                           mult_21_C241_n271, CI => mult_21_C241_n269, CO => 
                           mult_21_C241_n264, S => mult_21_C241_n265);
   mult_21_C241_U201 : ADFULD1 port map( A => mult_21_C241_n267, B => 
                           mult_21_C241_n294, CI => mult_21_C241_n292, CO => 
                           mult_21_C241_n262, S => mult_21_C241_n263);
   mult_21_C241_U200 : ADFULD1 port map( A => mult_21_C241_n290, B => 
                           mult_21_C241_n265, CI => mult_21_C241_n263, CO => 
                           mult_21_C241_n260, S => mult_21_C241_n261);
   mult_21_C241_U199 : ADHALFDL port map( A => mult_21_C241_n286, B => 
                           mult_21_C241_n1197, CO => mult_21_C241_n258, S => 
                           mult_21_C241_n259);
   mult_21_C241_U198 : ADFULD1 port map( A => mult_21_C241_n1167, B => 
                           mult_21_C241_n1029, CI => mult_21_C241_n1139, CO => 
                           mult_21_C241_n256, S => mult_21_C241_n257);
   mult_21_C241_U197 : ADFULD1 port map( A => mult_21_C241_n1113, B => 
                           mult_21_C241_n987, CI => mult_21_C241_n1089, CO => 
                           mult_21_C241_n254, S => mult_21_C241_n255);
   mult_21_C241_U196 : ADFULD1 port map( A => mult_21_C241_n959, B => 
                           mult_21_C241_n969, CI => mult_21_C241_n963, CO => 
                           mult_21_C241_n252, S => mult_21_C241_n253);
   mult_21_C241_U195 : ADFULD1 port map( A => mult_21_C241_n977, B => 
                           mult_21_C241_n1067, CI => mult_21_C241_n999, CO => 
                           mult_21_C241_n250, S => mult_21_C241_n251);
   mult_21_C241_U194 : ADFULD1 port map( A => mult_21_C241_n1047, B => 
                           mult_21_C241_n1013, CI => mult_21_C241_n259, CO => 
                           mult_21_C241_n248, S => mult_21_C241_n249);
   mult_21_C241_U193 : ADFULD1 port map( A => mult_21_C241_n278, B => 
                           mult_21_C241_n284, CI => mult_21_C241_n282, CO => 
                           mult_21_C241_n246, S => mult_21_C241_n247);
   mult_21_C241_U192 : ADFULD1 port map( A => mult_21_C241_n280, B => 
                           mult_21_C241_n276, CI => mult_21_C241_n251, CO => 
                           mult_21_C241_n244, S => mult_21_C241_n245);
   mult_21_C241_U191 : ADFULD1 port map( A => mult_21_C241_n253, B => 
                           mult_21_C241_n255, CI => mult_21_C241_n257, CO => 
                           mult_21_C241_n242, S => mult_21_C241_n243);
   mult_21_C241_U190 : ADFULD1 port map( A => mult_21_C241_n274, B => 
                           mult_21_C241_n249, CI => mult_21_C241_n272, CO => 
                           mult_21_C241_n240, S => mult_21_C241_n241);
   mult_21_C241_U189 : ADFULD1 port map( A => mult_21_C241_n270, B => 
                           mult_21_C241_n247, CI => mult_21_C241_n245, CO => 
                           mult_21_C241_n238, S => mult_21_C241_n239);
   mult_21_C241_U188 : ADFULD1 port map( A => mult_21_C241_n268, B => 
                           mult_21_C241_n243, CI => mult_21_C241_n241, CO => 
                           mult_21_C241_n236, S => mult_21_C241_n237);
   mult_21_C241_U187 : ADFULD1 port map( A => mult_21_C241_n239, B => 
                           mult_21_C241_n266, CI => mult_21_C241_n264, CO => 
                           mult_21_C241_n234, S => mult_21_C241_n235);
   mult_21_C241_U186 : ADFULD1 port map( A => mult_21_C241_n262, B => 
                           mult_21_C241_n237, CI => mult_21_C241_n235, CO => 
                           mult_21_C241_n232, S => mult_21_C241_n233);
   mult_21_C241_U185 : ADHALFDL port map( A => mult_21_C241_n1196, B => 
                           mult_21_C241_n939, CO => mult_21_C241_n230, S => 
                           mult_21_C241_n231);
   mult_21_C241_U184 : ADFULD1 port map( A => mult_21_C241_n1028, B => 
                           mult_21_C241_n956, CI => mult_21_C241_n958, CO => 
                           mult_21_C241_n228, S => mult_21_C241_n229);
   mult_21_C241_U183 : ADFULD1 port map( A => mult_21_C241_n1166, B => 
                           mult_21_C241_n1012, CI => mult_21_C241_n231, CO => 
                           mult_21_C241_n226, S => mult_21_C241_n227);
   mult_21_C241_U182 : ADFULD1 port map( A => mult_21_C241_n962, B => 
                           mult_21_C241_n1138, CI => mult_21_C241_n968, CO => 
                           mult_21_C241_n224, S => mult_21_C241_n225);
   mult_21_C241_U181 : ADFULD1 port map( A => mult_21_C241_n986, B => 
                           mult_21_C241_n976, CI => mult_21_C241_n998, CO => 
                           mult_21_C241_n222, S => mult_21_C241_n223);
   mult_21_C241_U180 : ADFULD1 port map( A => mult_21_C241_n1046, B => 
                           mult_21_C241_n1112, CI => mult_21_C241_n1066, CO => 
                           mult_21_C241_n220, S => mult_21_C241_n221);
   mult_21_C241_U179 : ADFULD1 port map( A => mult_21_C241_n258, B => 
                           mult_21_C241_n1088, CI => mult_21_C241_n250, CO => 
                           mult_21_C241_n218, S => mult_21_C241_n219);
   mult_21_C241_U178 : ADFULD1 port map( A => mult_21_C241_n256, B => 
                           mult_21_C241_n252, CI => mult_21_C241_n254, CO => 
                           mult_21_C241_n216, S => mult_21_C241_n217);
   mult_21_C241_U177 : ADFULD1 port map( A => mult_21_C241_n221, B => 
                           mult_21_C241_n229, CI => mult_21_C241_n227, CO => 
                           mult_21_C241_n214, S => mult_21_C241_n215);
   mult_21_C241_U176 : ADFULD1 port map( A => mult_21_C241_n225, B => 
                           mult_21_C241_n223, CI => mult_21_C241_n248, CO => 
                           mult_21_C241_n212, S => mult_21_C241_n213);
   mult_21_C241_U175 : ADFULD1 port map( A => mult_21_C241_n244, B => 
                           mult_21_C241_n246, CI => mult_21_C241_n219, CO => 
                           mult_21_C241_n210, S => mult_21_C241_n211);
   mult_21_C241_U174 : ADFULD1 port map( A => mult_21_C241_n217, B => 
                           mult_21_C241_n242, CI => mult_21_C241_n215, CO => 
                           mult_21_C241_n208, S => mult_21_C241_n209);
   mult_21_C241_U173 : ADFULD1 port map( A => mult_21_C241_n240, B => 
                           mult_21_C241_n213, CI => mult_21_C241_n238, CO => 
                           mult_21_C241_n206, S => mult_21_C241_n207);
   mult_21_C241_U172 : ADFULD1 port map( A => mult_21_C241_n209, B => 
                           mult_21_C241_n211, CI => mult_21_C241_n236, CO => 
                           mult_21_C241_n204, S => mult_21_C241_n205);
   mult_21_C241_U171 : ADFULD1 port map( A => mult_21_C241_n234, B => 
                           mult_21_C241_n207, CI => mult_21_C241_n205, CO => 
                           mult_21_C241_n202, S => mult_21_C241_n203);
   mult_21_C241_U155 : ADHALFDL port map( A => mult_21_C241_n1226, B => N2914, 
                           CO => mult_21_C241_n186, S => N3233);
   mult_21_C241_U154 : ADHALFDL port map( A => mult_21_C241_n186, B => 
                           mult_21_C241_n1225, CO => mult_21_C241_n185, S => 
                           N3234);
   mult_21_C241_U153 : ADFULD1 port map( A => mult_21_C241_n651, B => 
                           mult_21_C241_n1194, CI => mult_21_C241_n185, CO => 
                           mult_21_C241_n184, S => N3235);
   mult_21_C241_U152 : ADFULD1 port map( A => mult_21_C241_n649, B => 
                           mult_21_C241_n1193, CI => mult_21_C241_n184, CO => 
                           mult_21_C241_n183, S => N3236);
   mult_21_C241_U151 : ADFULD1 port map( A => mult_21_C241_n645, B => 
                           mult_21_C241_n648, CI => mult_21_C241_n183, CO => 
                           mult_21_C241_n182, S => N3237);
   mult_21_C241_U150 : ADFULD1 port map( A => mult_21_C241_n641, B => 
                           mult_21_C241_n644, CI => mult_21_C241_n182, CO => 
                           mult_21_C241_n181, S => N3238);
   mult_21_C241_U149 : ADFULD1 port map( A => mult_21_C241_n635, B => 
                           mult_21_C241_n640, CI => mult_21_C241_n181, CO => 
                           mult_21_C241_n180, S => N3239);
   mult_21_C241_U148 : ADFULD1 port map( A => mult_21_C241_n629, B => 
                           mult_21_C241_n634, CI => mult_21_C241_n180, CO => 
                           mult_21_C241_n179, S => N3240);
   mult_21_C241_U147 : ADFULD1 port map( A => mult_21_C241_n621, B => 
                           mult_21_C241_n628, CI => mult_21_C241_n179, CO => 
                           mult_21_C241_n178, S => N3241);
   mult_21_C241_U146 : ADFULD1 port map( A => mult_21_C241_n613, B => 
                           mult_21_C241_n620, CI => mult_21_C241_n178, CO => 
                           mult_21_C241_n177, S => N3242);
   mult_21_C241_U145 : ADFULD1 port map( A => mult_21_C241_n603, B => 
                           mult_21_C241_n612, CI => mult_21_C241_n177, CO => 
                           mult_21_C241_n176, S => N3243);
   mult_21_C241_U144 : ADFULD1 port map( A => mult_21_C241_n593, B => 
                           mult_21_C241_n602, CI => mult_21_C241_n176, CO => 
                           mult_21_C241_n175, S => N3244);
   mult_21_C241_U143 : ADFULD1 port map( A => mult_21_C241_n581, B => 
                           mult_21_C241_n592, CI => mult_21_C241_n175, CO => 
                           mult_21_C241_n174, S => N3245);
   mult_21_C241_U142 : ADFULD1 port map( A => mult_21_C241_n569, B => 
                           mult_21_C241_n580, CI => mult_21_C241_n174, CO => 
                           mult_21_C241_n173, S => N3246);
   mult_21_C241_U141 : ADFULD1 port map( A => mult_21_C241_n555, B => 
                           mult_21_C241_n568, CI => mult_21_C241_n173, CO => 
                           mult_21_C241_n172, S => N3247);
   mult_21_C241_U140 : ADFULD1 port map( A => mult_21_C241_n541, B => 
                           mult_21_C241_n554, CI => mult_21_C241_n172, CO => 
                           mult_21_C241_n171, S => N3248);
   mult_21_C241_U139 : ADFULD1 port map( A => mult_21_C241_n525, B => 
                           mult_21_C241_n540, CI => mult_21_C241_n171, CO => 
                           mult_21_C241_n170, S => N3249);
   mult_21_C241_U138 : ADFULD1 port map( A => mult_21_C241_n509, B => 
                           mult_21_C241_n524, CI => mult_21_C241_n170, CO => 
                           mult_21_C241_n169, S => N3250);
   mult_21_C241_U137 : ADFULD1 port map( A => mult_21_C241_n491, B => 
                           mult_21_C241_n508, CI => mult_21_C241_n169, CO => 
                           mult_21_C241_n168, S => N3251);
   mult_21_C241_U136 : ADFULD1 port map( A => mult_21_C241_n473, B => 
                           mult_21_C241_n490, CI => mult_21_C241_n168, CO => 
                           mult_21_C241_n167, S => N3252);
   mult_21_C241_U135 : ADFULD1 port map( A => mult_21_C241_n453, B => 
                           mult_21_C241_n472, CI => mult_21_C241_n167, CO => 
                           mult_21_C241_n166, S => N3253);
   mult_21_C241_U134 : ADFULD1 port map( A => mult_21_C241_n433, B => 
                           mult_21_C241_n452, CI => mult_21_C241_n166, CO => 
                           mult_21_C241_n165, S => N3254);
   mult_21_C241_U133 : ADFULD1 port map( A => mult_21_C241_n411, B => 
                           mult_21_C241_n432, CI => mult_21_C241_n165, CO => 
                           mult_21_C241_n164, S => N3255);
   mult_21_C241_U132 : ADFULD1 port map( A => mult_21_C241_n389, B => 
                           mult_21_C241_n410, CI => mult_21_C241_n164, CO => 
                           mult_21_C241_n163, S => N3256);
   mult_21_C241_U131 : ADFULD1 port map( A => mult_21_C241_n365, B => 
                           mult_21_C241_n388, CI => mult_21_C241_n163, CO => 
                           mult_21_C241_n162, S => N3257);
   mult_21_C241_U130 : ADFULD1 port map( A => mult_21_C241_n341, B => 
                           mult_21_C241_n364, CI => mult_21_C241_n162, CO => 
                           mult_21_C241_n161, S => N3258);
   mult_21_C241_U129 : ADFULD1 port map( A => mult_21_C241_n315, B => 
                           mult_21_C241_n340, CI => mult_21_C241_n161, CO => 
                           mult_21_C241_n160, S => N3259);
   mult_21_C241_U128 : ADFULD1 port map( A => mult_21_C241_n289, B => 
                           mult_21_C241_n314, CI => mult_21_C241_n160, CO => 
                           mult_21_C241_n159, S => N3260);
   mult_21_C241_U127 : ADFULD1 port map( A => mult_21_C241_n261, B => 
                           mult_21_C241_n288, CI => mult_21_C241_n159, CO => 
                           mult_21_C241_n158, S => N3261);
   mult_21_C241_U126 : ADFULD1 port map( A => mult_21_C241_n233, B => 
                           mult_21_C241_n260, CI => mult_21_C241_n158, CO => 
                           mult_21_C241_n157, S => N3262);
   mult_21_C241_U125 : ADFULD1 port map( A => mult_21_C241_n203, B => 
                           mult_21_C241_n232, CI => mult_21_C241_n157, CO => 
                           mult_21_C241_n156, S => N3263);
   mult_21_C243_U1396 : AOI21D1 port map( A1 => N2972, A2 => N2973, B => 
                           mult_21_C243_n1421, Z => mult_21_C243_n940);
   mult_21_C243_U1395 : OAI21D1 port map( A1 => N2975, A2 => N2974, B => 
                           mult_21_C243_n1422, Z => mult_21_C243_n104);
   mult_21_C243_U1394 : AOI21D1 port map( A1 => N2974, A2 => N2975, B => 
                           mult_21_C243_n1422, Z => mult_21_C243_n939);
   mult_21_C243_U1393 : AOI21D1 port map( A1 => N2946, A2 => N2947, B => 
                           mult_21_C243_n1395, Z => mult_21_C243_n953);
   mult_21_C243_U1392 : AOI21D1 port map( A1 => N2948, A2 => N2949, B => 
                           mult_21_C243_n1397, Z => mult_21_C243_n952);
   mult_21_C243_U1391 : AOI21D1 port map( A1 => N2950, A2 => N2951, B => 
                           mult_21_C243_n1399, Z => mult_21_C243_n951);
   mult_21_C243_U1390 : AOI21D1 port map( A1 => N2952, A2 => N2953, B => 
                           mult_21_C243_n1401, Z => mult_21_C243_n950);
   mult_21_C243_U1389 : AOI21D1 port map( A1 => N2954, A2 => N2955, B => 
                           mult_21_C243_n1403, Z => mult_21_C243_n949);
   mult_21_C243_U1388 : AOI21D1 port map( A1 => N2956, A2 => N2957, B => 
                           mult_21_C243_n1405, Z => mult_21_C243_n948);
   mult_21_C243_U1387 : AOI21D1 port map( A1 => N2958, A2 => N2959, B => 
                           mult_21_C243_n1407, Z => mult_21_C243_n947);
   mult_21_C243_U1386 : EXOR2D1 port map( A1 => N2975, A2 => N2974, Z => 
                           mult_21_C243_n1451);
   mult_21_C243_U1385 : MUXB2DL port map( A0 => N3105, A1 => N3106, SL => 
                           mult_21_C243_n1451, Z => mult_21_C243_n652);
   mult_21_C243_U1384 : NAN2D1 port map( A1 => N3105, A2 => mult_21_C243_n1451,
                           Z => mult_21_C243_n653);
   mult_21_C243_U1383 : EXOR2D1 port map( A1 => N2973, A2 => N2972, Z => 
                           mult_21_C243_n1450);
   mult_21_C243_U1382 : MUXB2DL port map( A0 => N3107, A1 => N3108, SL => 
                           mult_21_C243_n1450, Z => mult_21_C243_n654);
   mult_21_C243_U1381 : MUXB2DL port map( A0 => mult_21_C243_n1388, A1 => N3107
                           , SL => mult_21_C243_n1450, Z => mult_21_C243_n655);
   mult_21_C243_U1380 : MUXB2DL port map( A0 => N3105, A1 => N3106, SL => 
                           mult_21_C243_n1450, Z => mult_21_C243_n656);
   mult_21_C243_U1379 : NAN2D1 port map( A1 => N3105, A2 => mult_21_C243_n1450,
                           Z => mult_21_C243_n657);
   mult_21_C243_U1378 : EXOR2D1 port map( A1 => N2971, A2 => N2970, Z => 
                           mult_21_C243_n1449);
   mult_21_C243_U1377 : MUXB2DL port map( A0 => N3109, A1 => N3110, SL => 
                           mult_21_C243_n1449, Z => mult_21_C243_n658);
   mult_21_C243_U1376 : MUXB2DL port map( A0 => mult_21_C243_n1386, A1 => N3109
                           , SL => mult_21_C243_n1449, Z => mult_21_C243_n659);
   mult_21_C243_U1375 : MUXB2DL port map( A0 => N3107, A1 => N3108, SL => 
                           mult_21_C243_n1449, Z => mult_21_C243_n660);
   mult_21_C243_U1374 : MUXB2DL port map( A0 => mult_21_C243_n1388, A1 => N3107
                           , SL => mult_21_C243_n1449, Z => mult_21_C243_n661);
   mult_21_C243_U1373 : MUXB2DL port map( A0 => N3105, A1 => N3106, SL => 
                           mult_21_C243_n1449, Z => mult_21_C243_n662);
   mult_21_C243_U1372 : NAN2D1 port map( A1 => N3105, A2 => mult_21_C243_n1449,
                           Z => mult_21_C243_n663);
   mult_21_C243_U1371 : EXOR2D1 port map( A1 => N2969, A2 => N2968, Z => 
                           mult_21_C243_n1448);
   mult_21_C243_U1370 : MUXB2DL port map( A0 => N3111, A1 => N3112, SL => 
                           mult_21_C243_n1448, Z => mult_21_C243_n664);
   mult_21_C243_U1369 : MUXB2DL port map( A0 => N3110, A1 => N3111, SL => 
                           mult_21_C243_n1448, Z => mult_21_C243_n665);
   mult_21_C243_U1368 : MUXB2DL port map( A0 => N3109, A1 => N3110, SL => 
                           mult_21_C243_n1448, Z => mult_21_C243_n666);
   mult_21_C243_U1367 : MUXB2DL port map( A0 => mult_21_C243_n1386, A1 => N3109
                           , SL => mult_21_C243_n1448, Z => mult_21_C243_n667);
   mult_21_C243_U1366 : MUXB2DL port map( A0 => N3107, A1 => N3108, SL => 
                           mult_21_C243_n1448, Z => mult_21_C243_n668);
   mult_21_C243_U1365 : MUXB2DL port map( A0 => mult_21_C243_n1388, A1 => N3107
                           , SL => mult_21_C243_n1448, Z => mult_21_C243_n669);
   mult_21_C243_U1364 : MUXB2DL port map( A0 => N3105, A1 => N3106, SL => 
                           mult_21_C243_n1448, Z => mult_21_C243_n670);
   mult_21_C243_U1363 : NAN2D1 port map( A1 => N3105, A2 => mult_21_C243_n1448,
                           Z => mult_21_C243_n671);
   mult_21_C243_U1362 : MUXB2DL port map( A0 => N3113, A1 => N3114, SL => 
                           mult_21_C243_n1447, Z => mult_21_C243_n672);
   mult_21_C243_U1361 : MUXB2DL port map( A0 => N3112, A1 => N3113, SL => 
                           mult_21_C243_n1447, Z => mult_21_C243_n673);
   mult_21_C243_U1360 : MUXB2DL port map( A0 => N3111, A1 => N3112, SL => 
                           mult_21_C243_n1447, Z => mult_21_C243_n674);
   mult_21_C243_U1359 : MUXB2DL port map( A0 => N3110, A1 => N3111, SL => 
                           mult_21_C243_n1447, Z => mult_21_C243_n675);
   mult_21_C243_U1358 : MUXB2DL port map( A0 => N3109, A1 => N3110, SL => 
                           mult_21_C243_n1447, Z => mult_21_C243_n676);
   mult_21_C243_U1357 : MUXB2DL port map( A0 => mult_21_C243_n1386, A1 => N3109
                           , SL => mult_21_C243_n1447, Z => mult_21_C243_n677);
   mult_21_C243_U1356 : MUXB2DL port map( A0 => N3107, A1 => N3108, SL => 
                           mult_21_C243_n1447, Z => mult_21_C243_n678);
   mult_21_C243_U1355 : MUXB2DL port map( A0 => mult_21_C243_n1388, A1 => N3107
                           , SL => mult_21_C243_n1447, Z => mult_21_C243_n679);
   mult_21_C243_U1354 : AOI21D1 port map( A1 => N2960, A2 => N2961, B => 
                           mult_21_C243_n1409, Z => mult_21_C243_n946);
   mult_21_C243_U1353 : MUXB2DL port map( A0 => N3105, A1 => N3106, SL => 
                           mult_21_C243_n1447, Z => mult_21_C243_n680);
   mult_21_C243_U1352 : NAN2D1 port map( A1 => N3105, A2 => mult_21_C243_n1447,
                           Z => mult_21_C243_n681);
   mult_21_C243_U1351 : MUXB2DL port map( A0 => N3115, A1 => N3116, SL => 
                           mult_21_C243_n1446, Z => mult_21_C243_n682);
   mult_21_C243_U1350 : MUXB2DL port map( A0 => N3114, A1 => N3115, SL => 
                           mult_21_C243_n1446, Z => mult_21_C243_n683);
   mult_21_C243_U1349 : MUXB2DL port map( A0 => N3113, A1 => N3114, SL => 
                           mult_21_C243_n1446, Z => mult_21_C243_n684);
   mult_21_C243_U1348 : MUXB2DL port map( A0 => N3112, A1 => N3113, SL => 
                           mult_21_C243_n1446, Z => mult_21_C243_n685);
   mult_21_C243_U1347 : MUXB2DL port map( A0 => N3111, A1 => N3112, SL => 
                           mult_21_C243_n1446, Z => mult_21_C243_n686);
   mult_21_C243_U1346 : MUXB2DL port map( A0 => N3110, A1 => N3111, SL => 
                           mult_21_C243_n1446, Z => mult_21_C243_n687);
   mult_21_C243_U1345 : MUXB2DL port map( A0 => N3109, A1 => N3110, SL => 
                           mult_21_C243_n1446, Z => mult_21_C243_n688);
   mult_21_C243_U1344 : MUXB2DL port map( A0 => mult_21_C243_n1386, A1 => N3109
                           , SL => mult_21_C243_n1446, Z => mult_21_C243_n689);
   mult_21_C243_U1343 : MUXB2DL port map( A0 => N3107, A1 => N3108, SL => 
                           mult_21_C243_n1446, Z => mult_21_C243_n690);
   mult_21_C243_U1342 : MUXB2DL port map( A0 => mult_21_C243_n1388, A1 => N3107
                           , SL => mult_21_C243_n1446, Z => mult_21_C243_n691);
   mult_21_C243_U1341 : MUXB2DL port map( A0 => N3105, A1 => N3106, SL => 
                           mult_21_C243_n1446, Z => mult_21_C243_n692);
   mult_21_C243_U1340 : NAN2D1 port map( A1 => N3105, A2 => mult_21_C243_n1446,
                           Z => mult_21_C243_n693);
   mult_21_C243_U1339 : MUXB2DL port map( A0 => N3117, A1 => N3118, SL => 
                           mult_21_C243_n1445, Z => mult_21_C243_n694);
   mult_21_C243_U1338 : MUXB2DL port map( A0 => N3116, A1 => N3117, SL => 
                           mult_21_C243_n1445, Z => mult_21_C243_n695);
   mult_21_C243_U1337 : MUXB2DL port map( A0 => N3115, A1 => N3116, SL => 
                           mult_21_C243_n1445, Z => mult_21_C243_n696);
   mult_21_C243_U1336 : MUXB2DL port map( A0 => N3114, A1 => N3115, SL => 
                           mult_21_C243_n1445, Z => mult_21_C243_n697);
   mult_21_C243_U1335 : MUXB2DL port map( A0 => N3113, A1 => N3114, SL => 
                           mult_21_C243_n1445, Z => mult_21_C243_n698);
   mult_21_C243_U1334 : MUXB2DL port map( A0 => N3112, A1 => N3113, SL => 
                           mult_21_C243_n1445, Z => mult_21_C243_n699);
   mult_21_C243_U1333 : MUXB2DL port map( A0 => N3111, A1 => N3112, SL => 
                           mult_21_C243_n1445, Z => mult_21_C243_n700);
   mult_21_C243_U1332 : MUXB2DL port map( A0 => N3110, A1 => N3111, SL => 
                           mult_21_C243_n1445, Z => mult_21_C243_n701);
   mult_21_C243_U1331 : MUXB2DL port map( A0 => N3109, A1 => N3110, SL => 
                           mult_21_C243_n1445, Z => mult_21_C243_n702);
   mult_21_C243_U1330 : MUXB2DL port map( A0 => mult_21_C243_n1386, A1 => N3109
                           , SL => mult_21_C243_n1445, Z => mult_21_C243_n703);
   mult_21_C243_U1329 : MUXB2DL port map( A0 => N3107, A1 => N3108, SL => 
                           mult_21_C243_n1445, Z => mult_21_C243_n704);
   mult_21_C243_U1328 : MUXB2DL port map( A0 => mult_21_C243_n1388, A1 => N3107
                           , SL => mult_21_C243_n1445, Z => mult_21_C243_n705);
   mult_21_C243_U1327 : MUXB2DL port map( A0 => N3105, A1 => N3106, SL => 
                           mult_21_C243_n1445, Z => mult_21_C243_n706);
   mult_21_C243_U1326 : NAN2D1 port map( A1 => N3105, A2 => mult_21_C243_n1445,
                           Z => mult_21_C243_n707);
   mult_21_C243_U1325 : MUXB2DL port map( A0 => N3119, A1 => N3120, SL => 
                           mult_21_C243_n1444, Z => mult_21_C243_n708);
   mult_21_C243_U1324 : MUXB2DL port map( A0 => N3118, A1 => N3119, SL => 
                           mult_21_C243_n1444, Z => mult_21_C243_n709);
   mult_21_C243_U1323 : MUXB2DL port map( A0 => N3117, A1 => N3118, SL => 
                           mult_21_C243_n1444, Z => mult_21_C243_n710);
   mult_21_C243_U1322 : MUXB2DL port map( A0 => N3116, A1 => N3117, SL => 
                           mult_21_C243_n1444, Z => mult_21_C243_n711);
   mult_21_C243_U1321 : MUXB2DL port map( A0 => N3115, A1 => N3116, SL => 
                           mult_21_C243_n1444, Z => mult_21_C243_n712);
   mult_21_C243_U1320 : MUXB2DL port map( A0 => N3114, A1 => N3115, SL => 
                           mult_21_C243_n1444, Z => mult_21_C243_n713);
   mult_21_C243_U1319 : MUXB2DL port map( A0 => N3113, A1 => N3114, SL => 
                           mult_21_C243_n1444, Z => mult_21_C243_n714);
   mult_21_C243_U1318 : MUXB2DL port map( A0 => N3112, A1 => N3113, SL => 
                           mult_21_C243_n1444, Z => mult_21_C243_n715);
   mult_21_C243_U1317 : MUXB2DL port map( A0 => N3111, A1 => N3112, SL => 
                           mult_21_C243_n1444, Z => mult_21_C243_n716);
   mult_21_C243_U1316 : MUXB2DL port map( A0 => N3110, A1 => N3111, SL => 
                           mult_21_C243_n1444, Z => mult_21_C243_n717);
   mult_21_C243_U1315 : MUXB2DL port map( A0 => N3109, A1 => N3110, SL => 
                           mult_21_C243_n1444, Z => mult_21_C243_n718);
   mult_21_C243_U1314 : MUXB2DL port map( A0 => mult_21_C243_n1386, A1 => N3109
                           , SL => mult_21_C243_n1444, Z => mult_21_C243_n719);
   mult_21_C243_U1313 : MUXB2DL port map( A0 => N3107, A1 => N3108, SL => 
                           mult_21_C243_n1444, Z => mult_21_C243_n720);
   mult_21_C243_U1312 : MUXB2DL port map( A0 => mult_21_C243_n1388, A1 => N3107
                           , SL => mult_21_C243_n1444, Z => mult_21_C243_n721);
   mult_21_C243_U1311 : MUXB2DL port map( A0 => N3105, A1 => N3106, SL => 
                           mult_21_C243_n1444, Z => mult_21_C243_n722);
   mult_21_C243_U1310 : NAN2D1 port map( A1 => N3105, A2 => mult_21_C243_n1444,
                           Z => mult_21_C243_n723);
   mult_21_C243_U1309 : MUXB2DL port map( A0 => N3121, A1 => N3122, SL => 
                           mult_21_C243_n1443, Z => mult_21_C243_n724);
   mult_21_C243_U1308 : MUXB2DL port map( A0 => N3120, A1 => N3121, SL => 
                           mult_21_C243_n1443, Z => mult_21_C243_n725);
   mult_21_C243_U1307 : MUXB2DL port map( A0 => N3119, A1 => N3120, SL => 
                           mult_21_C243_n1443, Z => mult_21_C243_n726);
   mult_21_C243_U1306 : MUXB2DL port map( A0 => N3118, A1 => N3119, SL => 
                           mult_21_C243_n1443, Z => mult_21_C243_n727);
   mult_21_C243_U1305 : MUXB2DL port map( A0 => N3117, A1 => N3118, SL => 
                           mult_21_C243_n1443, Z => mult_21_C243_n728);
   mult_21_C243_U1304 : MUXB2DL port map( A0 => N3116, A1 => N3117, SL => 
                           mult_21_C243_n1443, Z => mult_21_C243_n729);
   mult_21_C243_U1303 : MUXB2DL port map( A0 => N3115, A1 => N3116, SL => 
                           mult_21_C243_n1443, Z => mult_21_C243_n730);
   mult_21_C243_U1302 : MUXB2DL port map( A0 => N3114, A1 => N3115, SL => 
                           mult_21_C243_n1443, Z => mult_21_C243_n731);
   mult_21_C243_U1301 : MUXB2DL port map( A0 => N3113, A1 => N3114, SL => 
                           mult_21_C243_n1443, Z => mult_21_C243_n732);
   mult_21_C243_U1300 : MUXB2DL port map( A0 => N3112, A1 => N3113, SL => 
                           mult_21_C243_n1443, Z => mult_21_C243_n733);
   mult_21_C243_U1299 : MUXB2DL port map( A0 => N3111, A1 => N3112, SL => 
                           mult_21_C243_n1443, Z => mult_21_C243_n734);
   mult_21_C243_U1298 : MUXB2DL port map( A0 => N3110, A1 => N3111, SL => 
                           mult_21_C243_n1443, Z => mult_21_C243_n735);
   mult_21_C243_U1297 : MUXB2DL port map( A0 => N3109, A1 => N3110, SL => 
                           mult_21_C243_n1443, Z => mult_21_C243_n736);
   mult_21_C243_U1296 : MUXB2DL port map( A0 => mult_21_C243_n1386, A1 => N3109
                           , SL => mult_21_C243_n1443, Z => mult_21_C243_n737);
   mult_21_C243_U1295 : MUXB2DL port map( A0 => N3107, A1 => N3108, SL => 
                           mult_21_C243_n1443, Z => mult_21_C243_n738);
   mult_21_C243_U1294 : MUXB2DL port map( A0 => mult_21_C243_n1388, A1 => N3107
                           , SL => mult_21_C243_n1443, Z => mult_21_C243_n739);
   mult_21_C243_U1293 : MUXB2DL port map( A0 => N3105, A1 => N3106, SL => 
                           mult_21_C243_n1443, Z => mult_21_C243_n740);
   mult_21_C243_U1292 : NAN2D1 port map( A1 => N3105, A2 => mult_21_C243_n1443,
                           Z => mult_21_C243_n741);
   mult_21_C243_U1291 : MUXB2DL port map( A0 => N3123, A1 => N3124, SL => 
                           mult_21_C243_n1442, Z => mult_21_C243_n742);
   mult_21_C243_U1290 : MUXB2DL port map( A0 => N3122, A1 => N3123, SL => 
                           mult_21_C243_n1442, Z => mult_21_C243_n743);
   mult_21_C243_U1289 : MUXB2DL port map( A0 => N3121, A1 => N3122, SL => 
                           mult_21_C243_n1442, Z => mult_21_C243_n744);
   mult_21_C243_U1288 : MUXB2DL port map( A0 => N3120, A1 => N3121, SL => 
                           mult_21_C243_n1442, Z => mult_21_C243_n745);
   mult_21_C243_U1287 : MUXB2DL port map( A0 => N3119, A1 => N3120, SL => 
                           mult_21_C243_n1442, Z => mult_21_C243_n746);
   mult_21_C243_U1286 : MUXB2DL port map( A0 => N3118, A1 => N3119, SL => 
                           mult_21_C243_n1442, Z => mult_21_C243_n747);
   mult_21_C243_U1285 : MUXB2DL port map( A0 => N3117, A1 => N3118, SL => 
                           mult_21_C243_n1442, Z => mult_21_C243_n748);
   mult_21_C243_U1284 : MUXB2DL port map( A0 => N3116, A1 => N3117, SL => 
                           mult_21_C243_n1442, Z => mult_21_C243_n749);
   mult_21_C243_U1283 : AOI21D1 port map( A1 => N2962, A2 => N2963, B => 
                           mult_21_C243_n1411, Z => mult_21_C243_n945);
   mult_21_C243_U1282 : MUXB2DL port map( A0 => N3115, A1 => N3116, SL => 
                           mult_21_C243_n1442, Z => mult_21_C243_n750);
   mult_21_C243_U1281 : MUXB2DL port map( A0 => N3114, A1 => N3115, SL => 
                           mult_21_C243_n1442, Z => mult_21_C243_n751);
   mult_21_C243_U1280 : MUXB2DL port map( A0 => N3113, A1 => N3114, SL => 
                           mult_21_C243_n1442, Z => mult_21_C243_n752);
   mult_21_C243_U1279 : MUXB2DL port map( A0 => N3112, A1 => N3113, SL => 
                           mult_21_C243_n1442, Z => mult_21_C243_n753);
   mult_21_C243_U1278 : MUXB2DL port map( A0 => N3111, A1 => N3112, SL => 
                           mult_21_C243_n1442, Z => mult_21_C243_n754);
   mult_21_C243_U1277 : MUXB2DL port map( A0 => N3110, A1 => N3111, SL => 
                           mult_21_C243_n1442, Z => mult_21_C243_n755);
   mult_21_C243_U1276 : MUXB2DL port map( A0 => N3109, A1 => N3110, SL => 
                           mult_21_C243_n1442, Z => mult_21_C243_n756);
   mult_21_C243_U1275 : MUXB2DL port map( A0 => mult_21_C243_n1386, A1 => N3109
                           , SL => mult_21_C243_n1442, Z => mult_21_C243_n757);
   mult_21_C243_U1274 : MUXB2DL port map( A0 => N3107, A1 => N3108, SL => 
                           mult_21_C243_n1442, Z => mult_21_C243_n758);
   mult_21_C243_U1273 : MUXB2DL port map( A0 => N3106, A1 => N3107, SL => 
                           mult_21_C243_n1442, Z => mult_21_C243_n759);
   mult_21_C243_U1272 : MUXB2DL port map( A0 => N3105, A1 => N3106, SL => 
                           mult_21_C243_n1442, Z => mult_21_C243_n760);
   mult_21_C243_U1271 : NAN2D1 port map( A1 => N3105, A2 => mult_21_C243_n1442,
                           Z => mult_21_C243_n761);
   mult_21_C243_U1270 : MUXB2DL port map( A0 => N3125, A1 => N3126, SL => 
                           mult_21_C243_n1441, Z => mult_21_C243_n762);
   mult_21_C243_U1269 : MUXB2DL port map( A0 => N3124, A1 => N3125, SL => 
                           mult_21_C243_n1441, Z => mult_21_C243_n763);
   mult_21_C243_U1268 : MUXB2DL port map( A0 => N3123, A1 => N3124, SL => 
                           mult_21_C243_n1441, Z => mult_21_C243_n764);
   mult_21_C243_U1267 : MUXB2DL port map( A0 => N3122, A1 => N3123, SL => 
                           mult_21_C243_n1441, Z => mult_21_C243_n765);
   mult_21_C243_U1266 : MUXB2DL port map( A0 => N3121, A1 => N3122, SL => 
                           mult_21_C243_n1441, Z => mult_21_C243_n766);
   mult_21_C243_U1265 : MUXB2DL port map( A0 => N3120, A1 => N3121, SL => 
                           mult_21_C243_n1441, Z => mult_21_C243_n767);
   mult_21_C243_U1264 : MUXB2DL port map( A0 => N3119, A1 => N3120, SL => 
                           mult_21_C243_n1441, Z => mult_21_C243_n768);
   mult_21_C243_U1263 : MUXB2DL port map( A0 => N3118, A1 => N3119, SL => 
                           mult_21_C243_n1441, Z => mult_21_C243_n769);
   mult_21_C243_U1262 : MUXB2DL port map( A0 => N3117, A1 => N3118, SL => 
                           mult_21_C243_n1441, Z => mult_21_C243_n770);
   mult_21_C243_U1261 : MUXB2DL port map( A0 => N3116, A1 => N3117, SL => 
                           mult_21_C243_n1441, Z => mult_21_C243_n771);
   mult_21_C243_U1260 : MUXB2DL port map( A0 => N3115, A1 => N3116, SL => 
                           mult_21_C243_n1441, Z => mult_21_C243_n772);
   mult_21_C243_U1259 : MUXB2DL port map( A0 => N3114, A1 => N3115, SL => 
                           mult_21_C243_n1441, Z => mult_21_C243_n773);
   mult_21_C243_U1258 : MUXB2DL port map( A0 => N3113, A1 => N3114, SL => 
                           mult_21_C243_n1441, Z => mult_21_C243_n774);
   mult_21_C243_U1257 : MUXB2DL port map( A0 => N3112, A1 => N3113, SL => 
                           mult_21_C243_n1441, Z => mult_21_C243_n775);
   mult_21_C243_U1256 : MUXB2DL port map( A0 => N3111, A1 => N3112, SL => 
                           mult_21_C243_n1441, Z => mult_21_C243_n776);
   mult_21_C243_U1255 : MUXB2DL port map( A0 => N3110, A1 => N3111, SL => 
                           mult_21_C243_n1441, Z => mult_21_C243_n777);
   mult_21_C243_U1254 : MUXB2DL port map( A0 => N3109, A1 => N3110, SL => 
                           mult_21_C243_n1441, Z => mult_21_C243_n778);
   mult_21_C243_U1253 : MUXB2DL port map( A0 => N3108, A1 => N3109, SL => 
                           mult_21_C243_n1441, Z => mult_21_C243_n779);
   mult_21_C243_U1252 : MUXB2DL port map( A0 => N3107, A1 => N3108, SL => 
                           mult_21_C243_n1441, Z => mult_21_C243_n780);
   mult_21_C243_U1251 : MUXB2DL port map( A0 => mult_21_C243_n1388, A1 => N3107
                           , SL => mult_21_C243_n1441, Z => mult_21_C243_n781);
   mult_21_C243_U1250 : MUXB2DL port map( A0 => N3105, A1 => N3106, SL => 
                           mult_21_C243_n1441, Z => mult_21_C243_n782);
   mult_21_C243_U1249 : NAN2D1 port map( A1 => N3105, A2 => mult_21_C243_n1441,
                           Z => mult_21_C243_n783);
   mult_21_C243_U1248 : MUXB2DL port map( A0 => N3127, A1 => N3128, SL => 
                           mult_21_C243_n1379, Z => mult_21_C243_n784);
   mult_21_C243_U1247 : MUXB2DL port map( A0 => N3126, A1 => N3127, SL => 
                           mult_21_C243_n1379, Z => mult_21_C243_n785);
   mult_21_C243_U1246 : MUXB2DL port map( A0 => N3125, A1 => N3126, SL => 
                           mult_21_C243_n1379, Z => mult_21_C243_n786);
   mult_21_C243_U1245 : MUXB2DL port map( A0 => N3124, A1 => N3125, SL => 
                           mult_21_C243_n1379, Z => mult_21_C243_n787);
   mult_21_C243_U1244 : MUXB2DL port map( A0 => N3123, A1 => N3124, SL => 
                           mult_21_C243_n1379, Z => mult_21_C243_n788);
   mult_21_C243_U1243 : MUXB2DL port map( A0 => N3122, A1 => N3123, SL => 
                           mult_21_C243_n1379, Z => mult_21_C243_n789);
   mult_21_C243_U1242 : MUXB2DL port map( A0 => N3121, A1 => N3122, SL => 
                           mult_21_C243_n1379, Z => mult_21_C243_n790);
   mult_21_C243_U1241 : MUXB2DL port map( A0 => N3120, A1 => N3121, SL => 
                           mult_21_C243_n1379, Z => mult_21_C243_n791);
   mult_21_C243_U1240 : MUXB2DL port map( A0 => N3119, A1 => N3120, SL => 
                           mult_21_C243_n1379, Z => mult_21_C243_n792);
   mult_21_C243_U1239 : MUXB2DL port map( A0 => N3118, A1 => N3119, SL => 
                           mult_21_C243_n1379, Z => mult_21_C243_n793);
   mult_21_C243_U1238 : MUXB2DL port map( A0 => N3117, A1 => N3118, SL => 
                           mult_21_C243_n1379, Z => mult_21_C243_n794);
   mult_21_C243_U1237 : MUXB2DL port map( A0 => N3116, A1 => N3117, SL => 
                           mult_21_C243_n1379, Z => mult_21_C243_n795);
   mult_21_C243_U1236 : MUXB2DL port map( A0 => N3115, A1 => N3116, SL => 
                           mult_21_C243_n1379, Z => mult_21_C243_n796);
   mult_21_C243_U1235 : MUXB2DL port map( A0 => N3114, A1 => N3115, SL => 
                           mult_21_C243_n1379, Z => mult_21_C243_n797);
   mult_21_C243_U1234 : MUXB2DL port map( A0 => N3113, A1 => N3114, SL => 
                           mult_21_C243_n1379, Z => mult_21_C243_n798);
   mult_21_C243_U1233 : MUXB2DL port map( A0 => N3112, A1 => N3113, SL => 
                           mult_21_C243_n1379, Z => mult_21_C243_n799);
   mult_21_C243_U1232 : MUXB2DL port map( A0 => N3111, A1 => N3112, SL => 
                           mult_21_C243_n1379, Z => mult_21_C243_n800);
   mult_21_C243_U1231 : MUXB2DL port map( A0 => N3110, A1 => N3111, SL => 
                           mult_21_C243_n1379, Z => mult_21_C243_n801);
   mult_21_C243_U1230 : MUXB2DL port map( A0 => N3109, A1 => N3110, SL => 
                           mult_21_C243_n1379, Z => mult_21_C243_n802);
   mult_21_C243_U1229 : MUXB2DL port map( A0 => mult_21_C243_n1386, A1 => N3109
                           , SL => mult_21_C243_n1379, Z => mult_21_C243_n803);
   mult_21_C243_U1228 : MUXB2DL port map( A0 => N3107, A1 => N3108, SL => 
                           mult_21_C243_n1379, Z => mult_21_C243_n804);
   mult_21_C243_U1227 : MUXB2DL port map( A0 => N3106, A1 => N3107, SL => 
                           mult_21_C243_n1379, Z => mult_21_C243_n805);
   mult_21_C243_U1226 : MUXB2DL port map( A0 => N3105, A1 => N3106, SL => 
                           mult_21_C243_n1379, Z => mult_21_C243_n806);
   mult_21_C243_U1225 : NAN2D1 port map( A1 => N3105, A2 => mult_21_C243_n1379,
                           Z => mult_21_C243_n807);
   mult_21_C243_U1224 : MUXB2DL port map( A0 => N3129, A1 => N3130, SL => 
                           mult_21_C243_n1378, Z => mult_21_C243_n808);
   mult_21_C243_U1223 : MUXB2DL port map( A0 => N3128, A1 => N3129, SL => 
                           mult_21_C243_n1378, Z => mult_21_C243_n809);
   mult_21_C243_U1222 : AOI21D1 port map( A1 => N2964, A2 => N2965, B => 
                           mult_21_C243_n1413, Z => mult_21_C243_n944);
   mult_21_C243_U1221 : MUXB2DL port map( A0 => N3127, A1 => N3128, SL => 
                           mult_21_C243_n1378, Z => mult_21_C243_n810);
   mult_21_C243_U1220 : MUXB2DL port map( A0 => N3126, A1 => N3127, SL => 
                           mult_21_C243_n1378, Z => mult_21_C243_n811);
   mult_21_C243_U1219 : MUXB2DL port map( A0 => N3125, A1 => N3126, SL => 
                           mult_21_C243_n1378, Z => mult_21_C243_n812);
   mult_21_C243_U1218 : MUXB2DL port map( A0 => N3124, A1 => N3125, SL => 
                           mult_21_C243_n1378, Z => mult_21_C243_n813);
   mult_21_C243_U1217 : MUXB2DL port map( A0 => N3123, A1 => N3124, SL => 
                           mult_21_C243_n1378, Z => mult_21_C243_n814);
   mult_21_C243_U1216 : MUXB2DL port map( A0 => N3122, A1 => N3123, SL => 
                           mult_21_C243_n1378, Z => mult_21_C243_n815);
   mult_21_C243_U1215 : MUXB2DL port map( A0 => N3121, A1 => N3122, SL => 
                           mult_21_C243_n1378, Z => mult_21_C243_n816);
   mult_21_C243_U1214 : MUXB2DL port map( A0 => N3120, A1 => N3121, SL => 
                           mult_21_C243_n1378, Z => mult_21_C243_n817);
   mult_21_C243_U1213 : MUXB2DL port map( A0 => N3119, A1 => N3120, SL => 
                           mult_21_C243_n1378, Z => mult_21_C243_n818);
   mult_21_C243_U1212 : MUXB2DL port map( A0 => N3118, A1 => N3119, SL => 
                           mult_21_C243_n1378, Z => mult_21_C243_n819);
   mult_21_C243_U1211 : MUXB2DL port map( A0 => N3117, A1 => N3118, SL => 
                           mult_21_C243_n1378, Z => mult_21_C243_n820);
   mult_21_C243_U1210 : MUXB2DL port map( A0 => N3116, A1 => N3117, SL => 
                           mult_21_C243_n1378, Z => mult_21_C243_n821);
   mult_21_C243_U1209 : MUXB2DL port map( A0 => N3115, A1 => N3116, SL => 
                           mult_21_C243_n1378, Z => mult_21_C243_n822);
   mult_21_C243_U1208 : MUXB2DL port map( A0 => N3114, A1 => N3115, SL => 
                           mult_21_C243_n1378, Z => mult_21_C243_n823);
   mult_21_C243_U1207 : MUXB2DL port map( A0 => N3113, A1 => N3114, SL => 
                           mult_21_C243_n1378, Z => mult_21_C243_n824);
   mult_21_C243_U1206 : MUXB2DL port map( A0 => N3112, A1 => N3113, SL => 
                           mult_21_C243_n1378, Z => mult_21_C243_n825);
   mult_21_C243_U1205 : MUXB2DL port map( A0 => N3111, A1 => N3112, SL => 
                           mult_21_C243_n1378, Z => mult_21_C243_n826);
   mult_21_C243_U1204 : MUXB2DL port map( A0 => N3110, A1 => N3111, SL => 
                           mult_21_C243_n1378, Z => mult_21_C243_n827);
   mult_21_C243_U1203 : MUXB2DL port map( A0 => N3109, A1 => N3110, SL => 
                           mult_21_C243_n1378, Z => mult_21_C243_n828);
   mult_21_C243_U1202 : MUXB2DL port map( A0 => mult_21_C243_n1386, A1 => N3109
                           , SL => mult_21_C243_n1378, Z => mult_21_C243_n829);
   mult_21_C243_U1201 : MUXB2DL port map( A0 => N3107, A1 => N3108, SL => 
                           mult_21_C243_n1378, Z => mult_21_C243_n830);
   mult_21_C243_U1200 : MUXB2DL port map( A0 => mult_21_C243_n1388, A1 => N3107
                           , SL => mult_21_C243_n1378, Z => mult_21_C243_n831);
   mult_21_C243_U1199 : MUXB2DL port map( A0 => N3105, A1 => N3106, SL => 
                           mult_21_C243_n1378, Z => mult_21_C243_n832);
   mult_21_C243_U1198 : NAN2D1 port map( A1 => N3105, A2 => mult_21_C243_n1378,
                           Z => mult_21_C243_n833);
   mult_21_C243_U1197 : MUXB2DL port map( A0 => N3131, A1 => N3132, SL => 
                           mult_21_C243_n1385, Z => mult_21_C243_n834);
   mult_21_C243_U1196 : MUXB2DL port map( A0 => N3130, A1 => N3131, SL => 
                           mult_21_C243_n1385, Z => mult_21_C243_n835);
   mult_21_C243_U1195 : MUXB2DL port map( A0 => N3129, A1 => N3130, SL => 
                           mult_21_C243_n1385, Z => mult_21_C243_n836);
   mult_21_C243_U1194 : MUXB2DL port map( A0 => N3128, A1 => N3129, SL => 
                           mult_21_C243_n1385, Z => mult_21_C243_n837);
   mult_21_C243_U1193 : MUXB2DL port map( A0 => N3127, A1 => N3128, SL => 
                           mult_21_C243_n1385, Z => mult_21_C243_n838);
   mult_21_C243_U1192 : MUXB2DL port map( A0 => N3126, A1 => N3127, SL => 
                           mult_21_C243_n1385, Z => mult_21_C243_n839);
   mult_21_C243_U1191 : MUXB2DL port map( A0 => N3125, A1 => N3126, SL => 
                           mult_21_C243_n1385, Z => mult_21_C243_n840);
   mult_21_C243_U1190 : MUXB2DL port map( A0 => N3124, A1 => N3125, SL => 
                           mult_21_C243_n1385, Z => mult_21_C243_n841);
   mult_21_C243_U1189 : MUXB2DL port map( A0 => N3123, A1 => N3124, SL => 
                           mult_21_C243_n1385, Z => mult_21_C243_n842);
   mult_21_C243_U1188 : MUXB2DL port map( A0 => N3122, A1 => N3123, SL => 
                           mult_21_C243_n1385, Z => mult_21_C243_n843);
   mult_21_C243_U1187 : MUXB2DL port map( A0 => N3121, A1 => N3122, SL => 
                           mult_21_C243_n1385, Z => mult_21_C243_n844);
   mult_21_C243_U1186 : MUXB2DL port map( A0 => N3120, A1 => N3121, SL => 
                           mult_21_C243_n1385, Z => mult_21_C243_n845);
   mult_21_C243_U1185 : MUXB2DL port map( A0 => N3119, A1 => N3120, SL => 
                           mult_21_C243_n1385, Z => mult_21_C243_n846);
   mult_21_C243_U1184 : MUXB2DL port map( A0 => N3118, A1 => N3119, SL => 
                           mult_21_C243_n1385, Z => mult_21_C243_n847);
   mult_21_C243_U1183 : MUXB2DL port map( A0 => N3117, A1 => N3118, SL => 
                           mult_21_C243_n1385, Z => mult_21_C243_n848);
   mult_21_C243_U1182 : MUXB2DL port map( A0 => N3116, A1 => N3117, SL => 
                           mult_21_C243_n1385, Z => mult_21_C243_n849);
   mult_21_C243_U1181 : MUXB2DL port map( A0 => N3115, A1 => N3116, SL => 
                           mult_21_C243_n1385, Z => mult_21_C243_n850);
   mult_21_C243_U1180 : MUXB2DL port map( A0 => N3114, A1 => N3115, SL => 
                           mult_21_C243_n1385, Z => mult_21_C243_n851);
   mult_21_C243_U1179 : MUXB2DL port map( A0 => N3113, A1 => N3114, SL => 
                           mult_21_C243_n1385, Z => mult_21_C243_n852);
   mult_21_C243_U1178 : MUXB2DL port map( A0 => N3112, A1 => N3113, SL => 
                           mult_21_C243_n1385, Z => mult_21_C243_n853);
   mult_21_C243_U1177 : MUXB2DL port map( A0 => N3111, A1 => N3112, SL => 
                           mult_21_C243_n1385, Z => mult_21_C243_n854);
   mult_21_C243_U1176 : MUXB2DL port map( A0 => N3110, A1 => N3111, SL => 
                           mult_21_C243_n1385, Z => mult_21_C243_n855);
   mult_21_C243_U1175 : MUXB2DL port map( A0 => N3109, A1 => N3110, SL => 
                           mult_21_C243_n1385, Z => mult_21_C243_n856);
   mult_21_C243_U1174 : MUXB2DL port map( A0 => mult_21_C243_n1386, A1 => N3109
                           , SL => mult_21_C243_n1385, Z => mult_21_C243_n857);
   mult_21_C243_U1173 : MUXB2DL port map( A0 => N3107, A1 => N3108, SL => 
                           mult_21_C243_n1385, Z => mult_21_C243_n858);
   mult_21_C243_U1172 : MUXB2DL port map( A0 => mult_21_C243_n1388, A1 => N3107
                           , SL => mult_21_C243_n1385, Z => mult_21_C243_n859);
   mult_21_C243_U1171 : AOI21D1 port map( A1 => N2966, A2 => N2967, B => 
                           mult_21_C243_n1415, Z => mult_21_C243_n943);
   mult_21_C243_U1170 : MUXB2DL port map( A0 => N3105, A1 => N3106, SL => 
                           mult_21_C243_n1385, Z => mult_21_C243_n860);
   mult_21_C243_U1169 : NAN2D1 port map( A1 => N3105, A2 => mult_21_C243_n1385,
                           Z => mult_21_C243_n861);
   mult_21_C243_U1168 : MUXB2DL port map( A0 => N3132, A1 => N3133, SL => 
                           mult_21_C243_n1384, Z => mult_21_C243_n863);
   mult_21_C243_U1167 : MUXB2DL port map( A0 => N3131, A1 => N3132, SL => 
                           mult_21_C243_n1384, Z => mult_21_C243_n864);
   mult_21_C243_U1166 : MUXB2DL port map( A0 => N3130, A1 => N3131, SL => 
                           mult_21_C243_n1384, Z => mult_21_C243_n865);
   mult_21_C243_U1165 : MUXB2DL port map( A0 => N3129, A1 => N3130, SL => 
                           mult_21_C243_n1384, Z => mult_21_C243_n866);
   mult_21_C243_U1164 : MUXB2DL port map( A0 => N3128, A1 => N3129, SL => 
                           mult_21_C243_n1384, Z => mult_21_C243_n867);
   mult_21_C243_U1163 : MUXB2DL port map( A0 => N3127, A1 => N3128, SL => 
                           mult_21_C243_n1384, Z => mult_21_C243_n868);
   mult_21_C243_U1162 : MUXB2DL port map( A0 => N3126, A1 => N3127, SL => 
                           mult_21_C243_n1384, Z => mult_21_C243_n869);
   mult_21_C243_U1161 : MUXB2DL port map( A0 => N3125, A1 => N3126, SL => 
                           mult_21_C243_n1384, Z => mult_21_C243_n870);
   mult_21_C243_U1160 : MUXB2DL port map( A0 => N3124, A1 => N3125, SL => 
                           mult_21_C243_n1384, Z => mult_21_C243_n871);
   mult_21_C243_U1159 : MUXB2DL port map( A0 => N3123, A1 => N3124, SL => 
                           mult_21_C243_n1384, Z => mult_21_C243_n872);
   mult_21_C243_U1158 : MUXB2DL port map( A0 => N3122, A1 => N3123, SL => 
                           mult_21_C243_n1384, Z => mult_21_C243_n873);
   mult_21_C243_U1157 : MUXB2DL port map( A0 => N3121, A1 => N3122, SL => 
                           mult_21_C243_n1384, Z => mult_21_C243_n874);
   mult_21_C243_U1156 : MUXB2DL port map( A0 => N3120, A1 => N3121, SL => 
                           mult_21_C243_n1384, Z => mult_21_C243_n875);
   mult_21_C243_U1155 : MUXB2DL port map( A0 => N3119, A1 => N3120, SL => 
                           mult_21_C243_n1384, Z => mult_21_C243_n876);
   mult_21_C243_U1154 : MUXB2DL port map( A0 => N3118, A1 => N3119, SL => 
                           mult_21_C243_n1384, Z => mult_21_C243_n877);
   mult_21_C243_U1153 : MUXB2DL port map( A0 => N3117, A1 => N3118, SL => 
                           mult_21_C243_n1384, Z => mult_21_C243_n878);
   mult_21_C243_U1152 : MUXB2DL port map( A0 => N3116, A1 => N3117, SL => 
                           mult_21_C243_n1384, Z => mult_21_C243_n879);
   mult_21_C243_U1151 : MUXB2DL port map( A0 => N3115, A1 => N3116, SL => 
                           mult_21_C243_n1384, Z => mult_21_C243_n880);
   mult_21_C243_U1150 : MUXB2DL port map( A0 => N3114, A1 => N3115, SL => 
                           mult_21_C243_n1384, Z => mult_21_C243_n881);
   mult_21_C243_U1149 : MUXB2DL port map( A0 => N3113, A1 => N3114, SL => 
                           mult_21_C243_n1384, Z => mult_21_C243_n882);
   mult_21_C243_U1148 : MUXB2DL port map( A0 => N3112, A1 => N3113, SL => 
                           mult_21_C243_n1384, Z => mult_21_C243_n883);
   mult_21_C243_U1147 : MUXB2DL port map( A0 => N3111, A1 => N3112, SL => 
                           mult_21_C243_n1384, Z => mult_21_C243_n884);
   mult_21_C243_U1146 : MUXB2DL port map( A0 => N3110, A1 => N3111, SL => 
                           mult_21_C243_n1384, Z => mult_21_C243_n885);
   mult_21_C243_U1145 : MUXB2DL port map( A0 => N3109, A1 => N3110, SL => 
                           mult_21_C243_n1384, Z => mult_21_C243_n886);
   mult_21_C243_U1144 : MUXB2DL port map( A0 => mult_21_C243_n1386, A1 => N3109
                           , SL => mult_21_C243_n1384, Z => mult_21_C243_n887);
   mult_21_C243_U1143 : MUXB2DL port map( A0 => N3107, A1 => N3108, SL => 
                           mult_21_C243_n1384, Z => mult_21_C243_n888);
   mult_21_C243_U1142 : MUXB2DL port map( A0 => mult_21_C243_n1388, A1 => N3107
                           , SL => mult_21_C243_n1384, Z => mult_21_C243_n889);
   mult_21_C243_U1141 : OAI21D1 port map( A1 => N2969, A2 => N2968, B => 
                           mult_21_C243_n1417, Z => mult_21_C243_n89);
   mult_21_C243_U1140 : MUXB2DL port map( A0 => N3105, A1 => N3106, SL => 
                           mult_21_C243_n1384, Z => mult_21_C243_n890);
   mult_21_C243_U1139 : NAN2D1 port map( A1 => N3105, A2 => mult_21_C243_n1384,
                           Z => mult_21_C243_n891);
   mult_21_C243_U1138 : MUXB2DL port map( A0 => N3135, A1 => N3136, SL => 
                           mult_21_C243_n1390, Z => mult_21_C243_n892);
   mult_21_C243_U1137 : MUXB2DL port map( A0 => N3134, A1 => N3135, SL => N2945
                           , Z => mult_21_C243_n893);
   mult_21_C243_U1136 : MUXB2DL port map( A0 => N3133, A1 => N3134, SL => N2945
                           , Z => mult_21_C243_n894);
   mult_21_C243_U1135 : MUXB2DL port map( A0 => N3132, A1 => N3133, SL => N2945
                           , Z => mult_21_C243_n895);
   mult_21_C243_U1134 : MUXB2DL port map( A0 => N3131, A1 => N3132, SL => N2945
                           , Z => mult_21_C243_n896);
   mult_21_C243_U1133 : MUXB2DL port map( A0 => N3130, A1 => N3131, SL => N2945
                           , Z => mult_21_C243_n897);
   mult_21_C243_U1132 : MUXB2DL port map( A0 => N3129, A1 => N3130, SL => N2945
                           , Z => mult_21_C243_n898);
   mult_21_C243_U1131 : MUXB2DL port map( A0 => N3128, A1 => N3129, SL => N2945
                           , Z => mult_21_C243_n899);
   mult_21_C243_U1130 : MUXB2DL port map( A0 => N3127, A1 => N3128, SL => N2945
                           , Z => mult_21_C243_n900);
   mult_21_C243_U1129 : MUXB2DL port map( A0 => N3126, A1 => N3127, SL => N2945
                           , Z => mult_21_C243_n901);
   mult_21_C243_U1128 : MUXB2DL port map( A0 => N3125, A1 => N3126, SL => N2945
                           , Z => mult_21_C243_n902);
   mult_21_C243_U1127 : MUXB2DL port map( A0 => N3124, A1 => N3125, SL => N2945
                           , Z => mult_21_C243_n903);
   mult_21_C243_U1126 : MUXB2DL port map( A0 => N3123, A1 => N3124, SL => N2945
                           , Z => mult_21_C243_n904);
   mult_21_C243_U1125 : MUXB2DL port map( A0 => N3122, A1 => N3123, SL => N2945
                           , Z => mult_21_C243_n905);
   mult_21_C243_U1124 : MUXB2DL port map( A0 => N3121, A1 => N3122, SL => N2945
                           , Z => mult_21_C243_n906);
   mult_21_C243_U1123 : MUXB2DL port map( A0 => N3120, A1 => N3121, SL => N2945
                           , Z => mult_21_C243_n907);
   mult_21_C243_U1122 : MUXB2DL port map( A0 => N3119, A1 => N3120, SL => N2945
                           , Z => mult_21_C243_n908);
   mult_21_C243_U1121 : MUXB2DL port map( A0 => N3118, A1 => N3119, SL => N2945
                           , Z => mult_21_C243_n909);
   mult_21_C243_U1120 : AOI21D1 port map( A1 => N2968, A2 => N2969, B => 
                           mult_21_C243_n1417, Z => mult_21_C243_n942);
   mult_21_C243_U1119 : MUXB2DL port map( A0 => N3117, A1 => N3118, SL => 
                           mult_21_C243_n1390, Z => mult_21_C243_n910);
   mult_21_C243_U1118 : MUXB2DL port map( A0 => N3116, A1 => N3117, SL => 
                           mult_21_C243_n1390, Z => mult_21_C243_n911);
   mult_21_C243_U1117 : MUXB2DL port map( A0 => N3115, A1 => N3116, SL => 
                           mult_21_C243_n1390, Z => mult_21_C243_n912);
   mult_21_C243_U1116 : MUXB2DL port map( A0 => N3114, A1 => N3115, SL => 
                           mult_21_C243_n1390, Z => mult_21_C243_n913);
   mult_21_C243_U1115 : MUXB2DL port map( A0 => N3113, A1 => N3114, SL => 
                           mult_21_C243_n1390, Z => mult_21_C243_n914);
   mult_21_C243_U1114 : MUXB2DL port map( A0 => N3112, A1 => N3113, SL => 
                           mult_21_C243_n1390, Z => mult_21_C243_n915);
   mult_21_C243_U1113 : MUXB2DL port map( A0 => N3111, A1 => N3112, SL => 
                           mult_21_C243_n1390, Z => mult_21_C243_n916);
   mult_21_C243_U1112 : MUXB2DL port map( A0 => N3110, A1 => N3111, SL => 
                           mult_21_C243_n1390, Z => mult_21_C243_n917);
   mult_21_C243_U1111 : MUXB2DL port map( A0 => N3109, A1 => N3110, SL => 
                           mult_21_C243_n1390, Z => mult_21_C243_n918);
   mult_21_C243_U1110 : MUXB2DL port map( A0 => mult_21_C243_n1386, A1 => N3109
                           , SL => mult_21_C243_n1390, Z => mult_21_C243_n919);
   mult_21_C243_U1109 : MUXB2DL port map( A0 => N3107, A1 => mult_21_C243_n1386
                           , SL => mult_21_C243_n1390, Z => mult_21_C243_n920);
   mult_21_C243_U1108 : MUXB2DL port map( A0 => mult_21_C243_n1388, A1 => N3107
                           , SL => mult_21_C243_n1390, Z => mult_21_C243_n921);
   mult_21_C243_U1107 : MUXB2DL port map( A0 => N3105, A1 => mult_21_C243_n1388
                           , SL => mult_21_C243_n1390, Z => mult_21_C243_n922);
   mult_21_C243_U1106 : NAN2D1 port map( A1 => N3105, A2 => mult_21_C243_n1390,
                           Z => mult_21_C243_n923);
   mult_21_C243_U1105 : OAI21D1 port map( A1 => N2971, A2 => N2970, B => 
                           mult_21_C243_n1418, Z => mult_21_C243_n94);
   mult_21_C243_U1104 : AOI21D1 port map( A1 => N2970, A2 => N2971, B => 
                           mult_21_C243_n1418, Z => mult_21_C243_n941);
   mult_21_C243_U1103 : OAI21D1 port map( A1 => N2973, A2 => N2972, B => 
                           mult_21_C243_n1421, Z => mult_21_C243_n99);
   mult_21_C243_U1102 : EXOR2D1 port map( A1 => mult_21_C243_n230, A2 => 
                           mult_21_C243_n228, Z => mult_21_C243_n1440);
   mult_21_C243_U1101 : EXOR3D1 port map( A1 => mult_21_C243_n226, A2 => 
                           mult_21_C243_n224, A3 => mult_21_C243_n1440, Z => 
                           mult_21_C243_n1435);
   mult_21_C243_U1100 : EXOR2D1 port map( A1 => mult_21_C243_n222, A2 => 
                           mult_21_C243_n220, Z => mult_21_C243_n1439);
   mult_21_C243_U1099 : EXOR3D1 port map( A1 => mult_21_C243_n216, A2 => 
                           mult_21_C243_n1195, A3 => mult_21_C243_n1439, Z => 
                           mult_21_C243_n1436);
   mult_21_C243_U1098 : EXOR3D1 port map( A1 => mult_21_C243_n1165, A2 => 
                           mult_21_C243_n1137, A3 => mult_21_C243_n1045, Z => 
                           mult_21_C243_n1438);
   mult_21_C243_U1097 : EXOR3D1 port map( A1 => mult_21_C243_n1027, A2 => 
                           mult_21_C243_n1011, A3 => mult_21_C243_n1438, Z => 
                           mult_21_C243_n1437);
   mult_21_C243_U1096 : EXOR3D1 port map( A1 => mult_21_C243_n1435, A2 => 
                           mult_21_C243_n1436, A3 => mult_21_C243_n1437, Z => 
                           mult_21_C243_n1427);
   mult_21_C243_U1095 : EXOR2D1 port map( A1 => mult_21_C243_n985, A2 => 
                           mult_21_C243_n967, Z => mult_21_C243_n1434);
   mult_21_C243_U1094 : EXOR3D1 port map( A1 => mult_21_C243_n961, A2 => 
                           mult_21_C243_n218, A3 => mult_21_C243_n1434, Z => 
                           mult_21_C243_n1431);
   mult_21_C243_U1093 : EXNOR2D1 port map( A1 => mult_21_C243_n210, A2 => 
                           mult_21_C243_n1111, Z => mult_21_C243_n1433);
   mult_21_C243_U1092 : EXOR3D1 port map( A1 => mult_21_C243_n1087, A2 => 
                           mult_21_C243_n1065, A3 => mult_21_C243_n1433, Z => 
                           mult_21_C243_n1432);
   mult_21_C243_U1091 : EXOR3D1 port map( A1 => mult_21_C243_n1431, A2 => 
                           mult_21_C243_n204, A3 => mult_21_C243_n1432, Z => 
                           mult_21_C243_n1428);
   mult_21_C243_U1090 : EXNOR2D1 port map( A1 => mult_21_C243_n997, A2 => 
                           mult_21_C243_n975, Z => mult_21_C243_n1430);
   mult_21_C243_U1089 : EXOR3D1 port map( A1 => mult_21_C243_n957, A2 => 
                           mult_21_C243_n955, A3 => mult_21_C243_n1430, Z => 
                           mult_21_C243_n1429);
   mult_21_C243_U1088 : EXOR3D1 port map( A1 => mult_21_C243_n1427, A2 => 
                           mult_21_C243_n1428, A3 => mult_21_C243_n1429, Z => 
                           mult_21_C243_n1423);
   mult_21_C243_U1087 : EXOR2D1 port map( A1 => mult_21_C243_n202, A2 => 
                           mult_21_C243_n156, Z => mult_21_C243_n1424);
   mult_21_C243_U1086 : EXOR2D1 port map( A1 => mult_21_C243_n214, A2 => 
                           mult_21_C243_n212, Z => mult_21_C243_n1426);
   mult_21_C243_U1085 : EXOR3D1 port map( A1 => mult_21_C243_n208, A2 => 
                           mult_21_C243_n206, A3 => mult_21_C243_n1426, Z => 
                           mult_21_C243_n1425);
   mult_21_C243_U1084 : EXOR3D1 port map( A1 => mult_21_C243_n1423, A2 => 
                           mult_21_C243_n1424, A3 => mult_21_C243_n1425, Z => 
                           N3296);
   mult_21_C243_U1083 : INVD1 port map( A => N2976, Z => mult_21_C243_n1422);
   mult_21_C243_U1082 : INVD1 port map( A => N3108, Z => mult_21_C243_n1387);
   mult_21_C243_U1081 : INVD1 port map( A => N3106, Z => mult_21_C243_n1389);
   mult_21_C243_U1080 : INVD1 port map( A => N2945, Z => mult_21_C243_n1391);
   mult_21_C243_U1079 : MUXB2DL port map( A0 => N3134, A1 => N3133, SL => 
                           mult_21_C243_n1382, Z => mult_21_C243_n862);
   mult_21_C243_U1078 : INVD1 port map( A => N2974, Z => mult_21_C243_n1421);
   mult_21_C243_U1077 : INVD1 port map( A => N2972, Z => mult_21_C243_n1418);
   mult_21_C243_U1076 : INVD1 port map( A => N2970, Z => mult_21_C243_n1417);
   mult_21_C243_U1075 : OAI21D1 port map( A1 => N2967, A2 => N2966, B => 
                           mult_21_C243_n1415, Z => mult_21_C243_n84);
   mult_21_C243_U1074 : INVD1 port map( A => N2968, Z => mult_21_C243_n1415);
   mult_21_C243_U1073 : EXOR2D1 port map( A1 => N2967, A2 => N2966, Z => 
                           mult_21_C243_n1447);
   mult_21_C243_U1072 : OAI21D1 port map( A1 => N2965, A2 => N2964, B => 
                           mult_21_C243_n1413, Z => mult_21_C243_n80);
   mult_21_C243_U1071 : INVD1 port map( A => N2966, Z => mult_21_C243_n1413);
   mult_21_C243_U1070 : EXOR2D1 port map( A1 => N2965, A2 => N2964, Z => 
                           mult_21_C243_n1446);
   mult_21_C243_U1069 : OAI21D1 port map( A1 => N2963, A2 => N2962, B => 
                           mult_21_C243_n1411, Z => mult_21_C243_n73);
   mult_21_C243_U1068 : INVD1 port map( A => N2964, Z => mult_21_C243_n1411);
   mult_21_C243_U1067 : EXOR2D1 port map( A1 => N2963, A2 => N2962, Z => 
                           mult_21_C243_n1445);
   mult_21_C243_U1066 : OAI21D1 port map( A1 => N2961, A2 => N2960, B => 
                           mult_21_C243_n1409, Z => mult_21_C243_n66);
   mult_21_C243_U1065 : INVD1 port map( A => N2962, Z => mult_21_C243_n1409);
   mult_21_C243_U1064 : EXOR2D1 port map( A1 => N2961, A2 => N2960, Z => 
                           mult_21_C243_n1444);
   mult_21_C243_U1063 : OAI21D1 port map( A1 => N2959, A2 => N2958, B => 
                           mult_21_C243_n1407, Z => mult_21_C243_n58);
   mult_21_C243_U1062 : INVD1 port map( A => N2960, Z => mult_21_C243_n1407);
   mult_21_C243_U1061 : EXOR2D1 port map( A1 => N2959, A2 => N2958, Z => 
                           mult_21_C243_n1443);
   mult_21_C243_U1060 : OAI21D1 port map( A1 => N2957, A2 => N2956, B => 
                           mult_21_C243_n1405, Z => mult_21_C243_n50);
   mult_21_C243_U1059 : INVD1 port map( A => N2958, Z => mult_21_C243_n1405);
   mult_21_C243_U1058 : EXOR2D1 port map( A1 => N2957, A2 => N2956, Z => 
                           mult_21_C243_n1442);
   mult_21_C243_U1057 : OAI21D1 port map( A1 => N2954, A2 => N2955, B => 
                           mult_21_C243_n1403, Z => mult_21_C243_n42);
   mult_21_C243_U1056 : INVD1 port map( A => N2956, Z => mult_21_C243_n1403);
   mult_21_C243_U1055 : EXOR2D1 port map( A1 => N2955, A2 => N2954, Z => 
                           mult_21_C243_n1441);
   mult_21_C243_U1054 : INVD1 port map( A => N2954, Z => mult_21_C243_n1401);
   mult_21_C243_U1053 : INVD1 port map( A => N2952, Z => mult_21_C243_n1399);
   mult_21_C243_U1052 : INVD1 port map( A => N2950, Z => mult_21_C243_n1397);
   mult_21_C243_U1051 : INVD1 port map( A => N2948, Z => mult_21_C243_n1395);
   mult_21_C243_U1050 : INVD1 port map( A => mult_21_C243_n1387, Z => 
                           mult_21_C243_n1386);
   mult_21_C243_U1049 : EXNOR2D1 port map( A1 => N2949, A2 => N2948, Z => 
                           mult_21_C243_n1383);
   mult_21_C243_U1048 : INVD1 port map( A => mult_21_C243_n1389, Z => 
                           mult_21_C243_n1388);
   mult_21_C243_U1047 : EXNOR2D1 port map( A1 => N2947, A2 => N2946, Z => 
                           mult_21_C243_n1382);
   mult_21_C243_U1046 : INVD1 port map( A => N2946, Z => mult_21_C243_n1392);
   mult_21_C243_U1045 : INVD1 port map( A => mult_21_C243_n1391, Z => 
                           mult_21_C243_n1390);
   mult_21_C243_U1044 : INVD1 port map( A => mult_21_C243_n939, Z => 
                           mult_21_C243_n1420);
   mult_21_C243_U1043 : INVD1 port map( A => mult_21_C243_n940, Z => 
                           mult_21_C243_n1419);
   mult_21_C243_U1042 : INVD1 port map( A => mult_21_C243_n941, Z => 
                           mult_21_C243_n1416);
   mult_21_C243_U1041 : INVD1 port map( A => mult_21_C243_n942, Z => 
                           mult_21_C243_n1414);
   mult_21_C243_U1040 : INVD1 port map( A => mult_21_C243_n943, Z => 
                           mult_21_C243_n1412);
   mult_21_C243_U1039 : INVD1 port map( A => mult_21_C243_n944, Z => 
                           mult_21_C243_n1410);
   mult_21_C243_U1038 : INVD1 port map( A => mult_21_C243_n945, Z => 
                           mult_21_C243_n1408);
   mult_21_C243_U1037 : INVD1 port map( A => mult_21_C243_n946, Z => 
                           mult_21_C243_n1406);
   mult_21_C243_U1036 : INVD1 port map( A => mult_21_C243_n947, Z => 
                           mult_21_C243_n1404);
   mult_21_C243_U1035 : INVD1 port map( A => mult_21_C243_n948, Z => 
                           mult_21_C243_n1402);
   mult_21_C243_U1034 : INVD1 port map( A => mult_21_C243_n949, Z => 
                           mult_21_C243_n1400);
   mult_21_C243_U1033 : INVD1 port map( A => mult_21_C243_n950, Z => 
                           mult_21_C243_n1398);
   mult_21_C243_U1032 : INVD1 port map( A => mult_21_C243_n951, Z => 
                           mult_21_C243_n1396);
   mult_21_C243_U1031 : INVD1 port map( A => mult_21_C243_n952, Z => 
                           mult_21_C243_n1394);
   mult_21_C243_U1030 : INVD1 port map( A => mult_21_C243_n953, Z => 
                           mult_21_C243_n1393);
   mult_21_C243_U1029 : INVD1 port map( A => mult_21_C243_n1383, Z => 
                           mult_21_C243_n1385);
   mult_21_C243_U1028 : INVD1 port map( A => mult_21_C243_n1382, Z => 
                           mult_21_C243_n1384);
   mult_21_C243_U1027 : OAI21D1 port map( A1 => N2953, A2 => N2952, B => 
                           mult_21_C243_n1401, Z => mult_21_C243_n1381);
   mult_21_C243_U1026 : OAI21D1 port map( A1 => N2951, A2 => N2950, B => 
                           mult_21_C243_n1399, Z => mult_21_C243_n1380);
   mult_21_C243_U1025 : EXOR2D1 port map( A1 => N2953, A2 => N2952, Z => 
                           mult_21_C243_n1379);
   mult_21_C243_U1024 : EXOR2D1 port map( A1 => N2951, A2 => N2950, Z => 
                           mult_21_C243_n1378);
   mult_21_C243_U1023 : OAI21D1 port map( A1 => N2949, A2 => N2948, B => 
                           mult_21_C243_n1397, Z => mult_21_C243_n1377);
   mult_21_C243_U1022 : OAI21D1 port map( A1 => N2947, A2 => N2946, B => 
                           mult_21_C243_n1395, Z => mult_21_C243_n1376);
   mult_21_C243_U1021 : NAN2D1 port map( A1 => mult_21_C243_n1390, A2 => 
                           mult_21_C243_n1392, Z => mult_21_C243_n1375);
   mult_21_C243_U954 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n923, Z => 
                           mult_21_C243_n1226);
   mult_21_C243_U952 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n922, Z => 
                           mult_21_C243_n1225);
   mult_21_C243_U950 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n921, Z => 
                           mult_21_C243_n1224);
   mult_21_C243_U948 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n920, Z => 
                           mult_21_C243_n1223);
   mult_21_C243_U946 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n919, Z => 
                           mult_21_C243_n1222);
   mult_21_C243_U944 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n918, Z => 
                           mult_21_C243_n1221);
   mult_21_C243_U942 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n917, Z => 
                           mult_21_C243_n1220);
   mult_21_C243_U940 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n916, Z => 
                           mult_21_C243_n1219);
   mult_21_C243_U938 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n915, Z => 
                           mult_21_C243_n1218);
   mult_21_C243_U936 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n914, Z => 
                           mult_21_C243_n1217);
   mult_21_C243_U934 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n913, Z => 
                           mult_21_C243_n1216);
   mult_21_C243_U932 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n912, Z => 
                           mult_21_C243_n1215);
   mult_21_C243_U930 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n911, Z => 
                           mult_21_C243_n1214);
   mult_21_C243_U928 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n910, Z => 
                           mult_21_C243_n1213);
   mult_21_C243_U926 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n909, Z => 
                           mult_21_C243_n1212);
   mult_21_C243_U924 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n908, Z => 
                           mult_21_C243_n1211);
   mult_21_C243_U922 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n907, Z => 
                           mult_21_C243_n1210);
   mult_21_C243_U920 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n906, Z => 
                           mult_21_C243_n1209);
   mult_21_C243_U918 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n905, Z => 
                           mult_21_C243_n1208);
   mult_21_C243_U916 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n904, Z => 
                           mult_21_C243_n1207);
   mult_21_C243_U914 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n903, Z => 
                           mult_21_C243_n1206);
   mult_21_C243_U912 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n902, Z => 
                           mult_21_C243_n1205);
   mult_21_C243_U910 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n901, Z => 
                           mult_21_C243_n1204);
   mult_21_C243_U908 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n900, Z => 
                           mult_21_C243_n1203);
   mult_21_C243_U906 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n899, Z => 
                           mult_21_C243_n1202);
   mult_21_C243_U904 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n898, Z => 
                           mult_21_C243_n1201);
   mult_21_C243_U902 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n897, Z => 
                           mult_21_C243_n1200);
   mult_21_C243_U900 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n896, Z => 
                           mult_21_C243_n1199);
   mult_21_C243_U898 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n895, Z => 
                           mult_21_C243_n1198);
   mult_21_C243_U896 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n894, Z => 
                           mult_21_C243_n1197);
   mult_21_C243_U894 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n893, Z => 
                           mult_21_C243_n1196);
   mult_21_C243_U892 : MUXB2DL port map( A0 => mult_21_C243_n1375, A1 => 
                           mult_21_C243_n1392, SL => mult_21_C243_n892, Z => 
                           mult_21_C243_n1195);
   mult_21_C243_U889 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n891, Z => 
                           mult_21_C243_n1194);
   mult_21_C243_U887 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n890, Z => 
                           mult_21_C243_n1193);
   mult_21_C243_U885 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n889, Z => 
                           mult_21_C243_n1192);
   mult_21_C243_U883 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n888, Z => 
                           mult_21_C243_n1191);
   mult_21_C243_U881 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n887, Z => 
                           mult_21_C243_n1190);
   mult_21_C243_U879 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n886, Z => 
                           mult_21_C243_n1189);
   mult_21_C243_U877 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n885, Z => 
                           mult_21_C243_n1188);
   mult_21_C243_U875 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n884, Z => 
                           mult_21_C243_n1187);
   mult_21_C243_U873 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n883, Z => 
                           mult_21_C243_n1186);
   mult_21_C243_U871 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n882, Z => 
                           mult_21_C243_n1185);
   mult_21_C243_U869 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n881, Z => 
                           mult_21_C243_n1184);
   mult_21_C243_U867 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n880, Z => 
                           mult_21_C243_n1183);
   mult_21_C243_U865 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n879, Z => 
                           mult_21_C243_n1182);
   mult_21_C243_U863 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n878, Z => 
                           mult_21_C243_n1181);
   mult_21_C243_U861 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n877, Z => 
                           mult_21_C243_n1180);
   mult_21_C243_U859 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n876, Z => 
                           mult_21_C243_n1179);
   mult_21_C243_U857 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n875, Z => 
                           mult_21_C243_n1178);
   mult_21_C243_U855 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n874, Z => 
                           mult_21_C243_n1177);
   mult_21_C243_U853 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n873, Z => 
                           mult_21_C243_n1176);
   mult_21_C243_U851 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n872, Z => 
                           mult_21_C243_n1175);
   mult_21_C243_U849 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n871, Z => 
                           mult_21_C243_n1174);
   mult_21_C243_U847 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n870, Z => 
                           mult_21_C243_n1173);
   mult_21_C243_U845 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n869, Z => 
                           mult_21_C243_n1172);
   mult_21_C243_U843 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n868, Z => 
                           mult_21_C243_n1171);
   mult_21_C243_U841 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n867, Z => 
                           mult_21_C243_n1170);
   mult_21_C243_U839 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n866, Z => 
                           mult_21_C243_n1169);
   mult_21_C243_U837 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n865, Z => 
                           mult_21_C243_n1168);
   mult_21_C243_U835 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n864, Z => 
                           mult_21_C243_n1167);
   mult_21_C243_U833 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n863, Z => 
                           mult_21_C243_n1166);
   mult_21_C243_U831 : MUXB2DL port map( A0 => mult_21_C243_n1376, A1 => 
                           mult_21_C243_n1393, SL => mult_21_C243_n862, Z => 
                           mult_21_C243_n1165);
   mult_21_C243_U828 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n861, Z => 
                           mult_21_C243_n1164);
   mult_21_C243_U826 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n860, Z => 
                           mult_21_C243_n1163);
   mult_21_C243_U824 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n859, Z => 
                           mult_21_C243_n1162);
   mult_21_C243_U822 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n858, Z => 
                           mult_21_C243_n1161);
   mult_21_C243_U820 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n857, Z => 
                           mult_21_C243_n1160);
   mult_21_C243_U818 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n856, Z => 
                           mult_21_C243_n1159);
   mult_21_C243_U816 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n855, Z => 
                           mult_21_C243_n1158);
   mult_21_C243_U814 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n854, Z => 
                           mult_21_C243_n1157);
   mult_21_C243_U812 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n853, Z => 
                           mult_21_C243_n1156);
   mult_21_C243_U810 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n852, Z => 
                           mult_21_C243_n1155);
   mult_21_C243_U808 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n851, Z => 
                           mult_21_C243_n1154);
   mult_21_C243_U806 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n850, Z => 
                           mult_21_C243_n1153);
   mult_21_C243_U804 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n849, Z => 
                           mult_21_C243_n1152);
   mult_21_C243_U802 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n848, Z => 
                           mult_21_C243_n1151);
   mult_21_C243_U800 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n847, Z => 
                           mult_21_C243_n1150);
   mult_21_C243_U798 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n846, Z => 
                           mult_21_C243_n1149);
   mult_21_C243_U796 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n845, Z => 
                           mult_21_C243_n1148);
   mult_21_C243_U794 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n844, Z => 
                           mult_21_C243_n1147);
   mult_21_C243_U792 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n843, Z => 
                           mult_21_C243_n1146);
   mult_21_C243_U790 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n842, Z => 
                           mult_21_C243_n1145);
   mult_21_C243_U788 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n841, Z => 
                           mult_21_C243_n1144);
   mult_21_C243_U786 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n840, Z => 
                           mult_21_C243_n1143);
   mult_21_C243_U784 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n839, Z => 
                           mult_21_C243_n1142);
   mult_21_C243_U782 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n838, Z => 
                           mult_21_C243_n1141);
   mult_21_C243_U780 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n837, Z => 
                           mult_21_C243_n1140);
   mult_21_C243_U778 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n836, Z => 
                           mult_21_C243_n1139);
   mult_21_C243_U776 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n835, Z => 
                           mult_21_C243_n1138);
   mult_21_C243_U774 : MUXB2DL port map( A0 => mult_21_C243_n1377, A1 => 
                           mult_21_C243_n1394, SL => mult_21_C243_n834, Z => 
                           mult_21_C243_n1137);
   mult_21_C243_U771 : MUXB2DL port map( A0 => mult_21_C243_n1380, A1 => 
                           mult_21_C243_n1396, SL => mult_21_C243_n833, Z => 
                           mult_21_C243_n1136);
   mult_21_C243_U769 : MUXB2DL port map( A0 => mult_21_C243_n1380, A1 => 
                           mult_21_C243_n1396, SL => mult_21_C243_n832, Z => 
                           mult_21_C243_n1135);
   mult_21_C243_U767 : MUXB2DL port map( A0 => mult_21_C243_n1380, A1 => 
                           mult_21_C243_n1396, SL => mult_21_C243_n831, Z => 
                           mult_21_C243_n1134);
   mult_21_C243_U765 : MUXB2DL port map( A0 => mult_21_C243_n1380, A1 => 
                           mult_21_C243_n1396, SL => mult_21_C243_n830, Z => 
                           mult_21_C243_n1133);
   mult_21_C243_U763 : MUXB2DL port map( A0 => mult_21_C243_n1380, A1 => 
                           mult_21_C243_n1396, SL => mult_21_C243_n829, Z => 
                           mult_21_C243_n1132);
   mult_21_C243_U761 : MUXB2DL port map( A0 => mult_21_C243_n1380, A1 => 
                           mult_21_C243_n1396, SL => mult_21_C243_n828, Z => 
                           mult_21_C243_n1131);
   mult_21_C243_U759 : MUXB2DL port map( A0 => mult_21_C243_n1380, A1 => 
                           mult_21_C243_n1396, SL => mult_21_C243_n827, Z => 
                           mult_21_C243_n1130);
   mult_21_C243_U757 : MUXB2DL port map( A0 => mult_21_C243_n1380, A1 => 
                           mult_21_C243_n1396, SL => mult_21_C243_n826, Z => 
                           mult_21_C243_n1129);
   mult_21_C243_U755 : MUXB2DL port map( A0 => mult_21_C243_n1380, A1 => 
                           mult_21_C243_n1396, SL => mult_21_C243_n825, Z => 
                           mult_21_C243_n1128);
   mult_21_C243_U753 : MUXB2DL port map( A0 => mult_21_C243_n1380, A1 => 
                           mult_21_C243_n1396, SL => mult_21_C243_n824, Z => 
                           mult_21_C243_n1127);
   mult_21_C243_U751 : MUXB2DL port map( A0 => mult_21_C243_n1380, A1 => 
                           mult_21_C243_n1396, SL => mult_21_C243_n823, Z => 
                           mult_21_C243_n1126);
   mult_21_C243_U749 : MUXB2DL port map( A0 => mult_21_C243_n1380, A1 => 
                           mult_21_C243_n1396, SL => mult_21_C243_n822, Z => 
                           mult_21_C243_n1125);
   mult_21_C243_U747 : MUXB2DL port map( A0 => mult_21_C243_n1380, A1 => 
                           mult_21_C243_n1396, SL => mult_21_C243_n821, Z => 
                           mult_21_C243_n1124);
   mult_21_C243_U745 : MUXB2DL port map( A0 => mult_21_C243_n1380, A1 => 
                           mult_21_C243_n1396, SL => mult_21_C243_n820, Z => 
                           mult_21_C243_n1123);
   mult_21_C243_U743 : MUXB2DL port map( A0 => mult_21_C243_n1380, A1 => 
                           mult_21_C243_n1396, SL => mult_21_C243_n819, Z => 
                           mult_21_C243_n1122);
   mult_21_C243_U741 : MUXB2DL port map( A0 => mult_21_C243_n1380, A1 => 
                           mult_21_C243_n1396, SL => mult_21_C243_n818, Z => 
                           mult_21_C243_n1121);
   mult_21_C243_U739 : MUXB2DL port map( A0 => mult_21_C243_n1380, A1 => 
                           mult_21_C243_n1396, SL => mult_21_C243_n817, Z => 
                           mult_21_C243_n1120);
   mult_21_C243_U737 : MUXB2DL port map( A0 => mult_21_C243_n1380, A1 => 
                           mult_21_C243_n1396, SL => mult_21_C243_n816, Z => 
                           mult_21_C243_n1119);
   mult_21_C243_U735 : MUXB2DL port map( A0 => mult_21_C243_n1380, A1 => 
                           mult_21_C243_n1396, SL => mult_21_C243_n815, Z => 
                           mult_21_C243_n1118);
   mult_21_C243_U733 : MUXB2DL port map( A0 => mult_21_C243_n1380, A1 => 
                           mult_21_C243_n1396, SL => mult_21_C243_n814, Z => 
                           mult_21_C243_n1117);
   mult_21_C243_U731 : MUXB2DL port map( A0 => mult_21_C243_n1380, A1 => 
                           mult_21_C243_n1396, SL => mult_21_C243_n813, Z => 
                           mult_21_C243_n1116);
   mult_21_C243_U729 : MUXB2DL port map( A0 => mult_21_C243_n1380, A1 => 
                           mult_21_C243_n1396, SL => mult_21_C243_n812, Z => 
                           mult_21_C243_n1115);
   mult_21_C243_U727 : MUXB2DL port map( A0 => mult_21_C243_n1380, A1 => 
                           mult_21_C243_n1396, SL => mult_21_C243_n811, Z => 
                           mult_21_C243_n1114);
   mult_21_C243_U725 : MUXB2DL port map( A0 => mult_21_C243_n1380, A1 => 
                           mult_21_C243_n1396, SL => mult_21_C243_n810, Z => 
                           mult_21_C243_n1113);
   mult_21_C243_U723 : MUXB2DL port map( A0 => mult_21_C243_n1380, A1 => 
                           mult_21_C243_n1396, SL => mult_21_C243_n809, Z => 
                           mult_21_C243_n1112);
   mult_21_C243_U721 : MUXB2DL port map( A0 => mult_21_C243_n1380, A1 => 
                           mult_21_C243_n1396, SL => mult_21_C243_n808, Z => 
                           mult_21_C243_n1111);
   mult_21_C243_U718 : MUXB2DL port map( A0 => mult_21_C243_n1381, A1 => 
                           mult_21_C243_n1398, SL => mult_21_C243_n807, Z => 
                           mult_21_C243_n1110);
   mult_21_C243_U716 : MUXB2DL port map( A0 => mult_21_C243_n1381, A1 => 
                           mult_21_C243_n1398, SL => mult_21_C243_n806, Z => 
                           mult_21_C243_n1109);
   mult_21_C243_U714 : MUXB2DL port map( A0 => mult_21_C243_n1381, A1 => 
                           mult_21_C243_n1398, SL => mult_21_C243_n805, Z => 
                           mult_21_C243_n1108);
   mult_21_C243_U712 : MUXB2DL port map( A0 => mult_21_C243_n1381, A1 => 
                           mult_21_C243_n1398, SL => mult_21_C243_n804, Z => 
                           mult_21_C243_n1107);
   mult_21_C243_U710 : MUXB2DL port map( A0 => mult_21_C243_n1381, A1 => 
                           mult_21_C243_n1398, SL => mult_21_C243_n803, Z => 
                           mult_21_C243_n1106);
   mult_21_C243_U708 : MUXB2DL port map( A0 => mult_21_C243_n1381, A1 => 
                           mult_21_C243_n1398, SL => mult_21_C243_n802, Z => 
                           mult_21_C243_n1105);
   mult_21_C243_U706 : MUXB2DL port map( A0 => mult_21_C243_n1381, A1 => 
                           mult_21_C243_n1398, SL => mult_21_C243_n801, Z => 
                           mult_21_C243_n1104);
   mult_21_C243_U704 : MUXB2DL port map( A0 => mult_21_C243_n1381, A1 => 
                           mult_21_C243_n1398, SL => mult_21_C243_n800, Z => 
                           mult_21_C243_n1103);
   mult_21_C243_U702 : MUXB2DL port map( A0 => mult_21_C243_n1381, A1 => 
                           mult_21_C243_n1398, SL => mult_21_C243_n799, Z => 
                           mult_21_C243_n1102);
   mult_21_C243_U700 : MUXB2DL port map( A0 => mult_21_C243_n1381, A1 => 
                           mult_21_C243_n1398, SL => mult_21_C243_n798, Z => 
                           mult_21_C243_n1101);
   mult_21_C243_U698 : MUXB2DL port map( A0 => mult_21_C243_n1381, A1 => 
                           mult_21_C243_n1398, SL => mult_21_C243_n797, Z => 
                           mult_21_C243_n1100);
   mult_21_C243_U696 : MUXB2DL port map( A0 => mult_21_C243_n1381, A1 => 
                           mult_21_C243_n1398, SL => mult_21_C243_n796, Z => 
                           mult_21_C243_n1099);
   mult_21_C243_U694 : MUXB2DL port map( A0 => mult_21_C243_n1381, A1 => 
                           mult_21_C243_n1398, SL => mult_21_C243_n795, Z => 
                           mult_21_C243_n1098);
   mult_21_C243_U692 : MUXB2DL port map( A0 => mult_21_C243_n1381, A1 => 
                           mult_21_C243_n1398, SL => mult_21_C243_n794, Z => 
                           mult_21_C243_n1097);
   mult_21_C243_U690 : MUXB2DL port map( A0 => mult_21_C243_n1381, A1 => 
                           mult_21_C243_n1398, SL => mult_21_C243_n793, Z => 
                           mult_21_C243_n1096);
   mult_21_C243_U688 : MUXB2DL port map( A0 => mult_21_C243_n1381, A1 => 
                           mult_21_C243_n1398, SL => mult_21_C243_n792, Z => 
                           mult_21_C243_n1095);
   mult_21_C243_U686 : MUXB2DL port map( A0 => mult_21_C243_n1381, A1 => 
                           mult_21_C243_n1398, SL => mult_21_C243_n791, Z => 
                           mult_21_C243_n1094);
   mult_21_C243_U684 : MUXB2DL port map( A0 => mult_21_C243_n1381, A1 => 
                           mult_21_C243_n1398, SL => mult_21_C243_n790, Z => 
                           mult_21_C243_n1093);
   mult_21_C243_U682 : MUXB2DL port map( A0 => mult_21_C243_n1381, A1 => 
                           mult_21_C243_n1398, SL => mult_21_C243_n789, Z => 
                           mult_21_C243_n1092);
   mult_21_C243_U680 : MUXB2DL port map( A0 => mult_21_C243_n1381, A1 => 
                           mult_21_C243_n1398, SL => mult_21_C243_n788, Z => 
                           mult_21_C243_n1091);
   mult_21_C243_U678 : MUXB2DL port map( A0 => mult_21_C243_n1381, A1 => 
                           mult_21_C243_n1398, SL => mult_21_C243_n787, Z => 
                           mult_21_C243_n1090);
   mult_21_C243_U676 : MUXB2DL port map( A0 => mult_21_C243_n1381, A1 => 
                           mult_21_C243_n1398, SL => mult_21_C243_n786, Z => 
                           mult_21_C243_n1089);
   mult_21_C243_U674 : MUXB2DL port map( A0 => mult_21_C243_n1381, A1 => 
                           mult_21_C243_n1398, SL => mult_21_C243_n785, Z => 
                           mult_21_C243_n1088);
   mult_21_C243_U672 : MUXB2DL port map( A0 => mult_21_C243_n1381, A1 => 
                           mult_21_C243_n1398, SL => mult_21_C243_n784, Z => 
                           mult_21_C243_n1087);
   mult_21_C243_U669 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n1400, SL => mult_21_C243_n783, Z => 
                           mult_21_C243_n1086);
   mult_21_C243_U667 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n1400, SL => mult_21_C243_n782, Z => 
                           mult_21_C243_n1085);
   mult_21_C243_U665 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n1400, SL => mult_21_C243_n781, Z => 
                           mult_21_C243_n1084);
   mult_21_C243_U663 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n1400, SL => mult_21_C243_n780, Z => 
                           mult_21_C243_n1083);
   mult_21_C243_U661 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n1400, SL => mult_21_C243_n779, Z => 
                           mult_21_C243_n1082);
   mult_21_C243_U659 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n1400, SL => mult_21_C243_n778, Z => 
                           mult_21_C243_n1081);
   mult_21_C243_U657 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n1400, SL => mult_21_C243_n777, Z => 
                           mult_21_C243_n1080);
   mult_21_C243_U655 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n1400, SL => mult_21_C243_n776, Z => 
                           mult_21_C243_n1079);
   mult_21_C243_U653 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n1400, SL => mult_21_C243_n775, Z => 
                           mult_21_C243_n1078);
   mult_21_C243_U651 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n1400, SL => mult_21_C243_n774, Z => 
                           mult_21_C243_n1077);
   mult_21_C243_U649 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n1400, SL => mult_21_C243_n773, Z => 
                           mult_21_C243_n1076);
   mult_21_C243_U647 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n1400, SL => mult_21_C243_n772, Z => 
                           mult_21_C243_n1075);
   mult_21_C243_U645 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n1400, SL => mult_21_C243_n771, Z => 
                           mult_21_C243_n1074);
   mult_21_C243_U643 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n1400, SL => mult_21_C243_n770, Z => 
                           mult_21_C243_n1073);
   mult_21_C243_U641 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n1400, SL => mult_21_C243_n769, Z => 
                           mult_21_C243_n1072);
   mult_21_C243_U639 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n1400, SL => mult_21_C243_n768, Z => 
                           mult_21_C243_n1071);
   mult_21_C243_U637 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n1400, SL => mult_21_C243_n767, Z => 
                           mult_21_C243_n1070);
   mult_21_C243_U635 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n1400, SL => mult_21_C243_n766, Z => 
                           mult_21_C243_n1069);
   mult_21_C243_U633 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n1400, SL => mult_21_C243_n765, Z => 
                           mult_21_C243_n1068);
   mult_21_C243_U631 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n1400, SL => mult_21_C243_n764, Z => 
                           mult_21_C243_n1067);
   mult_21_C243_U629 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n1400, SL => mult_21_C243_n763, Z => 
                           mult_21_C243_n1066);
   mult_21_C243_U627 : MUXB2DL port map( A0 => mult_21_C243_n42, A1 => 
                           mult_21_C243_n1400, SL => mult_21_C243_n762, Z => 
                           mult_21_C243_n1065);
   mult_21_C243_U624 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n1402, SL => mult_21_C243_n761, Z => 
                           mult_21_C243_n1064);
   mult_21_C243_U622 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n1402, SL => mult_21_C243_n760, Z => 
                           mult_21_C243_n1063);
   mult_21_C243_U620 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n1402, SL => mult_21_C243_n759, Z => 
                           mult_21_C243_n1062);
   mult_21_C243_U618 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n1402, SL => mult_21_C243_n758, Z => 
                           mult_21_C243_n1061);
   mult_21_C243_U616 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n1402, SL => mult_21_C243_n757, Z => 
                           mult_21_C243_n1060);
   mult_21_C243_U614 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n1402, SL => mult_21_C243_n756, Z => 
                           mult_21_C243_n1059);
   mult_21_C243_U612 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n1402, SL => mult_21_C243_n755, Z => 
                           mult_21_C243_n1058);
   mult_21_C243_U610 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n1402, SL => mult_21_C243_n754, Z => 
                           mult_21_C243_n1057);
   mult_21_C243_U608 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n1402, SL => mult_21_C243_n753, Z => 
                           mult_21_C243_n1056);
   mult_21_C243_U606 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n1402, SL => mult_21_C243_n752, Z => 
                           mult_21_C243_n1055);
   mult_21_C243_U604 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n1402, SL => mult_21_C243_n751, Z => 
                           mult_21_C243_n1054);
   mult_21_C243_U602 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n1402, SL => mult_21_C243_n750, Z => 
                           mult_21_C243_n1053);
   mult_21_C243_U600 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n1402, SL => mult_21_C243_n749, Z => 
                           mult_21_C243_n1052);
   mult_21_C243_U598 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n1402, SL => mult_21_C243_n748, Z => 
                           mult_21_C243_n1051);
   mult_21_C243_U596 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n1402, SL => mult_21_C243_n747, Z => 
                           mult_21_C243_n1050);
   mult_21_C243_U594 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n1402, SL => mult_21_C243_n746, Z => 
                           mult_21_C243_n1049);
   mult_21_C243_U592 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n1402, SL => mult_21_C243_n745, Z => 
                           mult_21_C243_n1048);
   mult_21_C243_U590 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n1402, SL => mult_21_C243_n744, Z => 
                           mult_21_C243_n1047);
   mult_21_C243_U588 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n1402, SL => mult_21_C243_n743, Z => 
                           mult_21_C243_n1046);
   mult_21_C243_U586 : MUXB2DL port map( A0 => mult_21_C243_n50, A1 => 
                           mult_21_C243_n1402, SL => mult_21_C243_n742, Z => 
                           mult_21_C243_n1045);
   mult_21_C243_U583 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n1404, SL => mult_21_C243_n741, Z => 
                           mult_21_C243_n1044);
   mult_21_C243_U581 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n1404, SL => mult_21_C243_n740, Z => 
                           mult_21_C243_n1043);
   mult_21_C243_U579 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n1404, SL => mult_21_C243_n739, Z => 
                           mult_21_C243_n1042);
   mult_21_C243_U577 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n1404, SL => mult_21_C243_n738, Z => 
                           mult_21_C243_n1041);
   mult_21_C243_U575 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n1404, SL => mult_21_C243_n737, Z => 
                           mult_21_C243_n1040);
   mult_21_C243_U573 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n1404, SL => mult_21_C243_n736, Z => 
                           mult_21_C243_n1039);
   mult_21_C243_U571 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n1404, SL => mult_21_C243_n735, Z => 
                           mult_21_C243_n1038);
   mult_21_C243_U569 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n1404, SL => mult_21_C243_n734, Z => 
                           mult_21_C243_n1037);
   mult_21_C243_U567 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n1404, SL => mult_21_C243_n733, Z => 
                           mult_21_C243_n1036);
   mult_21_C243_U565 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n1404, SL => mult_21_C243_n732, Z => 
                           mult_21_C243_n1035);
   mult_21_C243_U563 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n1404, SL => mult_21_C243_n731, Z => 
                           mult_21_C243_n1034);
   mult_21_C243_U561 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n1404, SL => mult_21_C243_n730, Z => 
                           mult_21_C243_n1033);
   mult_21_C243_U559 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n1404, SL => mult_21_C243_n729, Z => 
                           mult_21_C243_n1032);
   mult_21_C243_U557 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n1404, SL => mult_21_C243_n728, Z => 
                           mult_21_C243_n1031);
   mult_21_C243_U555 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n1404, SL => mult_21_C243_n727, Z => 
                           mult_21_C243_n1030);
   mult_21_C243_U553 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n1404, SL => mult_21_C243_n726, Z => 
                           mult_21_C243_n1029);
   mult_21_C243_U551 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n1404, SL => mult_21_C243_n725, Z => 
                           mult_21_C243_n1028);
   mult_21_C243_U549 : MUXB2DL port map( A0 => mult_21_C243_n58, A1 => 
                           mult_21_C243_n1404, SL => mult_21_C243_n724, Z => 
                           mult_21_C243_n1027);
   mult_21_C243_U546 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n1406, SL => mult_21_C243_n723, Z => 
                           mult_21_C243_n1026);
   mult_21_C243_U544 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n1406, SL => mult_21_C243_n722, Z => 
                           mult_21_C243_n1025);
   mult_21_C243_U542 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n1406, SL => mult_21_C243_n721, Z => 
                           mult_21_C243_n1024);
   mult_21_C243_U540 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n1406, SL => mult_21_C243_n720, Z => 
                           mult_21_C243_n1023);
   mult_21_C243_U538 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n1406, SL => mult_21_C243_n719, Z => 
                           mult_21_C243_n1022);
   mult_21_C243_U536 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n1406, SL => mult_21_C243_n718, Z => 
                           mult_21_C243_n1021);
   mult_21_C243_U534 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n1406, SL => mult_21_C243_n717, Z => 
                           mult_21_C243_n1020);
   mult_21_C243_U532 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n1406, SL => mult_21_C243_n716, Z => 
                           mult_21_C243_n1019);
   mult_21_C243_U530 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n1406, SL => mult_21_C243_n715, Z => 
                           mult_21_C243_n1018);
   mult_21_C243_U528 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n1406, SL => mult_21_C243_n714, Z => 
                           mult_21_C243_n1017);
   mult_21_C243_U526 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n1406, SL => mult_21_C243_n713, Z => 
                           mult_21_C243_n1016);
   mult_21_C243_U524 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n1406, SL => mult_21_C243_n712, Z => 
                           mult_21_C243_n1015);
   mult_21_C243_U522 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n1406, SL => mult_21_C243_n711, Z => 
                           mult_21_C243_n1014);
   mult_21_C243_U520 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n1406, SL => mult_21_C243_n710, Z => 
                           mult_21_C243_n1013);
   mult_21_C243_U518 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n1406, SL => mult_21_C243_n709, Z => 
                           mult_21_C243_n1012);
   mult_21_C243_U516 : MUXB2DL port map( A0 => mult_21_C243_n66, A1 => 
                           mult_21_C243_n1406, SL => mult_21_C243_n708, Z => 
                           mult_21_C243_n1011);
   mult_21_C243_U513 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n1408, SL => mult_21_C243_n707, Z => 
                           mult_21_C243_n1010);
   mult_21_C243_U511 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n1408, SL => mult_21_C243_n706, Z => 
                           mult_21_C243_n1009);
   mult_21_C243_U509 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n1408, SL => mult_21_C243_n705, Z => 
                           mult_21_C243_n1008);
   mult_21_C243_U507 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n1408, SL => mult_21_C243_n704, Z => 
                           mult_21_C243_n1007);
   mult_21_C243_U505 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n1408, SL => mult_21_C243_n703, Z => 
                           mult_21_C243_n1006);
   mult_21_C243_U503 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n1408, SL => mult_21_C243_n702, Z => 
                           mult_21_C243_n1005);
   mult_21_C243_U501 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n1408, SL => mult_21_C243_n701, Z => 
                           mult_21_C243_n1004);
   mult_21_C243_U499 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n1408, SL => mult_21_C243_n700, Z => 
                           mult_21_C243_n1003);
   mult_21_C243_U497 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n1408, SL => mult_21_C243_n699, Z => 
                           mult_21_C243_n1002);
   mult_21_C243_U495 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n1408, SL => mult_21_C243_n698, Z => 
                           mult_21_C243_n1001);
   mult_21_C243_U493 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n1408, SL => mult_21_C243_n697, Z => 
                           mult_21_C243_n1000);
   mult_21_C243_U491 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n1408, SL => mult_21_C243_n696, Z => 
                           mult_21_C243_n999);
   mult_21_C243_U489 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n1408, SL => mult_21_C243_n695, Z => 
                           mult_21_C243_n998);
   mult_21_C243_U487 : MUXB2DL port map( A0 => mult_21_C243_n73, A1 => 
                           mult_21_C243_n1408, SL => mult_21_C243_n694, Z => 
                           mult_21_C243_n997);
   mult_21_C243_U484 : MUXB2DL port map( A0 => mult_21_C243_n80, A1 => 
                           mult_21_C243_n1410, SL => mult_21_C243_n693, Z => 
                           mult_21_C243_n996);
   mult_21_C243_U482 : MUXB2DL port map( A0 => mult_21_C243_n80, A1 => 
                           mult_21_C243_n1410, SL => mult_21_C243_n692, Z => 
                           mult_21_C243_n995);
   mult_21_C243_U480 : MUXB2DL port map( A0 => mult_21_C243_n80, A1 => 
                           mult_21_C243_n1410, SL => mult_21_C243_n691, Z => 
                           mult_21_C243_n994);
   mult_21_C243_U478 : MUXB2DL port map( A0 => mult_21_C243_n80, A1 => 
                           mult_21_C243_n1410, SL => mult_21_C243_n690, Z => 
                           mult_21_C243_n993);
   mult_21_C243_U476 : MUXB2DL port map( A0 => mult_21_C243_n80, A1 => 
                           mult_21_C243_n1410, SL => mult_21_C243_n689, Z => 
                           mult_21_C243_n992);
   mult_21_C243_U474 : MUXB2DL port map( A0 => mult_21_C243_n80, A1 => 
                           mult_21_C243_n1410, SL => mult_21_C243_n688, Z => 
                           mult_21_C243_n991);
   mult_21_C243_U472 : MUXB2DL port map( A0 => mult_21_C243_n80, A1 => 
                           mult_21_C243_n1410, SL => mult_21_C243_n687, Z => 
                           mult_21_C243_n990);
   mult_21_C243_U470 : MUXB2DL port map( A0 => mult_21_C243_n80, A1 => 
                           mult_21_C243_n1410, SL => mult_21_C243_n686, Z => 
                           mult_21_C243_n989);
   mult_21_C243_U468 : MUXB2DL port map( A0 => mult_21_C243_n80, A1 => 
                           mult_21_C243_n1410, SL => mult_21_C243_n685, Z => 
                           mult_21_C243_n988);
   mult_21_C243_U466 : MUXB2DL port map( A0 => mult_21_C243_n80, A1 => 
                           mult_21_C243_n1410, SL => mult_21_C243_n684, Z => 
                           mult_21_C243_n987);
   mult_21_C243_U464 : MUXB2DL port map( A0 => mult_21_C243_n80, A1 => 
                           mult_21_C243_n1410, SL => mult_21_C243_n683, Z => 
                           mult_21_C243_n986);
   mult_21_C243_U462 : MUXB2DL port map( A0 => mult_21_C243_n80, A1 => 
                           mult_21_C243_n1410, SL => mult_21_C243_n682, Z => 
                           mult_21_C243_n985);
   mult_21_C243_U459 : MUXB2DL port map( A0 => mult_21_C243_n84, A1 => 
                           mult_21_C243_n1412, SL => mult_21_C243_n681, Z => 
                           mult_21_C243_n984);
   mult_21_C243_U457 : MUXB2DL port map( A0 => mult_21_C243_n84, A1 => 
                           mult_21_C243_n1412, SL => mult_21_C243_n680, Z => 
                           mult_21_C243_n983);
   mult_21_C243_U455 : MUXB2DL port map( A0 => mult_21_C243_n84, A1 => 
                           mult_21_C243_n1412, SL => mult_21_C243_n679, Z => 
                           mult_21_C243_n982);
   mult_21_C243_U453 : MUXB2DL port map( A0 => mult_21_C243_n84, A1 => 
                           mult_21_C243_n1412, SL => mult_21_C243_n678, Z => 
                           mult_21_C243_n981);
   mult_21_C243_U451 : MUXB2DL port map( A0 => mult_21_C243_n84, A1 => 
                           mult_21_C243_n1412, SL => mult_21_C243_n677, Z => 
                           mult_21_C243_n980);
   mult_21_C243_U449 : MUXB2DL port map( A0 => mult_21_C243_n84, A1 => 
                           mult_21_C243_n1412, SL => mult_21_C243_n676, Z => 
                           mult_21_C243_n979);
   mult_21_C243_U447 : MUXB2DL port map( A0 => mult_21_C243_n84, A1 => 
                           mult_21_C243_n1412, SL => mult_21_C243_n675, Z => 
                           mult_21_C243_n978);
   mult_21_C243_U445 : MUXB2DL port map( A0 => mult_21_C243_n84, A1 => 
                           mult_21_C243_n1412, SL => mult_21_C243_n674, Z => 
                           mult_21_C243_n977);
   mult_21_C243_U443 : MUXB2DL port map( A0 => mult_21_C243_n84, A1 => 
                           mult_21_C243_n1412, SL => mult_21_C243_n673, Z => 
                           mult_21_C243_n976);
   mult_21_C243_U441 : MUXB2DL port map( A0 => mult_21_C243_n84, A1 => 
                           mult_21_C243_n1412, SL => mult_21_C243_n672, Z => 
                           mult_21_C243_n975);
   mult_21_C243_U438 : MUXB2DL port map( A0 => mult_21_C243_n89, A1 => 
                           mult_21_C243_n1414, SL => mult_21_C243_n671, Z => 
                           mult_21_C243_n974);
   mult_21_C243_U436 : MUXB2DL port map( A0 => mult_21_C243_n89, A1 => 
                           mult_21_C243_n1414, SL => mult_21_C243_n670, Z => 
                           mult_21_C243_n973);
   mult_21_C243_U434 : MUXB2DL port map( A0 => mult_21_C243_n89, A1 => 
                           mult_21_C243_n1414, SL => mult_21_C243_n669, Z => 
                           mult_21_C243_n972);
   mult_21_C243_U432 : MUXB2DL port map( A0 => mult_21_C243_n89, A1 => 
                           mult_21_C243_n1414, SL => mult_21_C243_n668, Z => 
                           mult_21_C243_n971);
   mult_21_C243_U430 : MUXB2DL port map( A0 => mult_21_C243_n89, A1 => 
                           mult_21_C243_n1414, SL => mult_21_C243_n667, Z => 
                           mult_21_C243_n970);
   mult_21_C243_U428 : MUXB2DL port map( A0 => mult_21_C243_n89, A1 => 
                           mult_21_C243_n1414, SL => mult_21_C243_n666, Z => 
                           mult_21_C243_n969);
   mult_21_C243_U426 : MUXB2DL port map( A0 => mult_21_C243_n89, A1 => 
                           mult_21_C243_n1414, SL => mult_21_C243_n665, Z => 
                           mult_21_C243_n968);
   mult_21_C243_U424 : MUXB2DL port map( A0 => mult_21_C243_n89, A1 => 
                           mult_21_C243_n1414, SL => mult_21_C243_n664, Z => 
                           mult_21_C243_n967);
   mult_21_C243_U421 : MUXB2DL port map( A0 => mult_21_C243_n94, A1 => 
                           mult_21_C243_n1416, SL => mult_21_C243_n663, Z => 
                           mult_21_C243_n966);
   mult_21_C243_U419 : MUXB2DL port map( A0 => mult_21_C243_n94, A1 => 
                           mult_21_C243_n1416, SL => mult_21_C243_n662, Z => 
                           mult_21_C243_n965);
   mult_21_C243_U417 : MUXB2DL port map( A0 => mult_21_C243_n94, A1 => 
                           mult_21_C243_n1416, SL => mult_21_C243_n661, Z => 
                           mult_21_C243_n964);
   mult_21_C243_U415 : MUXB2DL port map( A0 => mult_21_C243_n94, A1 => 
                           mult_21_C243_n1416, SL => mult_21_C243_n660, Z => 
                           mult_21_C243_n963);
   mult_21_C243_U413 : MUXB2DL port map( A0 => mult_21_C243_n94, A1 => 
                           mult_21_C243_n1416, SL => mult_21_C243_n659, Z => 
                           mult_21_C243_n962);
   mult_21_C243_U411 : MUXB2DL port map( A0 => mult_21_C243_n94, A1 => 
                           mult_21_C243_n1416, SL => mult_21_C243_n658, Z => 
                           mult_21_C243_n961);
   mult_21_C243_U408 : MUXB2DL port map( A0 => mult_21_C243_n99, A1 => 
                           mult_21_C243_n1419, SL => mult_21_C243_n657, Z => 
                           mult_21_C243_n960);
   mult_21_C243_U406 : MUXB2DL port map( A0 => mult_21_C243_n99, A1 => 
                           mult_21_C243_n1419, SL => mult_21_C243_n656, Z => 
                           mult_21_C243_n959);
   mult_21_C243_U404 : MUXB2DL port map( A0 => mult_21_C243_n99, A1 => 
                           mult_21_C243_n1419, SL => mult_21_C243_n655, Z => 
                           mult_21_C243_n958);
   mult_21_C243_U402 : MUXB2DL port map( A0 => mult_21_C243_n99, A1 => 
                           mult_21_C243_n1419, SL => mult_21_C243_n654, Z => 
                           mult_21_C243_n957);
   mult_21_C243_U399 : MUXB2DL port map( A0 => mult_21_C243_n104, A1 => 
                           mult_21_C243_n1420, SL => mult_21_C243_n653, Z => 
                           mult_21_C243_n956);
   mult_21_C243_U397 : MUXB2DL port map( A0 => mult_21_C243_n104, A1 => 
                           mult_21_C243_n1420, SL => mult_21_C243_n652, Z => 
                           mult_21_C243_n955);
   mult_21_C243_U395 : ADHALFDL port map( A => mult_21_C243_n1224, B => 
                           mult_21_C243_n953, CO => mult_21_C243_n650, S => 
                           mult_21_C243_n651);
   mult_21_C243_U394 : ADHALFDL port map( A => mult_21_C243_n650, B => 
                           mult_21_C243_n1223, CO => mult_21_C243_n648, S => 
                           mult_21_C243_n649);
   mult_21_C243_U393 : ADHALFDL port map( A => mult_21_C243_n1222, B => 
                           mult_21_C243_n952, CO => mult_21_C243_n646, S => 
                           mult_21_C243_n647);
   mult_21_C243_U392 : ADFULD1 port map( A => mult_21_C243_n1192, B => 
                           mult_21_C243_n1164, CI => mult_21_C243_n647, CO => 
                           mult_21_C243_n644, S => mult_21_C243_n645);
   mult_21_C243_U391 : ADHALFDL port map( A => mult_21_C243_n646, B => 
                           mult_21_C243_n1221, CO => mult_21_C243_n642, S => 
                           mult_21_C243_n643);
   mult_21_C243_U390 : ADFULD1 port map( A => mult_21_C243_n1163, B => 
                           mult_21_C243_n1191, CI => mult_21_C243_n643, CO => 
                           mult_21_C243_n640, S => mult_21_C243_n641);
   mult_21_C243_U389 : ADHALFDL port map( A => mult_21_C243_n1220, B => 
                           mult_21_C243_n951, CO => mult_21_C243_n638, S => 
                           mult_21_C243_n639);
   mult_21_C243_U388 : ADFULD1 port map( A => mult_21_C243_n1190, B => 
                           mult_21_C243_n1136, CI => mult_21_C243_n1162, CO => 
                           mult_21_C243_n636, S => mult_21_C243_n637);
   mult_21_C243_U387 : ADFULD1 port map( A => mult_21_C243_n642, B => 
                           mult_21_C243_n639, CI => mult_21_C243_n637, CO => 
                           mult_21_C243_n634, S => mult_21_C243_n635);
   mult_21_C243_U386 : ADHALFDL port map( A => mult_21_C243_n638, B => 
                           mult_21_C243_n1219, CO => mult_21_C243_n632, S => 
                           mult_21_C243_n633);
   mult_21_C243_U385 : ADFULD1 port map( A => mult_21_C243_n1135, B => 
                           mult_21_C243_n1189, CI => mult_21_C243_n1161, CO => 
                           mult_21_C243_n630, S => mult_21_C243_n631);
   mult_21_C243_U384 : ADFULD1 port map( A => mult_21_C243_n636, B => 
                           mult_21_C243_n633, CI => mult_21_C243_n631, CO => 
                           mult_21_C243_n628, S => mult_21_C243_n629);
   mult_21_C243_U383 : ADHALFDL port map( A => mult_21_C243_n1218, B => 
                           mult_21_C243_n950, CO => mult_21_C243_n626, S => 
                           mult_21_C243_n627);
   mult_21_C243_U382 : ADFULD1 port map( A => mult_21_C243_n1188, B => 
                           mult_21_C243_n1110, CI => mult_21_C243_n1134, CO => 
                           mult_21_C243_n624, S => mult_21_C243_n625);
   mult_21_C243_U381 : ADFULD1 port map( A => mult_21_C243_n627, B => 
                           mult_21_C243_n1160, CI => mult_21_C243_n632, CO => 
                           mult_21_C243_n622, S => mult_21_C243_n623);
   mult_21_C243_U380 : ADFULD1 port map( A => mult_21_C243_n625, B => 
                           mult_21_C243_n630, CI => mult_21_C243_n623, CO => 
                           mult_21_C243_n620, S => mult_21_C243_n621);
   mult_21_C243_U379 : ADHALFDL port map( A => mult_21_C243_n626, B => 
                           mult_21_C243_n1217, CO => mult_21_C243_n618, S => 
                           mult_21_C243_n619);
   mult_21_C243_U378 : ADFULD1 port map( A => mult_21_C243_n1109, B => 
                           mult_21_C243_n1133, CI => mult_21_C243_n1159, CO => 
                           mult_21_C243_n616, S => mult_21_C243_n617);
   mult_21_C243_U377 : ADFULD1 port map( A => mult_21_C243_n619, B => 
                           mult_21_C243_n1187, CI => mult_21_C243_n624, CO => 
                           mult_21_C243_n614, S => mult_21_C243_n615);
   mult_21_C243_U376 : ADFULD1 port map( A => mult_21_C243_n617, B => 
                           mult_21_C243_n622, CI => mult_21_C243_n615, CO => 
                           mult_21_C243_n612, S => mult_21_C243_n613);
   mult_21_C243_U375 : ADHALFDL port map( A => mult_21_C243_n1216, B => 
                           mult_21_C243_n949, CO => mult_21_C243_n610, S => 
                           mult_21_C243_n611);
   mult_21_C243_U374 : ADFULD1 port map( A => mult_21_C243_n1132, B => 
                           mult_21_C243_n1086, CI => mult_21_C243_n1186, CO => 
                           mult_21_C243_n608, S => mult_21_C243_n609);
   mult_21_C243_U373 : ADFULD1 port map( A => mult_21_C243_n1108, B => 
                           mult_21_C243_n1158, CI => mult_21_C243_n611, CO => 
                           mult_21_C243_n606, S => mult_21_C243_n607);
   mult_21_C243_U372 : ADFULD1 port map( A => mult_21_C243_n616, B => 
                           mult_21_C243_n618, CI => mult_21_C243_n609, CO => 
                           mult_21_C243_n604, S => mult_21_C243_n605);
   mult_21_C243_U371 : ADFULD1 port map( A => mult_21_C243_n614, B => 
                           mult_21_C243_n607, CI => mult_21_C243_n605, CO => 
                           mult_21_C243_n602, S => mult_21_C243_n603);
   mult_21_C243_U370 : ADHALFDL port map( A => mult_21_C243_n610, B => 
                           mult_21_C243_n1215, CO => mult_21_C243_n600, S => 
                           mult_21_C243_n601);
   mult_21_C243_U369 : ADFULD1 port map( A => mult_21_C243_n1085, B => 
                           mult_21_C243_n1131, CI => mult_21_C243_n1185, CO => 
                           mult_21_C243_n598, S => mult_21_C243_n599);
   mult_21_C243_U368 : ADFULD1 port map( A => mult_21_C243_n1107, B => 
                           mult_21_C243_n1157, CI => mult_21_C243_n601, CO => 
                           mult_21_C243_n596, S => mult_21_C243_n597);
   mult_21_C243_U367 : ADFULD1 port map( A => mult_21_C243_n606, B => 
                           mult_21_C243_n608, CI => mult_21_C243_n599, CO => 
                           mult_21_C243_n594, S => mult_21_C243_n595);
   mult_21_C243_U366 : ADFULD1 port map( A => mult_21_C243_n604, B => 
                           mult_21_C243_n597, CI => mult_21_C243_n595, CO => 
                           mult_21_C243_n592, S => mult_21_C243_n593);
   mult_21_C243_U365 : ADHALFDL port map( A => mult_21_C243_n1214, B => 
                           mult_21_C243_n948, CO => mult_21_C243_n590, S => 
                           mult_21_C243_n591);
   mult_21_C243_U364 : ADFULD1 port map( A => mult_21_C243_n1130, B => 
                           mult_21_C243_n1064, CI => mult_21_C243_n1184, CO => 
                           mult_21_C243_n588, S => mult_21_C243_n589);
   mult_21_C243_U363 : ADFULD1 port map( A => mult_21_C243_n1084, B => 
                           mult_21_C243_n1156, CI => mult_21_C243_n591, CO => 
                           mult_21_C243_n586, S => mult_21_C243_n587);
   mult_21_C243_U362 : ADFULD1 port map( A => mult_21_C243_n600, B => 
                           mult_21_C243_n1106, CI => mult_21_C243_n598, CO => 
                           mult_21_C243_n584, S => mult_21_C243_n585);
   mult_21_C243_U361 : ADFULD1 port map( A => mult_21_C243_n587, B => 
                           mult_21_C243_n589, CI => mult_21_C243_n596, CO => 
                           mult_21_C243_n582, S => mult_21_C243_n583);
   mult_21_C243_U360 : ADFULD1 port map( A => mult_21_C243_n585, B => 
                           mult_21_C243_n594, CI => mult_21_C243_n583, CO => 
                           mult_21_C243_n580, S => mult_21_C243_n581);
   mult_21_C243_U359 : ADHALFDL port map( A => mult_21_C243_n590, B => 
                           mult_21_C243_n1213, CO => mult_21_C243_n578, S => 
                           mult_21_C243_n579);
   mult_21_C243_U358 : ADFULD1 port map( A => mult_21_C243_n1183, B => 
                           mult_21_C243_n1105, CI => mult_21_C243_n1155, CO => 
                           mult_21_C243_n576, S => mult_21_C243_n577);
   mult_21_C243_U357 : ADFULD1 port map( A => mult_21_C243_n1063, B => 
                           mult_21_C243_n1129, CI => mult_21_C243_n1083, CO => 
                           mult_21_C243_n574, S => mult_21_C243_n575);
   mult_21_C243_U356 : ADFULD1 port map( A => mult_21_C243_n588, B => 
                           mult_21_C243_n579, CI => mult_21_C243_n586, CO => 
                           mult_21_C243_n572, S => mult_21_C243_n573);
   mult_21_C243_U355 : ADFULD1 port map( A => mult_21_C243_n577, B => 
                           mult_21_C243_n575, CI => mult_21_C243_n584, CO => 
                           mult_21_C243_n570, S => mult_21_C243_n571);
   mult_21_C243_U354 : ADFULD1 port map( A => mult_21_C243_n582, B => 
                           mult_21_C243_n573, CI => mult_21_C243_n571, CO => 
                           mult_21_C243_n568, S => mult_21_C243_n569);
   mult_21_C243_U353 : ADHALFDL port map( A => mult_21_C243_n1212, B => 
                           mult_21_C243_n947, CO => mult_21_C243_n566, S => 
                           mult_21_C243_n567);
   mult_21_C243_U352 : ADFULD1 port map( A => mult_21_C243_n1104, B => 
                           mult_21_C243_n1044, CI => mult_21_C243_n1182, CO => 
                           mult_21_C243_n564, S => mult_21_C243_n565);
   mult_21_C243_U351 : ADFULD1 port map( A => mult_21_C243_n1154, B => 
                           mult_21_C243_n1082, CI => mult_21_C243_n567, CO => 
                           mult_21_C243_n562, S => mult_21_C243_n563);
   mult_21_C243_U350 : ADFULD1 port map( A => mult_21_C243_n1062, B => 
                           mult_21_C243_n1128, CI => mult_21_C243_n578, CO => 
                           mult_21_C243_n560, S => mult_21_C243_n561);
   mult_21_C243_U349 : ADFULD1 port map( A => mult_21_C243_n574, B => 
                           mult_21_C243_n576, CI => mult_21_C243_n565, CO => 
                           mult_21_C243_n558, S => mult_21_C243_n559);
   mult_21_C243_U348 : ADFULD1 port map( A => mult_21_C243_n561, B => 
                           mult_21_C243_n563, CI => mult_21_C243_n572, CO => 
                           mult_21_C243_n556, S => mult_21_C243_n557);
   mult_21_C243_U347 : ADFULD1 port map( A => mult_21_C243_n570, B => 
                           mult_21_C243_n559, CI => mult_21_C243_n557, CO => 
                           mult_21_C243_n554, S => mult_21_C243_n555);
   mult_21_C243_U346 : ADHALFDL port map( A => mult_21_C243_n566, B => 
                           mult_21_C243_n1211, CO => mult_21_C243_n552, S => 
                           mult_21_C243_n553);
   mult_21_C243_U345 : ADFULD1 port map( A => mult_21_C243_n1043, B => 
                           mult_21_C243_n1103, CI => mult_21_C243_n1061, CO => 
                           mult_21_C243_n550, S => mult_21_C243_n551);
   mult_21_C243_U344 : ADFULD1 port map( A => mult_21_C243_n1181, B => 
                           mult_21_C243_n1081, CI => mult_21_C243_n1127, CO => 
                           mult_21_C243_n548, S => mult_21_C243_n549);
   mult_21_C243_U343 : ADFULD1 port map( A => mult_21_C243_n553, B => 
                           mult_21_C243_n1153, CI => mult_21_C243_n564, CO => 
                           mult_21_C243_n546, S => mult_21_C243_n547);
   mult_21_C243_U342 : ADFULD1 port map( A => mult_21_C243_n560, B => 
                           mult_21_C243_n562, CI => mult_21_C243_n549, CO => 
                           mult_21_C243_n544, S => mult_21_C243_n545);
   mult_21_C243_U341 : ADFULD1 port map( A => mult_21_C243_n547, B => 
                           mult_21_C243_n551, CI => mult_21_C243_n558, CO => 
                           mult_21_C243_n542, S => mult_21_C243_n543);
   mult_21_C243_U340 : ADFULD1 port map( A => mult_21_C243_n556, B => 
                           mult_21_C243_n545, CI => mult_21_C243_n543, CO => 
                           mult_21_C243_n540, S => mult_21_C243_n541);
   mult_21_C243_U339 : ADHALFDL port map( A => mult_21_C243_n1210, B => 
                           mult_21_C243_n946, CO => mult_21_C243_n538, S => 
                           mult_21_C243_n539);
   mult_21_C243_U338 : ADFULD1 port map( A => mult_21_C243_n1102, B => 
                           mult_21_C243_n1026, CI => mult_21_C243_n1180, CO => 
                           mult_21_C243_n536, S => mult_21_C243_n537);
   mult_21_C243_U337 : ADFULD1 port map( A => mult_21_C243_n1042, B => 
                           mult_21_C243_n1060, CI => mult_21_C243_n539, CO => 
                           mult_21_C243_n534, S => mult_21_C243_n535);
   mult_21_C243_U336 : ADFULD1 port map( A => mult_21_C243_n1080, B => 
                           mult_21_C243_n1152, CI => mult_21_C243_n1126, CO => 
                           mult_21_C243_n532, S => mult_21_C243_n533);
   mult_21_C243_U335 : ADFULD1 port map( A => mult_21_C243_n550, B => 
                           mult_21_C243_n552, CI => mult_21_C243_n548, CO => 
                           mult_21_C243_n530, S => mult_21_C243_n531);
   mult_21_C243_U334 : ADFULD1 port map( A => mult_21_C243_n533, B => 
                           mult_21_C243_n537, CI => mult_21_C243_n535, CO => 
                           mult_21_C243_n528, S => mult_21_C243_n529);
   mult_21_C243_U333 : ADFULD1 port map( A => mult_21_C243_n544, B => 
                           mult_21_C243_n546, CI => mult_21_C243_n531, CO => 
                           mult_21_C243_n526, S => mult_21_C243_n527);
   mult_21_C243_U332 : ADFULD1 port map( A => mult_21_C243_n542, B => 
                           mult_21_C243_n529, CI => mult_21_C243_n527, CO => 
                           mult_21_C243_n524, S => mult_21_C243_n525);
   mult_21_C243_U331 : ADHALFDL port map( A => mult_21_C243_n538, B => 
                           mult_21_C243_n1209, CO => mult_21_C243_n522, S => 
                           mult_21_C243_n523);
   mult_21_C243_U330 : ADFULD1 port map( A => mult_21_C243_n1179, B => 
                           mult_21_C243_n1079, CI => mult_21_C243_n1151, CO => 
                           mult_21_C243_n520, S => mult_21_C243_n521);
   mult_21_C243_U329 : ADFULD1 port map( A => mult_21_C243_n1025, B => 
                           mult_21_C243_n1041, CI => mult_21_C243_n1059, CO => 
                           mult_21_C243_n518, S => mult_21_C243_n519);
   mult_21_C243_U328 : ADFULD1 port map( A => mult_21_C243_n1101, B => 
                           mult_21_C243_n1125, CI => mult_21_C243_n523, CO => 
                           mult_21_C243_n516, S => mult_21_C243_n517);
   mult_21_C243_U327 : ADFULD1 port map( A => mult_21_C243_n534, B => 
                           mult_21_C243_n536, CI => mult_21_C243_n532, CO => 
                           mult_21_C243_n514, S => mult_21_C243_n515);
   mult_21_C243_U326 : ADFULD1 port map( A => mult_21_C243_n521, B => 
                           mult_21_C243_n519, CI => mult_21_C243_n517, CO => 
                           mult_21_C243_n512, S => mult_21_C243_n513);
   mult_21_C243_U325 : ADFULD1 port map( A => mult_21_C243_n528, B => 
                           mult_21_C243_n530, CI => mult_21_C243_n515, CO => 
                           mult_21_C243_n510, S => mult_21_C243_n511);
   mult_21_C243_U324 : ADFULD1 port map( A => mult_21_C243_n526, B => 
                           mult_21_C243_n513, CI => mult_21_C243_n511, CO => 
                           mult_21_C243_n508, S => mult_21_C243_n509);
   mult_21_C243_U323 : ADHALFDL port map( A => mult_21_C243_n1208, B => 
                           mult_21_C243_n945, CO => mult_21_C243_n506, S => 
                           mult_21_C243_n507);
   mult_21_C243_U322 : ADFULD1 port map( A => mult_21_C243_n1078, B => 
                           mult_21_C243_n1010, CI => mult_21_C243_n1024, CO => 
                           mult_21_C243_n504, S => mult_21_C243_n505);
   mult_21_C243_U321 : ADFULD1 port map( A => mult_21_C243_n1178, B => 
                           mult_21_C243_n1100, CI => mult_21_C243_n507, CO => 
                           mult_21_C243_n502, S => mult_21_C243_n503);
   mult_21_C243_U320 : ADFULD1 port map( A => mult_21_C243_n1040, B => 
                           mult_21_C243_n1150, CI => mult_21_C243_n1058, CO => 
                           mult_21_C243_n500, S => mult_21_C243_n501);
   mult_21_C243_U319 : ADFULD1 port map( A => mult_21_C243_n522, B => 
                           mult_21_C243_n1124, CI => mult_21_C243_n520, CO => 
                           mult_21_C243_n498, S => mult_21_C243_n499);
   mult_21_C243_U318 : ADFULD1 port map( A => mult_21_C243_n505, B => 
                           mult_21_C243_n518, CI => mult_21_C243_n501, CO => 
                           mult_21_C243_n496, S => mult_21_C243_n497);
   mult_21_C243_U317 : ADFULD1 port map( A => mult_21_C243_n516, B => 
                           mult_21_C243_n503, CI => mult_21_C243_n514, CO => 
                           mult_21_C243_n494, S => mult_21_C243_n495);
   mult_21_C243_U316 : ADFULD1 port map( A => mult_21_C243_n497, B => 
                           mult_21_C243_n499, CI => mult_21_C243_n512, CO => 
                           mult_21_C243_n492, S => mult_21_C243_n493);
   mult_21_C243_U315 : ADFULD1 port map( A => mult_21_C243_n510, B => 
                           mult_21_C243_n495, CI => mult_21_C243_n493, CO => 
                           mult_21_C243_n490, S => mult_21_C243_n491);
   mult_21_C243_U314 : ADHALFDL port map( A => mult_21_C243_n506, B => 
                           mult_21_C243_n1207, CO => mult_21_C243_n488, S => 
                           mult_21_C243_n489);
   mult_21_C243_U313 : ADFULD1 port map( A => mult_21_C243_n1009, B => 
                           mult_21_C243_n1077, CI => mult_21_C243_n1023, CO => 
                           mult_21_C243_n486, S => mult_21_C243_n487);
   mult_21_C243_U312 : ADFULD1 port map( A => mult_21_C243_n1177, B => 
                           mult_21_C243_n1099, CI => mult_21_C243_n1039, CO => 
                           mult_21_C243_n484, S => mult_21_C243_n485);
   mult_21_C243_U311 : ADFULD1 port map( A => mult_21_C243_n1057, B => 
                           mult_21_C243_n1149, CI => mult_21_C243_n1123, CO => 
                           mult_21_C243_n482, S => mult_21_C243_n483);
   mult_21_C243_U310 : ADFULD1 port map( A => mult_21_C243_n504, B => 
                           mult_21_C243_n489, CI => mult_21_C243_n502, CO => 
                           mult_21_C243_n480, S => mult_21_C243_n481);
   mult_21_C243_U309 : ADFULD1 port map( A => mult_21_C243_n483, B => 
                           mult_21_C243_n500, CI => mult_21_C243_n485, CO => 
                           mult_21_C243_n478, S => mult_21_C243_n479);
   mult_21_C243_U308 : ADFULD1 port map( A => mult_21_C243_n498, B => 
                           mult_21_C243_n487, CI => mult_21_C243_n496, CO => 
                           mult_21_C243_n476, S => mult_21_C243_n477);
   mult_21_C243_U307 : ADFULD1 port map( A => mult_21_C243_n479, B => 
                           mult_21_C243_n481, CI => mult_21_C243_n494, CO => 
                           mult_21_C243_n474, S => mult_21_C243_n475);
   mult_21_C243_U306 : ADFULD1 port map( A => mult_21_C243_n492, B => 
                           mult_21_C243_n477, CI => mult_21_C243_n475, CO => 
                           mult_21_C243_n472, S => mult_21_C243_n473);
   mult_21_C243_U305 : ADHALFDL port map( A => mult_21_C243_n1206, B => 
                           mult_21_C243_n944, CO => mult_21_C243_n470, S => 
                           mult_21_C243_n471);
   mult_21_C243_U304 : ADFULD1 port map( A => mult_21_C243_n1076, B => 
                           mult_21_C243_n996, CI => mult_21_C243_n1176, CO => 
                           mult_21_C243_n468, S => mult_21_C243_n469);
   mult_21_C243_U303 : ADFULD1 port map( A => mult_21_C243_n1008, B => 
                           mult_21_C243_n1038, CI => mult_21_C243_n471, CO => 
                           mult_21_C243_n466, S => mult_21_C243_n467);
   mult_21_C243_U302 : ADFULD1 port map( A => mult_21_C243_n1022, B => 
                           mult_21_C243_n1148, CI => mult_21_C243_n1056, CO => 
                           mult_21_C243_n464, S => mult_21_C243_n465);
   mult_21_C243_U301 : ADFULD1 port map( A => mult_21_C243_n1098, B => 
                           mult_21_C243_n1122, CI => mult_21_C243_n488, CO => 
                           mult_21_C243_n462, S => mult_21_C243_n463);
   mult_21_C243_U300 : ADFULD1 port map( A => mult_21_C243_n482, B => 
                           mult_21_C243_n486, CI => mult_21_C243_n484, CO => 
                           mult_21_C243_n460, S => mult_21_C243_n461);
   mult_21_C243_U299 : ADFULD1 port map( A => mult_21_C243_n465, B => 
                           mult_21_C243_n469, CI => mult_21_C243_n467, CO => 
                           mult_21_C243_n458, S => mult_21_C243_n459);
   mult_21_C243_U298 : ADFULD1 port map( A => mult_21_C243_n480, B => 
                           mult_21_C243_n463, CI => mult_21_C243_n478, CO => 
                           mult_21_C243_n456, S => mult_21_C243_n457);
   mult_21_C243_U297 : ADFULD1 port map( A => mult_21_C243_n459, B => 
                           mult_21_C243_n461, CI => mult_21_C243_n476, CO => 
                           mult_21_C243_n454, S => mult_21_C243_n455);
   mult_21_C243_U296 : ADFULD1 port map( A => mult_21_C243_n474, B => 
                           mult_21_C243_n457, CI => mult_21_C243_n455, CO => 
                           mult_21_C243_n452, S => mult_21_C243_n453);
   mult_21_C243_U295 : ADHALFDL port map( A => mult_21_C243_n470, B => 
                           mult_21_C243_n1205, CO => mult_21_C243_n450, S => 
                           mult_21_C243_n451);
   mult_21_C243_U294 : ADFULD1 port map( A => mult_21_C243_n1175, B => 
                           mult_21_C243_n1055, CI => mult_21_C243_n1147, CO => 
                           mult_21_C243_n448, S => mult_21_C243_n449);
   mult_21_C243_U293 : ADFULD1 port map( A => mult_21_C243_n1121, B => 
                           mult_21_C243_n1021, CI => mult_21_C243_n1097, CO => 
                           mult_21_C243_n446, S => mult_21_C243_n447);
   mult_21_C243_U292 : ADFULD1 port map( A => mult_21_C243_n995, B => 
                           mult_21_C243_n1075, CI => mult_21_C243_n1007, CO => 
                           mult_21_C243_n444, S => mult_21_C243_n445);
   mult_21_C243_U291 : ADFULD1 port map( A => mult_21_C243_n451, B => 
                           mult_21_C243_n1037, CI => mult_21_C243_n468, CO => 
                           mult_21_C243_n442, S => mult_21_C243_n443);
   mult_21_C243_U290 : ADFULD1 port map( A => mult_21_C243_n464, B => 
                           mult_21_C243_n466, CI => mult_21_C243_n462, CO => 
                           mult_21_C243_n440, S => mult_21_C243_n441);
   mult_21_C243_U289 : ADFULD1 port map( A => mult_21_C243_n449, B => 
                           mult_21_C243_n445, CI => mult_21_C243_n447, CO => 
                           mult_21_C243_n438, S => mult_21_C243_n439);
   mult_21_C243_U288 : ADFULD1 port map( A => mult_21_C243_n443, B => 
                           mult_21_C243_n460, CI => mult_21_C243_n458, CO => 
                           mult_21_C243_n436, S => mult_21_C243_n437);
   mult_21_C243_U287 : ADFULD1 port map( A => mult_21_C243_n439, B => 
                           mult_21_C243_n441, CI => mult_21_C243_n456, CO => 
                           mult_21_C243_n434, S => mult_21_C243_n435);
   mult_21_C243_U286 : ADFULD1 port map( A => mult_21_C243_n454, B => 
                           mult_21_C243_n437, CI => mult_21_C243_n435, CO => 
                           mult_21_C243_n432, S => mult_21_C243_n433);
   mult_21_C243_U285 : ADHALFDL port map( A => mult_21_C243_n1204, B => 
                           mult_21_C243_n943, CO => mult_21_C243_n430, S => 
                           mult_21_C243_n431);
   mult_21_C243_U284 : ADFULD1 port map( A => mult_21_C243_n1054, B => 
                           mult_21_C243_n984, CI => mult_21_C243_n994, CO => 
                           mult_21_C243_n428, S => mult_21_C243_n429);
   mult_21_C243_U283 : ADFULD1 port map( A => mult_21_C243_n1174, B => 
                           mult_21_C243_n1036, CI => mult_21_C243_n431, CO => 
                           mult_21_C243_n426, S => mult_21_C243_n427);
   mult_21_C243_U282 : ADFULD1 port map( A => mult_21_C243_n1006, B => 
                           mult_21_C243_n1146, CI => mult_21_C243_n1020, CO => 
                           mult_21_C243_n424, S => mult_21_C243_n425);
   mult_21_C243_U281 : ADFULD1 port map( A => mult_21_C243_n1074, B => 
                           mult_21_C243_n1120, CI => mult_21_C243_n1096, CO => 
                           mult_21_C243_n422, S => mult_21_C243_n423);
   mult_21_C243_U280 : ADFULD1 port map( A => mult_21_C243_n448, B => 
                           mult_21_C243_n450, CI => mult_21_C243_n446, CO => 
                           mult_21_C243_n420, S => mult_21_C243_n421);
   mult_21_C243_U279 : ADFULD1 port map( A => mult_21_C243_n429, B => 
                           mult_21_C243_n444, CI => mult_21_C243_n423, CO => 
                           mult_21_C243_n418, S => mult_21_C243_n419);
   mult_21_C243_U278 : ADFULD1 port map( A => mult_21_C243_n427, B => 
                           mult_21_C243_n425, CI => mult_21_C243_n442, CO => 
                           mult_21_C243_n416, S => mult_21_C243_n417);
   mult_21_C243_U277 : ADFULD1 port map( A => mult_21_C243_n421, B => 
                           mult_21_C243_n440, CI => mult_21_C243_n438, CO => 
                           mult_21_C243_n414, S => mult_21_C243_n415);
   mult_21_C243_U276 : ADFULD1 port map( A => mult_21_C243_n417, B => 
                           mult_21_C243_n419, CI => mult_21_C243_n436, CO => 
                           mult_21_C243_n412, S => mult_21_C243_n413);
   mult_21_C243_U275 : ADFULD1 port map( A => mult_21_C243_n434, B => 
                           mult_21_C243_n415, CI => mult_21_C243_n413, CO => 
                           mult_21_C243_n410, S => mult_21_C243_n411);
   mult_21_C243_U274 : ADHALFDL port map( A => mult_21_C243_n430, B => 
                           mult_21_C243_n1203, CO => mult_21_C243_n408, S => 
                           mult_21_C243_n409);
   mult_21_C243_U273 : ADFULD1 port map( A => mult_21_C243_n983, B => 
                           mult_21_C243_n1053, CI => mult_21_C243_n993, CO => 
                           mult_21_C243_n406, S => mult_21_C243_n407);
   mult_21_C243_U272 : ADFULD1 port map( A => mult_21_C243_n1173, B => 
                           mult_21_C243_n1035, CI => mult_21_C243_n1145, CO => 
                           mult_21_C243_n404, S => mult_21_C243_n405);
   mult_21_C243_U271 : ADFULD1 port map( A => mult_21_C243_n1005, B => 
                           mult_21_C243_n1119, CI => mult_21_C243_n1019, CO => 
                           mult_21_C243_n402, S => mult_21_C243_n403);
   mult_21_C243_U270 : ADFULD1 port map( A => mult_21_C243_n1073, B => 
                           mult_21_C243_n1095, CI => mult_21_C243_n409, CO => 
                           mult_21_C243_n400, S => mult_21_C243_n401);
   mult_21_C243_U269 : ADFULD1 port map( A => mult_21_C243_n426, B => 
                           mult_21_C243_n428, CI => mult_21_C243_n422, CO => 
                           mult_21_C243_n398, S => mult_21_C243_n399);
   mult_21_C243_U268 : ADFULD1 port map( A => mult_21_C243_n403, B => 
                           mult_21_C243_n424, CI => mult_21_C243_n405, CO => 
                           mult_21_C243_n396, S => mult_21_C243_n397);
   mult_21_C243_U267 : ADFULD1 port map( A => mult_21_C243_n401, B => 
                           mult_21_C243_n407, CI => mult_21_C243_n420, CO => 
                           mult_21_C243_n394, S => mult_21_C243_n395);
   mult_21_C243_U266 : ADFULD1 port map( A => mult_21_C243_n399, B => 
                           mult_21_C243_n418, CI => mult_21_C243_n416, CO => 
                           mult_21_C243_n392, S => mult_21_C243_n393);
   mult_21_C243_U265 : ADFULD1 port map( A => mult_21_C243_n395, B => 
                           mult_21_C243_n397, CI => mult_21_C243_n414, CO => 
                           mult_21_C243_n390, S => mult_21_C243_n391);
   mult_21_C243_U264 : ADFULD1 port map( A => mult_21_C243_n412, B => 
                           mult_21_C243_n393, CI => mult_21_C243_n391, CO => 
                           mult_21_C243_n388, S => mult_21_C243_n389);
   mult_21_C243_U263 : ADHALFDL port map( A => mult_21_C243_n1202, B => 
                           mult_21_C243_n942, CO => mult_21_C243_n386, S => 
                           mult_21_C243_n387);
   mult_21_C243_U262 : ADFULD1 port map( A => mult_21_C243_n1052, B => 
                           mult_21_C243_n974, CI => mult_21_C243_n1172, CO => 
                           mult_21_C243_n384, S => mult_21_C243_n385);
   mult_21_C243_U261 : ADFULD1 port map( A => mult_21_C243_n982, B => 
                           mult_21_C243_n1018, CI => mult_21_C243_n387, CO => 
                           mult_21_C243_n382, S => mult_21_C243_n383);
   mult_21_C243_U260 : ADFULD1 port map( A => mult_21_C243_n992, B => 
                           mult_21_C243_n1144, CI => mult_21_C243_n1118, CO => 
                           mult_21_C243_n380, S => mult_21_C243_n381);
   mult_21_C243_U259 : ADFULD1 port map( A => mult_21_C243_n1004, B => 
                           mult_21_C243_n1094, CI => mult_21_C243_n1034, CO => 
                           mult_21_C243_n378, S => mult_21_C243_n379);
   mult_21_C243_U258 : ADFULD1 port map( A => mult_21_C243_n408, B => 
                           mult_21_C243_n1072, CI => mult_21_C243_n406, CO => 
                           mult_21_C243_n376, S => mult_21_C243_n377);
   mult_21_C243_U257 : ADFULD1 port map( A => mult_21_C243_n402, B => 
                           mult_21_C243_n404, CI => mult_21_C243_n385, CO => 
                           mult_21_C243_n374, S => mult_21_C243_n375);
   mult_21_C243_U256 : ADFULD1 port map( A => mult_21_C243_n383, B => 
                           mult_21_C243_n379, CI => mult_21_C243_n381, CO => 
                           mult_21_C243_n372, S => mult_21_C243_n373);
   mult_21_C243_U255 : ADFULD1 port map( A => mult_21_C243_n398, B => 
                           mult_21_C243_n400, CI => mult_21_C243_n377, CO => 
                           mult_21_C243_n370, S => mult_21_C243_n371);
   mult_21_C243_U254 : ADFULD1 port map( A => mult_21_C243_n375, B => 
                           mult_21_C243_n396, CI => mult_21_C243_n373, CO => 
                           mult_21_C243_n368, S => mult_21_C243_n369);
   mult_21_C243_U253 : ADFULD1 port map( A => mult_21_C243_n371, B => 
                           mult_21_C243_n394, CI => mult_21_C243_n392, CO => 
                           mult_21_C243_n366, S => mult_21_C243_n367);
   mult_21_C243_U252 : ADFULD1 port map( A => mult_21_C243_n390, B => 
                           mult_21_C243_n369, CI => mult_21_C243_n367, CO => 
                           mult_21_C243_n364, S => mult_21_C243_n365);
   mult_21_C243_U251 : ADHALFDL port map( A => mult_21_C243_n386, B => 
                           mult_21_C243_n1201, CO => mult_21_C243_n362, S => 
                           mult_21_C243_n363);
   mult_21_C243_U250 : ADFULD1 port map( A => mult_21_C243_n1171, B => 
                           mult_21_C243_n1051, CI => mult_21_C243_n1143, CO => 
                           mult_21_C243_n360, S => mult_21_C243_n361);
   mult_21_C243_U249 : ADFULD1 port map( A => mult_21_C243_n973, B => 
                           mult_21_C243_n1003, CI => mult_21_C243_n981, CO => 
                           mult_21_C243_n358, S => mult_21_C243_n359);
   mult_21_C243_U248 : ADFULD1 port map( A => mult_21_C243_n991, B => 
                           mult_21_C243_n1117, CI => mult_21_C243_n1017, CO => 
                           mult_21_C243_n356, S => mult_21_C243_n357);
   mult_21_C243_U247 : ADFULD1 port map( A => mult_21_C243_n1033, B => 
                           mult_21_C243_n1093, CI => mult_21_C243_n1071, CO => 
                           mult_21_C243_n354, S => mult_21_C243_n355);
   mult_21_C243_U246 : ADFULD1 port map( A => mult_21_C243_n384, B => 
                           mult_21_C243_n363, CI => mult_21_C243_n382, CO => 
                           mult_21_C243_n352, S => mult_21_C243_n353);
   mult_21_C243_U245 : ADFULD1 port map( A => mult_21_C243_n378, B => 
                           mult_21_C243_n380, CI => mult_21_C243_n355, CO => 
                           mult_21_C243_n350, S => mult_21_C243_n351);
   mult_21_C243_U244 : ADFULD1 port map( A => mult_21_C243_n361, B => 
                           mult_21_C243_n357, CI => mult_21_C243_n359, CO => 
                           mult_21_C243_n348, S => mult_21_C243_n349);
   mult_21_C243_U243 : ADFULD1 port map( A => mult_21_C243_n374, B => 
                           mult_21_C243_n376, CI => mult_21_C243_n353, CO => 
                           mult_21_C243_n346, S => mult_21_C243_n347);
   mult_21_C243_U242 : ADFULD1 port map( A => mult_21_C243_n351, B => 
                           mult_21_C243_n372, CI => mult_21_C243_n349, CO => 
                           mult_21_C243_n344, S => mult_21_C243_n345);
   mult_21_C243_U241 : ADFULD1 port map( A => mult_21_C243_n347, B => 
                           mult_21_C243_n370, CI => mult_21_C243_n368, CO => 
                           mult_21_C243_n342, S => mult_21_C243_n343);
   mult_21_C243_U240 : ADFULD1 port map( A => mult_21_C243_n366, B => 
                           mult_21_C243_n345, CI => mult_21_C243_n343, CO => 
                           mult_21_C243_n340, S => mult_21_C243_n341);
   mult_21_C243_U239 : ADHALFDL port map( A => mult_21_C243_n1200, B => 
                           mult_21_C243_n941, CO => mult_21_C243_n338, S => 
                           mult_21_C243_n339);
   mult_21_C243_U238 : ADFULD1 port map( A => mult_21_C243_n1050, B => 
                           mult_21_C243_n966, CI => mult_21_C243_n972, CO => 
                           mult_21_C243_n336, S => mult_21_C243_n337);
   mult_21_C243_U237 : ADFULD1 port map( A => mult_21_C243_n980, B => 
                           mult_21_C243_n1032, CI => mult_21_C243_n339, CO => 
                           mult_21_C243_n334, S => mult_21_C243_n335);
   mult_21_C243_U236 : ADFULD1 port map( A => mult_21_C243_n990, B => 
                           mult_21_C243_n1170, CI => mult_21_C243_n1002, CO => 
                           mult_21_C243_n332, S => mult_21_C243_n333);
   mult_21_C243_U235 : ADFULD1 port map( A => mult_21_C243_n1016, B => 
                           mult_21_C243_n1142, CI => mult_21_C243_n1070, CO => 
                           mult_21_C243_n330, S => mult_21_C243_n331);
   mult_21_C243_U234 : ADFULD1 port map( A => mult_21_C243_n1092, B => 
                           mult_21_C243_n1116, CI => mult_21_C243_n362, CO => 
                           mult_21_C243_n328, S => mult_21_C243_n329);
   mult_21_C243_U233 : ADFULD1 port map( A => mult_21_C243_n354, B => 
                           mult_21_C243_n360, CI => mult_21_C243_n356, CO => 
                           mult_21_C243_n326, S => mult_21_C243_n327);
   mult_21_C243_U232 : ADFULD1 port map( A => mult_21_C243_n337, B => 
                           mult_21_C243_n358, CI => mult_21_C243_n331, CO => 
                           mult_21_C243_n324, S => mult_21_C243_n325);
   mult_21_C243_U231 : ADFULD1 port map( A => mult_21_C243_n333, B => 
                           mult_21_C243_n335, CI => mult_21_C243_n329, CO => 
                           mult_21_C243_n322, S => mult_21_C243_n323);
   mult_21_C243_U230 : ADFULD1 port map( A => mult_21_C243_n350, B => 
                           mult_21_C243_n352, CI => mult_21_C243_n348, CO => 
                           mult_21_C243_n320, S => mult_21_C243_n321);
   mult_21_C243_U229 : ADFULD1 port map( A => mult_21_C243_n325, B => 
                           mult_21_C243_n327, CI => mult_21_C243_n323, CO => 
                           mult_21_C243_n318, S => mult_21_C243_n319);
   mult_21_C243_U228 : ADFULD1 port map( A => mult_21_C243_n344, B => 
                           mult_21_C243_n346, CI => mult_21_C243_n321, CO => 
                           mult_21_C243_n316, S => mult_21_C243_n317);
   mult_21_C243_U227 : ADFULD1 port map( A => mult_21_C243_n342, B => 
                           mult_21_C243_n319, CI => mult_21_C243_n317, CO => 
                           mult_21_C243_n314, S => mult_21_C243_n315);
   mult_21_C243_U226 : ADHALFDL port map( A => mult_21_C243_n338, B => 
                           mult_21_C243_n1199, CO => mult_21_C243_n312, S => 
                           mult_21_C243_n313);
   mult_21_C243_U225 : ADFULD1 port map( A => mult_21_C243_n965, B => 
                           mult_21_C243_n1031, CI => mult_21_C243_n971, CO => 
                           mult_21_C243_n310, S => mult_21_C243_n311);
   mult_21_C243_U224 : ADFULD1 port map( A => mult_21_C243_n979, B => 
                           mult_21_C243_n1049, CI => mult_21_C243_n1169, CO => 
                           mult_21_C243_n308, S => mult_21_C243_n309);
   mult_21_C243_U223 : ADFULD1 port map( A => mult_21_C243_n1141, B => 
                           mult_21_C243_n1001, CI => mult_21_C243_n989, CO => 
                           mult_21_C243_n306, S => mult_21_C243_n307);
   mult_21_C243_U222 : ADFULD1 port map( A => mult_21_C243_n1015, B => 
                           mult_21_C243_n1115, CI => mult_21_C243_n1069, CO => 
                           mult_21_C243_n304, S => mult_21_C243_n305);
   mult_21_C243_U221 : ADFULD1 port map( A => mult_21_C243_n313, B => 
                           mult_21_C243_n1091, CI => mult_21_C243_n336, CO => 
                           mult_21_C243_n302, S => mult_21_C243_n303);
   mult_21_C243_U220 : ADFULD1 port map( A => mult_21_C243_n332, B => 
                           mult_21_C243_n330, CI => mult_21_C243_n334, CO => 
                           mult_21_C243_n300, S => mult_21_C243_n301);
   mult_21_C243_U219 : ADFULD1 port map( A => mult_21_C243_n305, B => 
                           mult_21_C243_n328, CI => mult_21_C243_n311, CO => 
                           mult_21_C243_n298, S => mult_21_C243_n299);
   mult_21_C243_U218 : ADFULD1 port map( A => mult_21_C243_n307, B => 
                           mult_21_C243_n309, CI => mult_21_C243_n326, CO => 
                           mult_21_C243_n296, S => mult_21_C243_n297);
   mult_21_C243_U217 : ADFULD1 port map( A => mult_21_C243_n324, B => 
                           mult_21_C243_n303, CI => mult_21_C243_n301, CO => 
                           mult_21_C243_n294, S => mult_21_C243_n295);
   mult_21_C243_U216 : ADFULD1 port map( A => mult_21_C243_n299, B => 
                           mult_21_C243_n322, CI => mult_21_C243_n320, CO => 
                           mult_21_C243_n292, S => mult_21_C243_n293);
   mult_21_C243_U215 : ADFULD1 port map( A => mult_21_C243_n318, B => 
                           mult_21_C243_n297, CI => mult_21_C243_n295, CO => 
                           mult_21_C243_n290, S => mult_21_C243_n291);
   mult_21_C243_U214 : ADFULD1 port map( A => mult_21_C243_n316, B => 
                           mult_21_C243_n293, CI => mult_21_C243_n291, CO => 
                           mult_21_C243_n288, S => mult_21_C243_n289);
   mult_21_C243_U213 : ADHALFDL port map( A => mult_21_C243_n1198, B => 
                           mult_21_C243_n940, CO => mult_21_C243_n286, S => 
                           mult_21_C243_n287);
   mult_21_C243_U212 : ADFULD1 port map( A => mult_21_C243_n1030, B => 
                           mult_21_C243_n960, CI => mult_21_C243_n1168, CO => 
                           mult_21_C243_n284, S => mult_21_C243_n285);
   mult_21_C243_U211 : ADFULD1 port map( A => mult_21_C243_n1140, B => 
                           mult_21_C243_n1000, CI => mult_21_C243_n287, CO => 
                           mult_21_C243_n282, S => mult_21_C243_n283);
   mult_21_C243_U210 : ADFULD1 port map( A => mult_21_C243_n964, B => 
                           mult_21_C243_n1114, CI => mult_21_C243_n970, CO => 
                           mult_21_C243_n280, S => mult_21_C243_n281);
   mult_21_C243_U209 : ADFULD1 port map( A => mult_21_C243_n978, B => 
                           mult_21_C243_n1090, CI => mult_21_C243_n988, CO => 
                           mult_21_C243_n278, S => mult_21_C243_n279);
   mult_21_C243_U208 : ADFULD1 port map( A => mult_21_C243_n1014, B => 
                           mult_21_C243_n1068, CI => mult_21_C243_n1048, CO => 
                           mult_21_C243_n276, S => mult_21_C243_n277);
   mult_21_C243_U207 : ADFULD1 port map( A => mult_21_C243_n304, B => 
                           mult_21_C243_n312, CI => mult_21_C243_n306, CO => 
                           mult_21_C243_n274, S => mult_21_C243_n275);
   mult_21_C243_U206 : ADFULD1 port map( A => mult_21_C243_n310, B => 
                           mult_21_C243_n308, CI => mult_21_C243_n285, CO => 
                           mult_21_C243_n272, S => mult_21_C243_n273);
   mult_21_C243_U205 : ADFULD1 port map( A => mult_21_C243_n283, B => 
                           mult_21_C243_n277, CI => mult_21_C243_n279, CO => 
                           mult_21_C243_n270, S => mult_21_C243_n271);
   mult_21_C243_U204 : ADFULD1 port map( A => mult_21_C243_n302, B => 
                           mult_21_C243_n281, CI => mult_21_C243_n300, CO => 
                           mult_21_C243_n268, S => mult_21_C243_n269);
   mult_21_C243_U203 : ADFULD1 port map( A => mult_21_C243_n275, B => 
                           mult_21_C243_n298, CI => mult_21_C243_n273, CO => 
                           mult_21_C243_n266, S => mult_21_C243_n267);
   mult_21_C243_U202 : ADFULD1 port map( A => mult_21_C243_n296, B => 
                           mult_21_C243_n271, CI => mult_21_C243_n269, CO => 
                           mult_21_C243_n264, S => mult_21_C243_n265);
   mult_21_C243_U201 : ADFULD1 port map( A => mult_21_C243_n267, B => 
                           mult_21_C243_n294, CI => mult_21_C243_n292, CO => 
                           mult_21_C243_n262, S => mult_21_C243_n263);
   mult_21_C243_U200 : ADFULD1 port map( A => mult_21_C243_n290, B => 
                           mult_21_C243_n265, CI => mult_21_C243_n263, CO => 
                           mult_21_C243_n260, S => mult_21_C243_n261);
   mult_21_C243_U199 : ADHALFDL port map( A => mult_21_C243_n286, B => 
                           mult_21_C243_n1197, CO => mult_21_C243_n258, S => 
                           mult_21_C243_n259);
   mult_21_C243_U198 : ADFULD1 port map( A => mult_21_C243_n1167, B => 
                           mult_21_C243_n1029, CI => mult_21_C243_n1139, CO => 
                           mult_21_C243_n256, S => mult_21_C243_n257);
   mult_21_C243_U197 : ADFULD1 port map( A => mult_21_C243_n1113, B => 
                           mult_21_C243_n987, CI => mult_21_C243_n1089, CO => 
                           mult_21_C243_n254, S => mult_21_C243_n255);
   mult_21_C243_U196 : ADFULD1 port map( A => mult_21_C243_n959, B => 
                           mult_21_C243_n969, CI => mult_21_C243_n963, CO => 
                           mult_21_C243_n252, S => mult_21_C243_n253);
   mult_21_C243_U195 : ADFULD1 port map( A => mult_21_C243_n977, B => 
                           mult_21_C243_n1067, CI => mult_21_C243_n999, CO => 
                           mult_21_C243_n250, S => mult_21_C243_n251);
   mult_21_C243_U194 : ADFULD1 port map( A => mult_21_C243_n1047, B => 
                           mult_21_C243_n1013, CI => mult_21_C243_n259, CO => 
                           mult_21_C243_n248, S => mult_21_C243_n249);
   mult_21_C243_U193 : ADFULD1 port map( A => mult_21_C243_n278, B => 
                           mult_21_C243_n284, CI => mult_21_C243_n282, CO => 
                           mult_21_C243_n246, S => mult_21_C243_n247);
   mult_21_C243_U192 : ADFULD1 port map( A => mult_21_C243_n280, B => 
                           mult_21_C243_n276, CI => mult_21_C243_n251, CO => 
                           mult_21_C243_n244, S => mult_21_C243_n245);
   mult_21_C243_U191 : ADFULD1 port map( A => mult_21_C243_n253, B => 
                           mult_21_C243_n255, CI => mult_21_C243_n257, CO => 
                           mult_21_C243_n242, S => mult_21_C243_n243);
   mult_21_C243_U190 : ADFULD1 port map( A => mult_21_C243_n274, B => 
                           mult_21_C243_n249, CI => mult_21_C243_n272, CO => 
                           mult_21_C243_n240, S => mult_21_C243_n241);
   mult_21_C243_U189 : ADFULD1 port map( A => mult_21_C243_n270, B => 
                           mult_21_C243_n247, CI => mult_21_C243_n245, CO => 
                           mult_21_C243_n238, S => mult_21_C243_n239);
   mult_21_C243_U188 : ADFULD1 port map( A => mult_21_C243_n268, B => 
                           mult_21_C243_n243, CI => mult_21_C243_n241, CO => 
                           mult_21_C243_n236, S => mult_21_C243_n237);
   mult_21_C243_U187 : ADFULD1 port map( A => mult_21_C243_n239, B => 
                           mult_21_C243_n266, CI => mult_21_C243_n264, CO => 
                           mult_21_C243_n234, S => mult_21_C243_n235);
   mult_21_C243_U186 : ADFULD1 port map( A => mult_21_C243_n262, B => 
                           mult_21_C243_n237, CI => mult_21_C243_n235, CO => 
                           mult_21_C243_n232, S => mult_21_C243_n233);
   mult_21_C243_U185 : ADHALFDL port map( A => mult_21_C243_n1196, B => 
                           mult_21_C243_n939, CO => mult_21_C243_n230, S => 
                           mult_21_C243_n231);
   mult_21_C243_U184 : ADFULD1 port map( A => mult_21_C243_n1028, B => 
                           mult_21_C243_n956, CI => mult_21_C243_n958, CO => 
                           mult_21_C243_n228, S => mult_21_C243_n229);
   mult_21_C243_U183 : ADFULD1 port map( A => mult_21_C243_n1166, B => 
                           mult_21_C243_n1012, CI => mult_21_C243_n231, CO => 
                           mult_21_C243_n226, S => mult_21_C243_n227);
   mult_21_C243_U182 : ADFULD1 port map( A => mult_21_C243_n962, B => 
                           mult_21_C243_n1138, CI => mult_21_C243_n968, CO => 
                           mult_21_C243_n224, S => mult_21_C243_n225);
   mult_21_C243_U181 : ADFULD1 port map( A => mult_21_C243_n986, B => 
                           mult_21_C243_n976, CI => mult_21_C243_n998, CO => 
                           mult_21_C243_n222, S => mult_21_C243_n223);
   mult_21_C243_U180 : ADFULD1 port map( A => mult_21_C243_n1046, B => 
                           mult_21_C243_n1112, CI => mult_21_C243_n1066, CO => 
                           mult_21_C243_n220, S => mult_21_C243_n221);
   mult_21_C243_U179 : ADFULD1 port map( A => mult_21_C243_n258, B => 
                           mult_21_C243_n1088, CI => mult_21_C243_n250, CO => 
                           mult_21_C243_n218, S => mult_21_C243_n219);
   mult_21_C243_U178 : ADFULD1 port map( A => mult_21_C243_n256, B => 
                           mult_21_C243_n252, CI => mult_21_C243_n254, CO => 
                           mult_21_C243_n216, S => mult_21_C243_n217);
   mult_21_C243_U177 : ADFULD1 port map( A => mult_21_C243_n221, B => 
                           mult_21_C243_n229, CI => mult_21_C243_n227, CO => 
                           mult_21_C243_n214, S => mult_21_C243_n215);
   mult_21_C243_U176 : ADFULD1 port map( A => mult_21_C243_n225, B => 
                           mult_21_C243_n223, CI => mult_21_C243_n248, CO => 
                           mult_21_C243_n212, S => mult_21_C243_n213);
   mult_21_C243_U175 : ADFULD1 port map( A => mult_21_C243_n244, B => 
                           mult_21_C243_n246, CI => mult_21_C243_n219, CO => 
                           mult_21_C243_n210, S => mult_21_C243_n211);
   mult_21_C243_U174 : ADFULD1 port map( A => mult_21_C243_n217, B => 
                           mult_21_C243_n242, CI => mult_21_C243_n215, CO => 
                           mult_21_C243_n208, S => mult_21_C243_n209);
   mult_21_C243_U173 : ADFULD1 port map( A => mult_21_C243_n240, B => 
                           mult_21_C243_n213, CI => mult_21_C243_n238, CO => 
                           mult_21_C243_n206, S => mult_21_C243_n207);
   mult_21_C243_U172 : ADFULD1 port map( A => mult_21_C243_n209, B => 
                           mult_21_C243_n211, CI => mult_21_C243_n236, CO => 
                           mult_21_C243_n204, S => mult_21_C243_n205);
   mult_21_C243_U171 : ADFULD1 port map( A => mult_21_C243_n234, B => 
                           mult_21_C243_n207, CI => mult_21_C243_n205, CO => 
                           mult_21_C243_n202, S => mult_21_C243_n203);
   mult_21_C243_U155 : ADHALFDL port map( A => mult_21_C243_n1226, B => N2946, 
                           CO => mult_21_C243_n186, S => N3265);
   mult_21_C243_U154 : ADHALFDL port map( A => mult_21_C243_n186, B => 
                           mult_21_C243_n1225, CO => mult_21_C243_n185, S => 
                           N3266);
   mult_21_C243_U153 : ADFULD1 port map( A => mult_21_C243_n651, B => 
                           mult_21_C243_n1194, CI => mult_21_C243_n185, CO => 
                           mult_21_C243_n184, S => N3267);
   mult_21_C243_U152 : ADFULD1 port map( A => mult_21_C243_n649, B => 
                           mult_21_C243_n1193, CI => mult_21_C243_n184, CO => 
                           mult_21_C243_n183, S => N3268);
   mult_21_C243_U151 : ADFULD1 port map( A => mult_21_C243_n645, B => 
                           mult_21_C243_n648, CI => mult_21_C243_n183, CO => 
                           mult_21_C243_n182, S => N3269);
   mult_21_C243_U150 : ADFULD1 port map( A => mult_21_C243_n641, B => 
                           mult_21_C243_n644, CI => mult_21_C243_n182, CO => 
                           mult_21_C243_n181, S => N3270);
   mult_21_C243_U149 : ADFULD1 port map( A => mult_21_C243_n635, B => 
                           mult_21_C243_n640, CI => mult_21_C243_n181, CO => 
                           mult_21_C243_n180, S => N3271);
   mult_21_C243_U148 : ADFULD1 port map( A => mult_21_C243_n629, B => 
                           mult_21_C243_n634, CI => mult_21_C243_n180, CO => 
                           mult_21_C243_n179, S => N3272);
   mult_21_C243_U147 : ADFULD1 port map( A => mult_21_C243_n621, B => 
                           mult_21_C243_n628, CI => mult_21_C243_n179, CO => 
                           mult_21_C243_n178, S => N3273);
   mult_21_C243_U146 : ADFULD1 port map( A => mult_21_C243_n613, B => 
                           mult_21_C243_n620, CI => mult_21_C243_n178, CO => 
                           mult_21_C243_n177, S => N3274);
   mult_21_C243_U145 : ADFULD1 port map( A => mult_21_C243_n603, B => 
                           mult_21_C243_n612, CI => mult_21_C243_n177, CO => 
                           mult_21_C243_n176, S => N3275);
   mult_21_C243_U144 : ADFULD1 port map( A => mult_21_C243_n593, B => 
                           mult_21_C243_n602, CI => mult_21_C243_n176, CO => 
                           mult_21_C243_n175, S => N3276);
   mult_21_C243_U143 : ADFULD1 port map( A => mult_21_C243_n581, B => 
                           mult_21_C243_n592, CI => mult_21_C243_n175, CO => 
                           mult_21_C243_n174, S => N3277);
   mult_21_C243_U142 : ADFULD1 port map( A => mult_21_C243_n569, B => 
                           mult_21_C243_n580, CI => mult_21_C243_n174, CO => 
                           mult_21_C243_n173, S => N3278);
   mult_21_C243_U141 : ADFULD1 port map( A => mult_21_C243_n555, B => 
                           mult_21_C243_n568, CI => mult_21_C243_n173, CO => 
                           mult_21_C243_n172, S => N3279);
   mult_21_C243_U140 : ADFULD1 port map( A => mult_21_C243_n541, B => 
                           mult_21_C243_n554, CI => mult_21_C243_n172, CO => 
                           mult_21_C243_n171, S => N3280);
   mult_21_C243_U139 : ADFULD1 port map( A => mult_21_C243_n525, B => 
                           mult_21_C243_n540, CI => mult_21_C243_n171, CO => 
                           mult_21_C243_n170, S => N3281);
   mult_21_C243_U138 : ADFULD1 port map( A => mult_21_C243_n509, B => 
                           mult_21_C243_n524, CI => mult_21_C243_n170, CO => 
                           mult_21_C243_n169, S => N3282);
   mult_21_C243_U137 : ADFULD1 port map( A => mult_21_C243_n491, B => 
                           mult_21_C243_n508, CI => mult_21_C243_n169, CO => 
                           mult_21_C243_n168, S => N3283);
   mult_21_C243_U136 : ADFULD1 port map( A => mult_21_C243_n473, B => 
                           mult_21_C243_n490, CI => mult_21_C243_n168, CO => 
                           mult_21_C243_n167, S => N3284);
   mult_21_C243_U135 : ADFULD1 port map( A => mult_21_C243_n453, B => 
                           mult_21_C243_n472, CI => mult_21_C243_n167, CO => 
                           mult_21_C243_n166, S => N3285);
   mult_21_C243_U134 : ADFULD1 port map( A => mult_21_C243_n433, B => 
                           mult_21_C243_n452, CI => mult_21_C243_n166, CO => 
                           mult_21_C243_n165, S => N3286);
   mult_21_C243_U133 : ADFULD1 port map( A => mult_21_C243_n411, B => 
                           mult_21_C243_n432, CI => mult_21_C243_n165, CO => 
                           mult_21_C243_n164, S => N3287);
   mult_21_C243_U132 : ADFULD1 port map( A => mult_21_C243_n389, B => 
                           mult_21_C243_n410, CI => mult_21_C243_n164, CO => 
                           mult_21_C243_n163, S => N3288);
   mult_21_C243_U131 : ADFULD1 port map( A => mult_21_C243_n365, B => 
                           mult_21_C243_n388, CI => mult_21_C243_n163, CO => 
                           mult_21_C243_n162, S => N3289);
   mult_21_C243_U130 : ADFULD1 port map( A => mult_21_C243_n341, B => 
                           mult_21_C243_n364, CI => mult_21_C243_n162, CO => 
                           mult_21_C243_n161, S => N3290);
   mult_21_C243_U129 : ADFULD1 port map( A => mult_21_C243_n315, B => 
                           mult_21_C243_n340, CI => mult_21_C243_n161, CO => 
                           mult_21_C243_n160, S => N3291);
   mult_21_C243_U128 : ADFULD1 port map( A => mult_21_C243_n289, B => 
                           mult_21_C243_n314, CI => mult_21_C243_n160, CO => 
                           mult_21_C243_n159, S => N3292);
   mult_21_C243_U127 : ADFULD1 port map( A => mult_21_C243_n261, B => 
                           mult_21_C243_n288, CI => mult_21_C243_n159, CO => 
                           mult_21_C243_n158, S => N3293);
   mult_21_C243_U126 : ADFULD1 port map( A => mult_21_C243_n233, B => 
                           mult_21_C243_n260, CI => mult_21_C243_n158, CO => 
                           mult_21_C243_n157, S => N3294);
   mult_21_C243_U125 : ADFULD1 port map( A => mult_21_C243_n203, B => 
                           mult_21_C243_n232, CI => mult_21_C243_n157, CO => 
                           mult_21_C243_n156, S => N3295);
   mult_21_C245_U1393 : AOI21D1 port map( A1 => N3004, A2 => N3005, B => 
                           mult_21_C245_n1418, Z => mult_21_C245_n940);
   mult_21_C245_U1392 : OAI21D1 port map( A1 => N3007, A2 => N3006, B => 
                           mult_21_C245_n1419, Z => mult_21_C245_n104);
   mult_21_C245_U1391 : AOI21D1 port map( A1 => N3006, A2 => N3007, B => 
                           mult_21_C245_n1419, Z => mult_21_C245_n939);
   mult_21_C245_U1390 : AOI21D1 port map( A1 => N2978, A2 => N2979, B => 
                           mult_21_C245_n1392, Z => mult_21_C245_n953);
   mult_21_C245_U1389 : AOI21D1 port map( A1 => N2980, A2 => N2981, B => 
                           mult_21_C245_n1394, Z => mult_21_C245_n952);
   mult_21_C245_U1388 : AOI21D1 port map( A1 => N2982, A2 => N2983, B => 
                           mult_21_C245_n1396, Z => mult_21_C245_n951);
   mult_21_C245_U1387 : AOI21D1 port map( A1 => N2984, A2 => N2985, B => 
                           mult_21_C245_n1398, Z => mult_21_C245_n950);
   mult_21_C245_U1386 : AOI21D1 port map( A1 => N2986, A2 => N2987, B => 
                           mult_21_C245_n1400, Z => mult_21_C245_n949);
   mult_21_C245_U1385 : AOI21D1 port map( A1 => N2988, A2 => N2989, B => 
                           mult_21_C245_n1402, Z => mult_21_C245_n948);
   mult_21_C245_U1384 : AOI21D1 port map( A1 => N2990, A2 => N2991, B => 
                           mult_21_C245_n1404, Z => mult_21_C245_n947);
   mult_21_C245_U1383 : EXOR2D1 port map( A1 => N3007, A2 => N3006, Z => 
                           mult_21_C245_n1448);
   mult_21_C245_U1382 : MUXB2DL port map( A0 => N3137, A1 => N3138, SL => 
                           mult_21_C245_n1448, Z => mult_21_C245_n652);
   mult_21_C245_U1381 : NAN2D1 port map( A1 => N3137, A2 => mult_21_C245_n1448,
                           Z => mult_21_C245_n653);
   mult_21_C245_U1380 : EXOR2D1 port map( A1 => N3005, A2 => N3004, Z => 
                           mult_21_C245_n1447);
   mult_21_C245_U1379 : MUXB2DL port map( A0 => N3139, A1 => N3140, SL => 
                           mult_21_C245_n1447, Z => mult_21_C245_n654);
   mult_21_C245_U1378 : MUXB2DL port map( A0 => mult_21_C245_n1387, A1 => N3139
                           , SL => mult_21_C245_n1447, Z => mult_21_C245_n655);
   mult_21_C245_U1377 : MUXB2DL port map( A0 => N3137, A1 => N3138, SL => 
                           mult_21_C245_n1447, Z => mult_21_C245_n656);
   mult_21_C245_U1376 : NAN2D1 port map( A1 => N3137, A2 => mult_21_C245_n1447,
                           Z => mult_21_C245_n657);
   mult_21_C245_U1375 : EXOR2D1 port map( A1 => N3003, A2 => N3002, Z => 
                           mult_21_C245_n1446);
   mult_21_C245_U1374 : MUXB2DL port map( A0 => N3141, A1 => N3142, SL => 
                           mult_21_C245_n1446, Z => mult_21_C245_n658);
   mult_21_C245_U1373 : MUXB2DL port map( A0 => mult_21_C245_n1385, A1 => N3141
                           , SL => mult_21_C245_n1446, Z => mult_21_C245_n659);
   mult_21_C245_U1372 : MUXB2DL port map( A0 => N3139, A1 => N3140, SL => 
                           mult_21_C245_n1446, Z => mult_21_C245_n660);
   mult_21_C245_U1371 : MUXB2DL port map( A0 => mult_21_C245_n1387, A1 => N3139
                           , SL => mult_21_C245_n1446, Z => mult_21_C245_n661);
   mult_21_C245_U1370 : MUXB2DL port map( A0 => N3137, A1 => N3138, SL => 
                           mult_21_C245_n1446, Z => mult_21_C245_n662);
   mult_21_C245_U1369 : NAN2D1 port map( A1 => N3137, A2 => mult_21_C245_n1446,
                           Z => mult_21_C245_n663);
   mult_21_C245_U1368 : EXOR2D1 port map( A1 => N3001, A2 => N3000, Z => 
                           mult_21_C245_n1445);
   mult_21_C245_U1367 : MUXB2DL port map( A0 => N3143, A1 => N3144, SL => 
                           mult_21_C245_n1445, Z => mult_21_C245_n664);
   mult_21_C245_U1366 : MUXB2DL port map( A0 => N3142, A1 => N3143, SL => 
                           mult_21_C245_n1445, Z => mult_21_C245_n665);
   mult_21_C245_U1365 : MUXB2DL port map( A0 => N3141, A1 => N3142, SL => 
                           mult_21_C245_n1445, Z => mult_21_C245_n666);
   mult_21_C245_U1364 : MUXB2DL port map( A0 => mult_21_C245_n1385, A1 => N3141
                           , SL => mult_21_C245_n1445, Z => mult_21_C245_n667);
   mult_21_C245_U1363 : MUXB2DL port map( A0 => N3139, A1 => N3140, SL => 
                           mult_21_C245_n1445, Z => mult_21_C245_n668);
   mult_21_C245_U1362 : MUXB2DL port map( A0 => mult_21_C245_n1387, A1 => N3139
                           , SL => mult_21_C245_n1445, Z => mult_21_C245_n669);
   mult_21_C245_U1361 : MUXB2DL port map( A0 => N3137, A1 => N3138, SL => 
                           mult_21_C245_n1445, Z => mult_21_C245_n670);
   mult_21_C245_U1360 : NAN2D1 port map( A1 => N3137, A2 => mult_21_C245_n1445,
                           Z => mult_21_C245_n671);
   mult_21_C245_U1359 : MUXB2DL port map( A0 => N3145, A1 => N3146, SL => 
                           mult_21_C245_n1444, Z => mult_21_C245_n672);
   mult_21_C245_U1358 : MUXB2DL port map( A0 => N3144, A1 => N3145, SL => 
                           mult_21_C245_n1444, Z => mult_21_C245_n673);
   mult_21_C245_U1357 : MUXB2DL port map( A0 => N3143, A1 => N3144, SL => 
                           mult_21_C245_n1444, Z => mult_21_C245_n674);
   mult_21_C245_U1356 : MUXB2DL port map( A0 => N3142, A1 => N3143, SL => 
                           mult_21_C245_n1444, Z => mult_21_C245_n675);
   mult_21_C245_U1355 : MUXB2DL port map( A0 => N3141, A1 => N3142, SL => 
                           mult_21_C245_n1444, Z => mult_21_C245_n676);
   mult_21_C245_U1354 : MUXB2DL port map( A0 => mult_21_C245_n1385, A1 => N3141
                           , SL => mult_21_C245_n1444, Z => mult_21_C245_n677);
   mult_21_C245_U1353 : MUXB2DL port map( A0 => N3139, A1 => N3140, SL => 
                           mult_21_C245_n1444, Z => mult_21_C245_n678);
   mult_21_C245_U1352 : MUXB2DL port map( A0 => mult_21_C245_n1387, A1 => N3139
                           , SL => mult_21_C245_n1444, Z => mult_21_C245_n679);
   mult_21_C245_U1351 : AOI21D1 port map( A1 => N2992, A2 => N2993, B => 
                           mult_21_C245_n1406, Z => mult_21_C245_n946);
   mult_21_C245_U1350 : MUXB2DL port map( A0 => N3137, A1 => N3138, SL => 
                           mult_21_C245_n1444, Z => mult_21_C245_n680);
   mult_21_C245_U1349 : NAN2D1 port map( A1 => N3137, A2 => mult_21_C245_n1444,
                           Z => mult_21_C245_n681);
   mult_21_C245_U1348 : MUXB2DL port map( A0 => N3147, A1 => N3148, SL => 
                           mult_21_C245_n1443, Z => mult_21_C245_n682);
   mult_21_C245_U1347 : MUXB2DL port map( A0 => N3146, A1 => N3147, SL => 
                           mult_21_C245_n1443, Z => mult_21_C245_n683);
   mult_21_C245_U1346 : MUXB2DL port map( A0 => N3145, A1 => N3146, SL => 
                           mult_21_C245_n1443, Z => mult_21_C245_n684);
   mult_21_C245_U1345 : MUXB2DL port map( A0 => N3144, A1 => N3145, SL => 
                           mult_21_C245_n1443, Z => mult_21_C245_n685);
   mult_21_C245_U1344 : MUXB2DL port map( A0 => N3143, A1 => N3144, SL => 
                           mult_21_C245_n1443, Z => mult_21_C245_n686);
   mult_21_C245_U1343 : MUXB2DL port map( A0 => N3142, A1 => N3143, SL => 
                           mult_21_C245_n1443, Z => mult_21_C245_n687);
   mult_21_C245_U1342 : MUXB2DL port map( A0 => N3141, A1 => N3142, SL => 
                           mult_21_C245_n1443, Z => mult_21_C245_n688);
   mult_21_C245_U1341 : MUXB2DL port map( A0 => mult_21_C245_n1385, A1 => N3141
                           , SL => mult_21_C245_n1443, Z => mult_21_C245_n689);
   mult_21_C245_U1340 : MUXB2DL port map( A0 => N3139, A1 => N3140, SL => 
                           mult_21_C245_n1443, Z => mult_21_C245_n690);
   mult_21_C245_U1339 : MUXB2DL port map( A0 => mult_21_C245_n1387, A1 => N3139
                           , SL => mult_21_C245_n1443, Z => mult_21_C245_n691);
   mult_21_C245_U1338 : MUXB2DL port map( A0 => N3137, A1 => N3138, SL => 
                           mult_21_C245_n1443, Z => mult_21_C245_n692);
   mult_21_C245_U1337 : NAN2D1 port map( A1 => N3137, A2 => mult_21_C245_n1443,
                           Z => mult_21_C245_n693);
   mult_21_C245_U1336 : MUXB2DL port map( A0 => N3149, A1 => N3150, SL => 
                           mult_21_C245_n1442, Z => mult_21_C245_n694);
   mult_21_C245_U1335 : MUXB2DL port map( A0 => N3148, A1 => N3149, SL => 
                           mult_21_C245_n1442, Z => mult_21_C245_n695);
   mult_21_C245_U1334 : MUXB2DL port map( A0 => N3147, A1 => N3148, SL => 
                           mult_21_C245_n1442, Z => mult_21_C245_n696);
   mult_21_C245_U1333 : MUXB2DL port map( A0 => N3146, A1 => N3147, SL => 
                           mult_21_C245_n1442, Z => mult_21_C245_n697);
   mult_21_C245_U1332 : MUXB2DL port map( A0 => N3145, A1 => N3146, SL => 
                           mult_21_C245_n1442, Z => mult_21_C245_n698);
   mult_21_C245_U1331 : MUXB2DL port map( A0 => N3144, A1 => N3145, SL => 
                           mult_21_C245_n1442, Z => mult_21_C245_n699);
   mult_21_C245_U1330 : MUXB2DL port map( A0 => N3143, A1 => N3144, SL => 
                           mult_21_C245_n1442, Z => mult_21_C245_n700);
   mult_21_C245_U1329 : MUXB2DL port map( A0 => N3142, A1 => N3143, SL => 
                           mult_21_C245_n1442, Z => mult_21_C245_n701);
   mult_21_C245_U1328 : MUXB2DL port map( A0 => N3141, A1 => N3142, SL => 
                           mult_21_C245_n1442, Z => mult_21_C245_n702);
   mult_21_C245_U1327 : MUXB2DL port map( A0 => mult_21_C245_n1385, A1 => N3141
                           , SL => mult_21_C245_n1442, Z => mult_21_C245_n703);
   mult_21_C245_U1326 : MUXB2DL port map( A0 => N3139, A1 => N3140, SL => 
                           mult_21_C245_n1442, Z => mult_21_C245_n704);
   mult_21_C245_U1325 : MUXB2DL port map( A0 => mult_21_C245_n1387, A1 => N3139
                           , SL => mult_21_C245_n1442, Z => mult_21_C245_n705);
   mult_21_C245_U1324 : MUXB2DL port map( A0 => N3137, A1 => N3138, SL => 
                           mult_21_C245_n1442, Z => mult_21_C245_n706);
   mult_21_C245_U1323 : NAN2D1 port map( A1 => N3137, A2 => mult_21_C245_n1442,
                           Z => mult_21_C245_n707);
   mult_21_C245_U1322 : MUXB2DL port map( A0 => N3151, A1 => N3152, SL => 
                           mult_21_C245_n1441, Z => mult_21_C245_n708);
   mult_21_C245_U1321 : MUXB2DL port map( A0 => N3150, A1 => N3151, SL => 
                           mult_21_C245_n1441, Z => mult_21_C245_n709);
   mult_21_C245_U1320 : MUXB2DL port map( A0 => N3149, A1 => N3150, SL => 
                           mult_21_C245_n1441, Z => mult_21_C245_n710);
   mult_21_C245_U1319 : MUXB2DL port map( A0 => N3148, A1 => N3149, SL => 
                           mult_21_C245_n1441, Z => mult_21_C245_n711);
   mult_21_C245_U1318 : MUXB2DL port map( A0 => N3147, A1 => N3148, SL => 
                           mult_21_C245_n1441, Z => mult_21_C245_n712);
   mult_21_C245_U1317 : MUXB2DL port map( A0 => N3146, A1 => N3147, SL => 
                           mult_21_C245_n1441, Z => mult_21_C245_n713);
   mult_21_C245_U1316 : MUXB2DL port map( A0 => N3145, A1 => N3146, SL => 
                           mult_21_C245_n1441, Z => mult_21_C245_n714);
   mult_21_C245_U1315 : MUXB2DL port map( A0 => N3144, A1 => N3145, SL => 
                           mult_21_C245_n1441, Z => mult_21_C245_n715);
   mult_21_C245_U1314 : MUXB2DL port map( A0 => N3143, A1 => N3144, SL => 
                           mult_21_C245_n1441, Z => mult_21_C245_n716);
   mult_21_C245_U1313 : MUXB2DL port map( A0 => N3142, A1 => N3143, SL => 
                           mult_21_C245_n1441, Z => mult_21_C245_n717);
   mult_21_C245_U1312 : MUXB2DL port map( A0 => N3141, A1 => N3142, SL => 
                           mult_21_C245_n1441, Z => mult_21_C245_n718);
   mult_21_C245_U1311 : MUXB2DL port map( A0 => mult_21_C245_n1385, A1 => N3141
                           , SL => mult_21_C245_n1441, Z => mult_21_C245_n719);
   mult_21_C245_U1310 : MUXB2DL port map( A0 => N3139, A1 => N3140, SL => 
                           mult_21_C245_n1441, Z => mult_21_C245_n720);
   mult_21_C245_U1309 : MUXB2DL port map( A0 => mult_21_C245_n1387, A1 => N3139
                           , SL => mult_21_C245_n1441, Z => mult_21_C245_n721);
   mult_21_C245_U1308 : MUXB2DL port map( A0 => N3137, A1 => N3138, SL => 
                           mult_21_C245_n1441, Z => mult_21_C245_n722);
   mult_21_C245_U1307 : NAN2D1 port map( A1 => N3137, A2 => mult_21_C245_n1441,
                           Z => mult_21_C245_n723);
   mult_21_C245_U1306 : MUXB2DL port map( A0 => N3153, A1 => N3154, SL => 
                           mult_21_C245_n1440, Z => mult_21_C245_n724);
   mult_21_C245_U1305 : MUXB2DL port map( A0 => N3152, A1 => N3153, SL => 
                           mult_21_C245_n1440, Z => mult_21_C245_n725);
   mult_21_C245_U1304 : MUXB2DL port map( A0 => N3151, A1 => N3152, SL => 
                           mult_21_C245_n1440, Z => mult_21_C245_n726);
   mult_21_C245_U1303 : MUXB2DL port map( A0 => N3150, A1 => N3151, SL => 
                           mult_21_C245_n1440, Z => mult_21_C245_n727);
   mult_21_C245_U1302 : MUXB2DL port map( A0 => N3149, A1 => N3150, SL => 
                           mult_21_C245_n1440, Z => mult_21_C245_n728);
   mult_21_C245_U1301 : MUXB2DL port map( A0 => N3148, A1 => N3149, SL => 
                           mult_21_C245_n1440, Z => mult_21_C245_n729);
   mult_21_C245_U1300 : MUXB2DL port map( A0 => N3147, A1 => N3148, SL => 
                           mult_21_C245_n1440, Z => mult_21_C245_n730);
   mult_21_C245_U1299 : MUXB2DL port map( A0 => N3146, A1 => N3147, SL => 
                           mult_21_C245_n1440, Z => mult_21_C245_n731);
   mult_21_C245_U1298 : MUXB2DL port map( A0 => N3145, A1 => N3146, SL => 
                           mult_21_C245_n1440, Z => mult_21_C245_n732);
   mult_21_C245_U1297 : MUXB2DL port map( A0 => N3144, A1 => N3145, SL => 
                           mult_21_C245_n1440, Z => mult_21_C245_n733);
   mult_21_C245_U1296 : MUXB2DL port map( A0 => N3143, A1 => N3144, SL => 
                           mult_21_C245_n1440, Z => mult_21_C245_n734);
   mult_21_C245_U1295 : MUXB2DL port map( A0 => N3142, A1 => N3143, SL => 
                           mult_21_C245_n1440, Z => mult_21_C245_n735);
   mult_21_C245_U1294 : MUXB2DL port map( A0 => N3141, A1 => N3142, SL => 
                           mult_21_C245_n1440, Z => mult_21_C245_n736);
   mult_21_C245_U1293 : MUXB2DL port map( A0 => mult_21_C245_n1385, A1 => N3141
                           , SL => mult_21_C245_n1440, Z => mult_21_C245_n737);
   mult_21_C245_U1292 : MUXB2DL port map( A0 => N3139, A1 => N3140, SL => 
                           mult_21_C245_n1440, Z => mult_21_C245_n738);
   mult_21_C245_U1291 : MUXB2DL port map( A0 => mult_21_C245_n1387, A1 => N3139
                           , SL => mult_21_C245_n1440, Z => mult_21_C245_n739);
   mult_21_C245_U1290 : MUXB2DL port map( A0 => N3137, A1 => N3138, SL => 
                           mult_21_C245_n1440, Z => mult_21_C245_n740);
   mult_21_C245_U1289 : NAN2D1 port map( A1 => N3137, A2 => mult_21_C245_n1440,
                           Z => mult_21_C245_n741);
   mult_21_C245_U1288 : MUXB2DL port map( A0 => N3155, A1 => N3156, SL => 
                           mult_21_C245_n1439, Z => mult_21_C245_n742);
   mult_21_C245_U1287 : MUXB2DL port map( A0 => N3154, A1 => N3155, SL => 
                           mult_21_C245_n1439, Z => mult_21_C245_n743);
   mult_21_C245_U1286 : MUXB2DL port map( A0 => N3153, A1 => N3154, SL => 
                           mult_21_C245_n1439, Z => mult_21_C245_n744);
   mult_21_C245_U1285 : MUXB2DL port map( A0 => N3152, A1 => N3153, SL => 
                           mult_21_C245_n1439, Z => mult_21_C245_n745);
   mult_21_C245_U1284 : MUXB2DL port map( A0 => N3151, A1 => N3152, SL => 
                           mult_21_C245_n1439, Z => mult_21_C245_n746);
   mult_21_C245_U1283 : MUXB2DL port map( A0 => N3150, A1 => N3151, SL => 
                           mult_21_C245_n1439, Z => mult_21_C245_n747);
   mult_21_C245_U1282 : MUXB2DL port map( A0 => N3149, A1 => N3150, SL => 
                           mult_21_C245_n1439, Z => mult_21_C245_n748);
   mult_21_C245_U1281 : MUXB2DL port map( A0 => N3148, A1 => N3149, SL => 
                           mult_21_C245_n1439, Z => mult_21_C245_n749);
   mult_21_C245_U1280 : AOI21D1 port map( A1 => N2994, A2 => N2995, B => 
                           mult_21_C245_n1408, Z => mult_21_C245_n945);
   mult_21_C245_U1279 : MUXB2DL port map( A0 => N3147, A1 => N3148, SL => 
                           mult_21_C245_n1439, Z => mult_21_C245_n750);
   mult_21_C245_U1278 : MUXB2DL port map( A0 => N3146, A1 => N3147, SL => 
                           mult_21_C245_n1439, Z => mult_21_C245_n751);
   mult_21_C245_U1277 : MUXB2DL port map( A0 => N3145, A1 => N3146, SL => 
                           mult_21_C245_n1439, Z => mult_21_C245_n752);
   mult_21_C245_U1276 : MUXB2DL port map( A0 => N3144, A1 => N3145, SL => 
                           mult_21_C245_n1439, Z => mult_21_C245_n753);
   mult_21_C245_U1275 : MUXB2DL port map( A0 => N3143, A1 => N3144, SL => 
                           mult_21_C245_n1439, Z => mult_21_C245_n754);
   mult_21_C245_U1274 : MUXB2DL port map( A0 => N3142, A1 => N3143, SL => 
                           mult_21_C245_n1439, Z => mult_21_C245_n755);
   mult_21_C245_U1273 : MUXB2DL port map( A0 => N3141, A1 => N3142, SL => 
                           mult_21_C245_n1439, Z => mult_21_C245_n756);
   mult_21_C245_U1272 : MUXB2DL port map( A0 => mult_21_C245_n1385, A1 => N3141
                           , SL => mult_21_C245_n1439, Z => mult_21_C245_n757);
   mult_21_C245_U1271 : MUXB2DL port map( A0 => N3139, A1 => N3140, SL => 
                           mult_21_C245_n1439, Z => mult_21_C245_n758);
   mult_21_C245_U1270 : MUXB2DL port map( A0 => N3138, A1 => N3139, SL => 
                           mult_21_C245_n1439, Z => mult_21_C245_n759);
   mult_21_C245_U1269 : MUXB2DL port map( A0 => N3137, A1 => N3138, SL => 
                           mult_21_C245_n1439, Z => mult_21_C245_n760);
   mult_21_C245_U1268 : NAN2D1 port map( A1 => N3137, A2 => mult_21_C245_n1439,
                           Z => mult_21_C245_n761);
   mult_21_C245_U1267 : MUXB2DL port map( A0 => N3157, A1 => N3158, SL => 
                           mult_21_C245_n1438, Z => mult_21_C245_n762);
   mult_21_C245_U1266 : MUXB2DL port map( A0 => N3156, A1 => N3157, SL => 
                           mult_21_C245_n1438, Z => mult_21_C245_n763);
   mult_21_C245_U1265 : MUXB2DL port map( A0 => N3155, A1 => N3156, SL => 
                           mult_21_C245_n1438, Z => mult_21_C245_n764);
   mult_21_C245_U1264 : MUXB2DL port map( A0 => N3154, A1 => N3155, SL => 
                           mult_21_C245_n1438, Z => mult_21_C245_n765);
   mult_21_C245_U1263 : MUXB2DL port map( A0 => N3153, A1 => N3154, SL => 
                           mult_21_C245_n1438, Z => mult_21_C245_n766);
   mult_21_C245_U1262 : MUXB2DL port map( A0 => N3152, A1 => N3153, SL => 
                           mult_21_C245_n1438, Z => mult_21_C245_n767);
   mult_21_C245_U1261 : MUXB2DL port map( A0 => N3151, A1 => N3152, SL => 
                           mult_21_C245_n1438, Z => mult_21_C245_n768);
   mult_21_C245_U1260 : MUXB2DL port map( A0 => N3150, A1 => N3151, SL => 
                           mult_21_C245_n1438, Z => mult_21_C245_n769);
   mult_21_C245_U1259 : MUXB2DL port map( A0 => N3149, A1 => N3150, SL => 
                           mult_21_C245_n1438, Z => mult_21_C245_n770);
   mult_21_C245_U1258 : MUXB2DL port map( A0 => N3148, A1 => N3149, SL => 
                           mult_21_C245_n1438, Z => mult_21_C245_n771);
   mult_21_C245_U1257 : MUXB2DL port map( A0 => N3147, A1 => N3148, SL => 
                           mult_21_C245_n1438, Z => mult_21_C245_n772);
   mult_21_C245_U1256 : MUXB2DL port map( A0 => N3146, A1 => N3147, SL => 
                           mult_21_C245_n1438, Z => mult_21_C245_n773);
   mult_21_C245_U1255 : MUXB2DL port map( A0 => N3145, A1 => N3146, SL => 
                           mult_21_C245_n1438, Z => mult_21_C245_n774);
   mult_21_C245_U1254 : MUXB2DL port map( A0 => N3144, A1 => N3145, SL => 
                           mult_21_C245_n1438, Z => mult_21_C245_n775);
   mult_21_C245_U1253 : MUXB2DL port map( A0 => N3143, A1 => N3144, SL => 
                           mult_21_C245_n1438, Z => mult_21_C245_n776);
   mult_21_C245_U1252 : MUXB2DL port map( A0 => N3142, A1 => N3143, SL => 
                           mult_21_C245_n1438, Z => mult_21_C245_n777);
   mult_21_C245_U1251 : MUXB2DL port map( A0 => N3141, A1 => N3142, SL => 
                           mult_21_C245_n1438, Z => mult_21_C245_n778);
   mult_21_C245_U1250 : MUXB2DL port map( A0 => N3140, A1 => N3141, SL => 
                           mult_21_C245_n1438, Z => mult_21_C245_n779);
   mult_21_C245_U1249 : MUXB2DL port map( A0 => N3139, A1 => N3140, SL => 
                           mult_21_C245_n1438, Z => mult_21_C245_n780);
   mult_21_C245_U1248 : MUXB2DL port map( A0 => mult_21_C245_n1387, A1 => N3139
                           , SL => mult_21_C245_n1438, Z => mult_21_C245_n781);
   mult_21_C245_U1247 : MUXB2DL port map( A0 => N3137, A1 => N3138, SL => 
                           mult_21_C245_n1438, Z => mult_21_C245_n782);
   mult_21_C245_U1246 : NAN2D1 port map( A1 => N3137, A2 => mult_21_C245_n1438,
                           Z => mult_21_C245_n783);
   mult_21_C245_U1245 : MUXB2DL port map( A0 => N3159, A1 => N3160, SL => 
                           mult_21_C245_n1377, Z => mult_21_C245_n784);
   mult_21_C245_U1244 : MUXB2DL port map( A0 => N3158, A1 => N3159, SL => 
                           mult_21_C245_n1377, Z => mult_21_C245_n785);
   mult_21_C245_U1243 : MUXB2DL port map( A0 => N3157, A1 => N3158, SL => 
                           mult_21_C245_n1377, Z => mult_21_C245_n786);
   mult_21_C245_U1242 : MUXB2DL port map( A0 => N3156, A1 => N3157, SL => 
                           mult_21_C245_n1377, Z => mult_21_C245_n787);
   mult_21_C245_U1241 : MUXB2DL port map( A0 => N3155, A1 => N3156, SL => 
                           mult_21_C245_n1377, Z => mult_21_C245_n788);
   mult_21_C245_U1240 : MUXB2DL port map( A0 => N3154, A1 => N3155, SL => 
                           mult_21_C245_n1377, Z => mult_21_C245_n789);
   mult_21_C245_U1239 : MUXB2DL port map( A0 => N3153, A1 => N3154, SL => 
                           mult_21_C245_n1377, Z => mult_21_C245_n790);
   mult_21_C245_U1238 : MUXB2DL port map( A0 => N3152, A1 => N3153, SL => 
                           mult_21_C245_n1377, Z => mult_21_C245_n791);
   mult_21_C245_U1237 : MUXB2DL port map( A0 => N3151, A1 => N3152, SL => 
                           mult_21_C245_n1377, Z => mult_21_C245_n792);
   mult_21_C245_U1236 : MUXB2DL port map( A0 => N3150, A1 => N3151, SL => 
                           mult_21_C245_n1377, Z => mult_21_C245_n793);
   mult_21_C245_U1235 : MUXB2DL port map( A0 => N3149, A1 => N3150, SL => 
                           mult_21_C245_n1377, Z => mult_21_C245_n794);
   mult_21_C245_U1234 : MUXB2DL port map( A0 => N3148, A1 => N3149, SL => 
                           mult_21_C245_n1377, Z => mult_21_C245_n795);
   mult_21_C245_U1233 : MUXB2DL port map( A0 => N3147, A1 => N3148, SL => 
                           mult_21_C245_n1377, Z => mult_21_C245_n796);
   mult_21_C245_U1232 : MUXB2DL port map( A0 => N3146, A1 => N3147, SL => 
                           mult_21_C245_n1377, Z => mult_21_C245_n797);
   mult_21_C245_U1231 : MUXB2DL port map( A0 => N3145, A1 => N3146, SL => 
                           mult_21_C245_n1377, Z => mult_21_C245_n798);
   mult_21_C245_U1230 : MUXB2DL port map( A0 => N3144, A1 => N3145, SL => 
                           mult_21_C245_n1377, Z => mult_21_C245_n799);
   mult_21_C245_U1229 : MUXB2DL port map( A0 => N3143, A1 => N3144, SL => 
                           mult_21_C245_n1377, Z => mult_21_C245_n800);
   mult_21_C245_U1228 : MUXB2DL port map( A0 => N3142, A1 => N3143, SL => 
                           mult_21_C245_n1377, Z => mult_21_C245_n801);
   mult_21_C245_U1227 : MUXB2DL port map( A0 => N3141, A1 => N3142, SL => 
                           mult_21_C245_n1377, Z => mult_21_C245_n802);
   mult_21_C245_U1226 : MUXB2DL port map( A0 => mult_21_C245_n1385, A1 => N3141
                           , SL => mult_21_C245_n1377, Z => mult_21_C245_n803);
   mult_21_C245_U1225 : MUXB2DL port map( A0 => N3139, A1 => N3140, SL => 
                           mult_21_C245_n1377, Z => mult_21_C245_n804);
   mult_21_C245_U1224 : MUXB2DL port map( A0 => N3138, A1 => N3139, SL => 
                           mult_21_C245_n1377, Z => mult_21_C245_n805);
   mult_21_C245_U1223 : MUXB2DL port map( A0 => N3137, A1 => N3138, SL => 
                           mult_21_C245_n1377, Z => mult_21_C245_n806);
   mult_21_C245_U1222 : NAN2D1 port map( A1 => N3137, A2 => mult_21_C245_n1377,
                           Z => mult_21_C245_n807);
   mult_21_C245_U1221 : MUXB2DL port map( A0 => N3161, A1 => N3162, SL => 
                           mult_21_C245_n1376, Z => mult_21_C245_n808);
   mult_21_C245_U1220 : MUXB2DL port map( A0 => N3160, A1 => N3161, SL => 
                           mult_21_C245_n1376, Z => mult_21_C245_n809);
   mult_21_C245_U1219 : AOI21D1 port map( A1 => N2996, A2 => N2997, B => 
                           mult_21_C245_n1410, Z => mult_21_C245_n944);
   mult_21_C245_U1218 : MUXB2DL port map( A0 => N3159, A1 => N3160, SL => 
                           mult_21_C245_n1376, Z => mult_21_C245_n810);
   mult_21_C245_U1217 : MUXB2DL port map( A0 => N3158, A1 => N3159, SL => 
                           mult_21_C245_n1376, Z => mult_21_C245_n811);
   mult_21_C245_U1216 : MUXB2DL port map( A0 => N3157, A1 => N3158, SL => 
                           mult_21_C245_n1376, Z => mult_21_C245_n812);
   mult_21_C245_U1215 : MUXB2DL port map( A0 => N3156, A1 => N3157, SL => 
                           mult_21_C245_n1376, Z => mult_21_C245_n813);
   mult_21_C245_U1214 : MUXB2DL port map( A0 => N3155, A1 => N3156, SL => 
                           mult_21_C245_n1376, Z => mult_21_C245_n814);
   mult_21_C245_U1213 : MUXB2DL port map( A0 => N3154, A1 => N3155, SL => 
                           mult_21_C245_n1376, Z => mult_21_C245_n815);
   mult_21_C245_U1212 : MUXB2DL port map( A0 => N3153, A1 => N3154, SL => 
                           mult_21_C245_n1376, Z => mult_21_C245_n816);
   mult_21_C245_U1211 : MUXB2DL port map( A0 => N3152, A1 => N3153, SL => 
                           mult_21_C245_n1376, Z => mult_21_C245_n817);
   mult_21_C245_U1210 : MUXB2DL port map( A0 => N3151, A1 => N3152, SL => 
                           mult_21_C245_n1376, Z => mult_21_C245_n818);
   mult_21_C245_U1209 : MUXB2DL port map( A0 => N3150, A1 => N3151, SL => 
                           mult_21_C245_n1376, Z => mult_21_C245_n819);
   mult_21_C245_U1208 : MUXB2DL port map( A0 => N3149, A1 => N3150, SL => 
                           mult_21_C245_n1376, Z => mult_21_C245_n820);
   mult_21_C245_U1207 : MUXB2DL port map( A0 => N3148, A1 => N3149, SL => 
                           mult_21_C245_n1376, Z => mult_21_C245_n821);
   mult_21_C245_U1206 : MUXB2DL port map( A0 => N3147, A1 => N3148, SL => 
                           mult_21_C245_n1376, Z => mult_21_C245_n822);
   mult_21_C245_U1205 : MUXB2DL port map( A0 => N3146, A1 => N3147, SL => 
                           mult_21_C245_n1376, Z => mult_21_C245_n823);
   mult_21_C245_U1204 : MUXB2DL port map( A0 => N3145, A1 => N3146, SL => 
                           mult_21_C245_n1376, Z => mult_21_C245_n824);
   mult_21_C245_U1203 : MUXB2DL port map( A0 => N3144, A1 => N3145, SL => 
                           mult_21_C245_n1376, Z => mult_21_C245_n825);
   mult_21_C245_U1202 : MUXB2DL port map( A0 => N3143, A1 => N3144, SL => 
                           mult_21_C245_n1376, Z => mult_21_C245_n826);
   mult_21_C245_U1201 : MUXB2DL port map( A0 => N3142, A1 => N3143, SL => 
                           mult_21_C245_n1376, Z => mult_21_C245_n827);
   mult_21_C245_U1200 : MUXB2DL port map( A0 => N3141, A1 => N3142, SL => 
                           mult_21_C245_n1376, Z => mult_21_C245_n828);
   mult_21_C245_U1199 : MUXB2DL port map( A0 => mult_21_C245_n1385, A1 => N3141
                           , SL => mult_21_C245_n1376, Z => mult_21_C245_n829);
   mult_21_C245_U1198 : MUXB2DL port map( A0 => N3139, A1 => N3140, SL => 
                           mult_21_C245_n1376, Z => mult_21_C245_n830);
   mult_21_C245_U1197 : MUXB2DL port map( A0 => mult_21_C245_n1387, A1 => N3139
                           , SL => mult_21_C245_n1376, Z => mult_21_C245_n831);
   mult_21_C245_U1196 : MUXB2DL port map( A0 => N3137, A1 => N3138, SL => 
                           mult_21_C245_n1376, Z => mult_21_C245_n832);
   mult_21_C245_U1195 : NAN2D1 port map( A1 => N3137, A2 => mult_21_C245_n1376,
                           Z => mult_21_C245_n833);
   mult_21_C245_U1194 : MUXB2DL port map( A0 => N3163, A1 => N3164, SL => 
                           mult_21_C245_n1375, Z => mult_21_C245_n834);
   mult_21_C245_U1193 : MUXB2DL port map( A0 => N3162, A1 => N3163, SL => 
                           mult_21_C245_n1375, Z => mult_21_C245_n835);
   mult_21_C245_U1192 : MUXB2DL port map( A0 => N3161, A1 => N3162, SL => 
                           mult_21_C245_n1375, Z => mult_21_C245_n836);
   mult_21_C245_U1191 : MUXB2DL port map( A0 => N3160, A1 => N3161, SL => 
                           mult_21_C245_n1375, Z => mult_21_C245_n837);
   mult_21_C245_U1190 : MUXB2DL port map( A0 => N3159, A1 => N3160, SL => 
                           mult_21_C245_n1375, Z => mult_21_C245_n838);
   mult_21_C245_U1189 : MUXB2DL port map( A0 => N3158, A1 => N3159, SL => 
                           mult_21_C245_n1375, Z => mult_21_C245_n839);
   mult_21_C245_U1188 : MUXB2DL port map( A0 => N3157, A1 => N3158, SL => 
                           mult_21_C245_n1375, Z => mult_21_C245_n840);
   mult_21_C245_U1187 : MUXB2DL port map( A0 => N3156, A1 => N3157, SL => 
                           mult_21_C245_n1375, Z => mult_21_C245_n841);
   mult_21_C245_U1186 : MUXB2DL port map( A0 => N3155, A1 => N3156, SL => 
                           mult_21_C245_n1375, Z => mult_21_C245_n842);
   mult_21_C245_U1185 : MUXB2DL port map( A0 => N3154, A1 => N3155, SL => 
                           mult_21_C245_n1375, Z => mult_21_C245_n843);
   mult_21_C245_U1184 : MUXB2DL port map( A0 => N3153, A1 => N3154, SL => 
                           mult_21_C245_n1375, Z => mult_21_C245_n844);
   mult_21_C245_U1183 : MUXB2DL port map( A0 => N3152, A1 => N3153, SL => 
                           mult_21_C245_n1375, Z => mult_21_C245_n845);
   mult_21_C245_U1182 : MUXB2DL port map( A0 => N3151, A1 => N3152, SL => 
                           mult_21_C245_n1375, Z => mult_21_C245_n846);
   mult_21_C245_U1181 : MUXB2DL port map( A0 => N3150, A1 => N3151, SL => 
                           mult_21_C245_n1375, Z => mult_21_C245_n847);
   mult_21_C245_U1180 : MUXB2DL port map( A0 => N3149, A1 => N3150, SL => 
                           mult_21_C245_n1375, Z => mult_21_C245_n848);
   mult_21_C245_U1179 : MUXB2DL port map( A0 => N3148, A1 => N3149, SL => 
                           mult_21_C245_n1375, Z => mult_21_C245_n849);
   mult_21_C245_U1178 : MUXB2DL port map( A0 => N3147, A1 => N3148, SL => 
                           mult_21_C245_n1375, Z => mult_21_C245_n850);
   mult_21_C245_U1177 : MUXB2DL port map( A0 => N3146, A1 => N3147, SL => 
                           mult_21_C245_n1375, Z => mult_21_C245_n851);
   mult_21_C245_U1176 : MUXB2DL port map( A0 => N3145, A1 => N3146, SL => 
                           mult_21_C245_n1375, Z => mult_21_C245_n852);
   mult_21_C245_U1175 : MUXB2DL port map( A0 => N3144, A1 => N3145, SL => 
                           mult_21_C245_n1375, Z => mult_21_C245_n853);
   mult_21_C245_U1174 : MUXB2DL port map( A0 => N3143, A1 => N3144, SL => 
                           mult_21_C245_n1375, Z => mult_21_C245_n854);
   mult_21_C245_U1173 : MUXB2DL port map( A0 => N3142, A1 => N3143, SL => 
                           mult_21_C245_n1375, Z => mult_21_C245_n855);
   mult_21_C245_U1172 : MUXB2DL port map( A0 => N3141, A1 => N3142, SL => 
                           mult_21_C245_n1375, Z => mult_21_C245_n856);
   mult_21_C245_U1171 : MUXB2DL port map( A0 => mult_21_C245_n1385, A1 => N3141
                           , SL => mult_21_C245_n1375, Z => mult_21_C245_n857);
   mult_21_C245_U1170 : MUXB2DL port map( A0 => N3139, A1 => N3140, SL => 
                           mult_21_C245_n1375, Z => mult_21_C245_n858);
   mult_21_C245_U1169 : MUXB2DL port map( A0 => mult_21_C245_n1387, A1 => N3139
                           , SL => mult_21_C245_n1375, Z => mult_21_C245_n859);
   mult_21_C245_U1168 : AOI21D1 port map( A1 => N2998, A2 => N2999, B => 
                           mult_21_C245_n1412, Z => mult_21_C245_n943);
   mult_21_C245_U1167 : MUXB2DL port map( A0 => N3137, A1 => N3138, SL => 
                           mult_21_C245_n1375, Z => mult_21_C245_n860);
   mult_21_C245_U1166 : NAN2D1 port map( A1 => N3137, A2 => mult_21_C245_n1375,
                           Z => mult_21_C245_n861);
   mult_21_C245_U1165 : MUXB2DL port map( A0 => N3164, A1 => N3165, SL => 
                           mult_21_C245_n1384, Z => mult_21_C245_n863);
   mult_21_C245_U1164 : MUXB2DL port map( A0 => N3163, A1 => N3164, SL => 
                           mult_21_C245_n1384, Z => mult_21_C245_n864);
   mult_21_C245_U1163 : MUXB2DL port map( A0 => N3162, A1 => N3163, SL => 
                           mult_21_C245_n1384, Z => mult_21_C245_n865);
   mult_21_C245_U1162 : MUXB2DL port map( A0 => N3161, A1 => N3162, SL => 
                           mult_21_C245_n1384, Z => mult_21_C245_n866);
   mult_21_C245_U1161 : MUXB2DL port map( A0 => N3160, A1 => N3161, SL => 
                           mult_21_C245_n1384, Z => mult_21_C245_n867);
   mult_21_C245_U1160 : MUXB2DL port map( A0 => N3159, A1 => N3160, SL => 
                           mult_21_C245_n1384, Z => mult_21_C245_n868);
   mult_21_C245_U1159 : MUXB2DL port map( A0 => N3158, A1 => N3159, SL => 
                           mult_21_C245_n1384, Z => mult_21_C245_n869);
   mult_21_C245_U1158 : MUXB2DL port map( A0 => N3157, A1 => N3158, SL => 
                           mult_21_C245_n1384, Z => mult_21_C245_n870);
   mult_21_C245_U1157 : MUXB2DL port map( A0 => N3156, A1 => N3157, SL => 
                           mult_21_C245_n1384, Z => mult_21_C245_n871);
   mult_21_C245_U1156 : MUXB2DL port map( A0 => N3155, A1 => N3156, SL => 
                           mult_21_C245_n1384, Z => mult_21_C245_n872);
   mult_21_C245_U1155 : MUXB2DL port map( A0 => N3154, A1 => N3155, SL => 
                           mult_21_C245_n1384, Z => mult_21_C245_n873);
   mult_21_C245_U1154 : MUXB2DL port map( A0 => N3153, A1 => N3154, SL => 
                           mult_21_C245_n1384, Z => mult_21_C245_n874);
   mult_21_C245_U1153 : MUXB2DL port map( A0 => N3152, A1 => N3153, SL => 
                           mult_21_C245_n1384, Z => mult_21_C245_n875);
   mult_21_C245_U1152 : MUXB2DL port map( A0 => N3151, A1 => N3152, SL => 
                           mult_21_C245_n1384, Z => mult_21_C245_n876);
   mult_21_C245_U1151 : MUXB2DL port map( A0 => N3150, A1 => N3151, SL => 
                           mult_21_C245_n1384, Z => mult_21_C245_n877);
   mult_21_C245_U1150 : MUXB2DL port map( A0 => N3149, A1 => N3150, SL => 
                           mult_21_C245_n1384, Z => mult_21_C245_n878);
   mult_21_C245_U1149 : MUXB2DL port map( A0 => N3148, A1 => N3149, SL => 
                           mult_21_C245_n1384, Z => mult_21_C245_n879);
   mult_21_C245_U1148 : MUXB2DL port map( A0 => N3147, A1 => N3148, SL => 
                           mult_21_C245_n1384, Z => mult_21_C245_n880);
   mult_21_C245_U1147 : MUXB2DL port map( A0 => N3146, A1 => N3147, SL => 
                           mult_21_C245_n1384, Z => mult_21_C245_n881);
   mult_21_C245_U1146 : MUXB2DL port map( A0 => N3145, A1 => N3146, SL => 
                           mult_21_C245_n1384, Z => mult_21_C245_n882);
   mult_21_C245_U1145 : MUXB2DL port map( A0 => N3144, A1 => N3145, SL => 
                           mult_21_C245_n1384, Z => mult_21_C245_n883);
   mult_21_C245_U1144 : MUXB2DL port map( A0 => N3143, A1 => N3144, SL => 
                           mult_21_C245_n1384, Z => mult_21_C245_n884);
   mult_21_C245_U1143 : MUXB2DL port map( A0 => N3142, A1 => N3143, SL => 
                           mult_21_C245_n1384, Z => mult_21_C245_n885);
   mult_21_C245_U1142 : MUXB2DL port map( A0 => N3141, A1 => N3142, SL => 
                           mult_21_C245_n1384, Z => mult_21_C245_n886);
   mult_21_C245_U1141 : MUXB2DL port map( A0 => mult_21_C245_n1385, A1 => N3141
                           , SL => mult_21_C245_n1384, Z => mult_21_C245_n887);
   mult_21_C245_U1140 : MUXB2DL port map( A0 => N3139, A1 => N3140, SL => 
                           mult_21_C245_n1384, Z => mult_21_C245_n888);
   mult_21_C245_U1139 : MUXB2DL port map( A0 => mult_21_C245_n1387, A1 => N3139
                           , SL => mult_21_C245_n1384, Z => mult_21_C245_n889);
   mult_21_C245_U1138 : OAI21D1 port map( A1 => N3001, A2 => N3000, B => 
                           mult_21_C245_n1414, Z => mult_21_C245_n89);
   mult_21_C245_U1137 : MUXB2DL port map( A0 => N3137, A1 => N3138, SL => 
                           mult_21_C245_n1384, Z => mult_21_C245_n890);
   mult_21_C245_U1136 : NAN2D1 port map( A1 => N3137, A2 => mult_21_C245_n1384,
                           Z => mult_21_C245_n891);
   mult_21_C245_U1135 : MUXB2DL port map( A0 => N3167, A1 => N3168, SL => N2977
                           , Z => mult_21_C245_n892);
   mult_21_C245_U1134 : MUXB2DL port map( A0 => N3166, A1 => N3167, SL => N2977
                           , Z => mult_21_C245_n893);
   mult_21_C245_U1133 : MUXB2DL port map( A0 => N3165, A1 => N3166, SL => N2977
                           , Z => mult_21_C245_n894);
   mult_21_C245_U1132 : MUXB2DL port map( A0 => N3164, A1 => N3165, SL => N2977
                           , Z => mult_21_C245_n895);
   mult_21_C245_U1131 : MUXB2DL port map( A0 => N3163, A1 => N3164, SL => N2977
                           , Z => mult_21_C245_n896);
   mult_21_C245_U1130 : MUXB2DL port map( A0 => N3162, A1 => N3163, SL => N2977
                           , Z => mult_21_C245_n897);
   mult_21_C245_U1129 : MUXB2DL port map( A0 => N3161, A1 => N3162, SL => N2977
                           , Z => mult_21_C245_n898);
   mult_21_C245_U1128 : MUXB2DL port map( A0 => N3160, A1 => N3161, SL => N2977
                           , Z => mult_21_C245_n899);
   mult_21_C245_U1127 : MUXB2DL port map( A0 => N3159, A1 => N3160, SL => N2977
                           , Z => mult_21_C245_n900);
   mult_21_C245_U1126 : MUXB2DL port map( A0 => N3158, A1 => N3159, SL => N2977
                           , Z => mult_21_C245_n901);
   mult_21_C245_U1125 : MUXB2DL port map( A0 => N3157, A1 => N3158, SL => N2977
                           , Z => mult_21_C245_n902);
   mult_21_C245_U1124 : MUXB2DL port map( A0 => N3156, A1 => N3157, SL => N2977
                           , Z => mult_21_C245_n903);
   mult_21_C245_U1123 : MUXB2DL port map( A0 => N3155, A1 => N3156, SL => N2977
                           , Z => mult_21_C245_n904);
   mult_21_C245_U1122 : MUXB2DL port map( A0 => N3154, A1 => N3155, SL => N2977
                           , Z => mult_21_C245_n905);
   mult_21_C245_U1121 : MUXB2DL port map( A0 => N3153, A1 => N3154, SL => N2977
                           , Z => mult_21_C245_n906);
   mult_21_C245_U1120 : MUXB2DL port map( A0 => N3152, A1 => N3153, SL => N2977
                           , Z => mult_21_C245_n907);
   mult_21_C245_U1119 : MUXB2DL port map( A0 => N3151, A1 => N3152, SL => N2977
                           , Z => mult_21_C245_n908);
   mult_21_C245_U1118 : MUXB2DL port map( A0 => N3150, A1 => N3151, SL => N2977
                           , Z => mult_21_C245_n909);
   mult_21_C245_U1117 : AOI21D1 port map( A1 => N3000, A2 => N3001, B => 
                           mult_21_C245_n1414, Z => mult_21_C245_n942);
   mult_21_C245_U1116 : MUXB2DL port map( A0 => N3149, A1 => N3150, SL => N2977
                           , Z => mult_21_C245_n910);
   mult_21_C245_U1115 : MUXB2DL port map( A0 => N3148, A1 => N3149, SL => N2977
                           , Z => mult_21_C245_n911);
   mult_21_C245_U1114 : MUXB2DL port map( A0 => N3147, A1 => N3148, SL => N2977
                           , Z => mult_21_C245_n912);
   mult_21_C245_U1113 : MUXB2DL port map( A0 => N3146, A1 => N3147, SL => N2977
                           , Z => mult_21_C245_n913);
   mult_21_C245_U1112 : MUXB2DL port map( A0 => N3145, A1 => N3146, SL => N2977
                           , Z => mult_21_C245_n914);
   mult_21_C245_U1111 : MUXB2DL port map( A0 => N3144, A1 => N3145, SL => N2977
                           , Z => mult_21_C245_n915);
   mult_21_C245_U1110 : MUXB2DL port map( A0 => N3143, A1 => N3144, SL => N2977
                           , Z => mult_21_C245_n916);
   mult_21_C245_U1109 : MUXB2DL port map( A0 => N3142, A1 => N3143, SL => N2977
                           , Z => mult_21_C245_n917);
   mult_21_C245_U1108 : MUXB2DL port map( A0 => N3141, A1 => N3142, SL => N2977
                           , Z => mult_21_C245_n918);
   mult_21_C245_U1107 : MUXB2DL port map( A0 => mult_21_C245_n1385, A1 => N3141
                           , SL => N2977, Z => mult_21_C245_n919);
   mult_21_C245_U1106 : MUXB2DL port map( A0 => N3139, A1 => mult_21_C245_n1385
                           , SL => N2977, Z => mult_21_C245_n920);
   mult_21_C245_U1105 : MUXB2DL port map( A0 => mult_21_C245_n1387, A1 => N3139
                           , SL => N2977, Z => mult_21_C245_n921);
   mult_21_C245_U1104 : MUXB2DL port map( A0 => N3137, A1 => mult_21_C245_n1387
                           , SL => N2977, Z => mult_21_C245_n922);
   mult_21_C245_U1103 : NAN2D1 port map( A1 => N3137, A2 => N2977, Z => 
                           mult_21_C245_n923);
   mult_21_C245_U1102 : OAI21D1 port map( A1 => N3003, A2 => N3002, B => 
                           mult_21_C245_n1415, Z => mult_21_C245_n94);
   mult_21_C245_U1101 : AOI21D1 port map( A1 => N3002, A2 => N3003, B => 
                           mult_21_C245_n1415, Z => mult_21_C245_n941);
   mult_21_C245_U1100 : OAI21D1 port map( A1 => N3005, A2 => N3004, B => 
                           mult_21_C245_n1418, Z => mult_21_C245_n99);
   mult_21_C245_U1099 : EXOR2D1 port map( A1 => mult_21_C245_n230, A2 => 
                           mult_21_C245_n228, Z => mult_21_C245_n1437);
   mult_21_C245_U1098 : EXOR3D1 port map( A1 => mult_21_C245_n226, A2 => 
                           mult_21_C245_n224, A3 => mult_21_C245_n1437, Z => 
                           mult_21_C245_n1432);
   mult_21_C245_U1097 : EXOR2D1 port map( A1 => mult_21_C245_n222, A2 => 
                           mult_21_C245_n220, Z => mult_21_C245_n1436);
   mult_21_C245_U1096 : EXOR3D1 port map( A1 => mult_21_C245_n216, A2 => 
                           mult_21_C245_n1195, A3 => mult_21_C245_n1436, Z => 
                           mult_21_C245_n1433);
   mult_21_C245_U1095 : EXOR3D1 port map( A1 => mult_21_C245_n1165, A2 => 
                           mult_21_C245_n1137, A3 => mult_21_C245_n1045, Z => 
                           mult_21_C245_n1435);
   mult_21_C245_U1094 : EXOR3D1 port map( A1 => mult_21_C245_n1027, A2 => 
                           mult_21_C245_n1011, A3 => mult_21_C245_n1435, Z => 
                           mult_21_C245_n1434);
   mult_21_C245_U1093 : EXOR3D1 port map( A1 => mult_21_C245_n1432, A2 => 
                           mult_21_C245_n1433, A3 => mult_21_C245_n1434, Z => 
                           mult_21_C245_n1424);
   mult_21_C245_U1092 : EXOR2D1 port map( A1 => mult_21_C245_n985, A2 => 
                           mult_21_C245_n967, Z => mult_21_C245_n1431);
   mult_21_C245_U1091 : EXOR3D1 port map( A1 => mult_21_C245_n961, A2 => 
                           mult_21_C245_n218, A3 => mult_21_C245_n1431, Z => 
                           mult_21_C245_n1428);
   mult_21_C245_U1090 : EXNOR2D1 port map( A1 => mult_21_C245_n210, A2 => 
                           mult_21_C245_n1111, Z => mult_21_C245_n1430);
   mult_21_C245_U1089 : EXOR3D1 port map( A1 => mult_21_C245_n1087, A2 => 
                           mult_21_C245_n1065, A3 => mult_21_C245_n1430, Z => 
                           mult_21_C245_n1429);
   mult_21_C245_U1088 : EXOR3D1 port map( A1 => mult_21_C245_n1428, A2 => 
                           mult_21_C245_n204, A3 => mult_21_C245_n1429, Z => 
                           mult_21_C245_n1425);
   mult_21_C245_U1087 : EXNOR2D1 port map( A1 => mult_21_C245_n997, A2 => 
                           mult_21_C245_n975, Z => mult_21_C245_n1427);
   mult_21_C245_U1086 : EXOR3D1 port map( A1 => mult_21_C245_n957, A2 => 
                           mult_21_C245_n955, A3 => mult_21_C245_n1427, Z => 
                           mult_21_C245_n1426);
   mult_21_C245_U1085 : EXOR3D1 port map( A1 => mult_21_C245_n1424, A2 => 
                           mult_21_C245_n1425, A3 => mult_21_C245_n1426, Z => 
                           mult_21_C245_n1420);
   mult_21_C245_U1084 : EXOR2D1 port map( A1 => mult_21_C245_n202, A2 => 
                           mult_21_C245_n156, Z => mult_21_C245_n1421);
   mult_21_C245_U1083 : EXOR2D1 port map( A1 => mult_21_C245_n214, A2 => 
                           mult_21_C245_n212, Z => mult_21_C245_n1423);
   mult_21_C245_U1082 : EXOR3D1 port map( A1 => mult_21_C245_n208, A2 => 
                           mult_21_C245_n206, A3 => mult_21_C245_n1423, Z => 
                           mult_21_C245_n1422);
   mult_21_C245_U1081 : EXOR3D1 port map( A1 => mult_21_C245_n1420, A2 => 
                           mult_21_C245_n1421, A3 => mult_21_C245_n1422, Z => 
                           N3328);
   mult_21_C245_U1080 : INVD1 port map( A => N3008, Z => mult_21_C245_n1419);
   mult_21_C245_U1079 : INVD1 port map( A => N3140, Z => mult_21_C245_n1386);
   mult_21_C245_U1078 : INVD1 port map( A => N3138, Z => mult_21_C245_n1388);
   mult_21_C245_U1077 : MUXB2DL port map( A0 => N3166, A1 => N3165, SL => 
                           mult_21_C245_n1383, Z => mult_21_C245_n862);
   mult_21_C245_U1076 : INVD1 port map( A => N3006, Z => mult_21_C245_n1418);
   mult_21_C245_U1075 : INVD1 port map( A => N3004, Z => mult_21_C245_n1415);
   mult_21_C245_U1074 : INVD1 port map( A => N3002, Z => mult_21_C245_n1414);
   mult_21_C245_U1073 : OAI21D1 port map( A1 => N2999, A2 => N2998, B => 
                           mult_21_C245_n1412, Z => mult_21_C245_n84);
   mult_21_C245_U1072 : INVD1 port map( A => N3000, Z => mult_21_C245_n1412);
   mult_21_C245_U1071 : EXOR2D1 port map( A1 => N2999, A2 => N2998, Z => 
                           mult_21_C245_n1444);
   mult_21_C245_U1070 : OAI21D1 port map( A1 => N2997, A2 => N2996, B => 
                           mult_21_C245_n1410, Z => mult_21_C245_n80);
   mult_21_C245_U1069 : INVD1 port map( A => N2998, Z => mult_21_C245_n1410);
   mult_21_C245_U1068 : EXOR2D1 port map( A1 => N2997, A2 => N2996, Z => 
                           mult_21_C245_n1443);
   mult_21_C245_U1067 : OAI21D1 port map( A1 => N2995, A2 => N2994, B => 
                           mult_21_C245_n1408, Z => mult_21_C245_n73);
   mult_21_C245_U1066 : INVD1 port map( A => N2996, Z => mult_21_C245_n1408);
   mult_21_C245_U1065 : EXOR2D1 port map( A1 => N2995, A2 => N2994, Z => 
                           mult_21_C245_n1442);
   mult_21_C245_U1064 : OAI21D1 port map( A1 => N2993, A2 => N2992, B => 
                           mult_21_C245_n1406, Z => mult_21_C245_n66);
   mult_21_C245_U1063 : INVD1 port map( A => N2994, Z => mult_21_C245_n1406);
   mult_21_C245_U1062 : EXOR2D1 port map( A1 => N2993, A2 => N2992, Z => 
                           mult_21_C245_n1441);
   mult_21_C245_U1061 : OAI21D1 port map( A1 => N2991, A2 => N2990, B => 
                           mult_21_C245_n1404, Z => mult_21_C245_n58);
   mult_21_C245_U1060 : INVD1 port map( A => N2992, Z => mult_21_C245_n1404);
   mult_21_C245_U1059 : EXOR2D1 port map( A1 => N2991, A2 => N2990, Z => 
                           mult_21_C245_n1440);
   mult_21_C245_U1058 : OAI21D1 port map( A1 => N2989, A2 => N2988, B => 
                           mult_21_C245_n1402, Z => mult_21_C245_n50);
   mult_21_C245_U1057 : INVD1 port map( A => N2990, Z => mult_21_C245_n1402);
   mult_21_C245_U1056 : EXOR2D1 port map( A1 => N2989, A2 => N2988, Z => 
                           mult_21_C245_n1439);
   mult_21_C245_U1055 : OAI21D1 port map( A1 => N2986, A2 => N2987, B => 
                           mult_21_C245_n1400, Z => mult_21_C245_n42);
   mult_21_C245_U1054 : INVD1 port map( A => N2988, Z => mult_21_C245_n1400);
   mult_21_C245_U1053 : EXOR2D1 port map( A1 => N2987, A2 => N2986, Z => 
                           mult_21_C245_n1438);
   mult_21_C245_U1052 : INVD1 port map( A => N2986, Z => mult_21_C245_n1398);
   mult_21_C245_U1051 : INVD1 port map( A => N2984, Z => mult_21_C245_n1396);
   mult_21_C245_U1050 : INVD1 port map( A => N2982, Z => mult_21_C245_n1394);
   mult_21_C245_U1049 : INVD1 port map( A => N2980, Z => mult_21_C245_n1392);
   mult_21_C245_U1048 : INVD1 port map( A => mult_21_C245_n1386, Z => 
                           mult_21_C245_n1385);
   mult_21_C245_U1047 : INVD1 port map( A => mult_21_C245_n1388, Z => 
                           mult_21_C245_n1387);
   mult_21_C245_U1046 : EXNOR2D1 port map( A1 => N2979, A2 => N2978, Z => 
                           mult_21_C245_n1383);
   mult_21_C245_U1045 : INVD1 port map( A => N2978, Z => mult_21_C245_n1389);
   mult_21_C245_U1044 : INVD1 port map( A => mult_21_C245_n939, Z => 
                           mult_21_C245_n1417);
   mult_21_C245_U1043 : INVD1 port map( A => mult_21_C245_n940, Z => 
                           mult_21_C245_n1416);
   mult_21_C245_U1042 : INVD1 port map( A => mult_21_C245_n941, Z => 
                           mult_21_C245_n1413);
   mult_21_C245_U1041 : INVD1 port map( A => mult_21_C245_n942, Z => 
                           mult_21_C245_n1411);
   mult_21_C245_U1040 : INVD1 port map( A => mult_21_C245_n943, Z => 
                           mult_21_C245_n1409);
   mult_21_C245_U1039 : INVD1 port map( A => mult_21_C245_n944, Z => 
                           mult_21_C245_n1407);
   mult_21_C245_U1038 : INVD1 port map( A => mult_21_C245_n945, Z => 
                           mult_21_C245_n1405);
   mult_21_C245_U1037 : INVD1 port map( A => mult_21_C245_n946, Z => 
                           mult_21_C245_n1403);
   mult_21_C245_U1036 : INVD1 port map( A => mult_21_C245_n947, Z => 
                           mult_21_C245_n1401);
   mult_21_C245_U1035 : INVD1 port map( A => mult_21_C245_n948, Z => 
                           mult_21_C245_n1399);
   mult_21_C245_U1034 : INVD1 port map( A => mult_21_C245_n949, Z => 
                           mult_21_C245_n1397);
   mult_21_C245_U1033 : INVD1 port map( A => mult_21_C245_n950, Z => 
                           mult_21_C245_n1395);
   mult_21_C245_U1032 : INVD1 port map( A => mult_21_C245_n951, Z => 
                           mult_21_C245_n1393);
   mult_21_C245_U1031 : INVD1 port map( A => mult_21_C245_n952, Z => 
                           mult_21_C245_n1391);
   mult_21_C245_U1030 : INVD1 port map( A => mult_21_C245_n953, Z => 
                           mult_21_C245_n1390);
   mult_21_C245_U1029 : INVD1 port map( A => mult_21_C245_n1383, Z => 
                           mult_21_C245_n1384);
   mult_21_C245_U1028 : OAI21D1 port map( A1 => N2985, A2 => N2984, B => 
                           mult_21_C245_n1398, Z => mult_21_C245_n1382);
   mult_21_C245_U1027 : OAI21D1 port map( A1 => N2983, A2 => N2982, B => 
                           mult_21_C245_n1396, Z => mult_21_C245_n1381);
   mult_21_C245_U1026 : OAI21D1 port map( A1 => N2981, A2 => N2980, B => 
                           mult_21_C245_n1394, Z => mult_21_C245_n1380);
   mult_21_C245_U1025 : OAI21D1 port map( A1 => N2979, A2 => N2978, B => 
                           mult_21_C245_n1392, Z => mult_21_C245_n1379);
   mult_21_C245_U1024 : NAN2D1 port map( A1 => N2977, A2 => mult_21_C245_n1389,
                           Z => mult_21_C245_n1378);
   mult_21_C245_U1023 : EXOR2D1 port map( A1 => N2985, A2 => N2984, Z => 
                           mult_21_C245_n1377);
   mult_21_C245_U1022 : EXOR2D1 port map( A1 => N2983, A2 => N2982, Z => 
                           mult_21_C245_n1376);
   mult_21_C245_U1021 : EXOR2D1 port map( A1 => N2981, A2 => N2980, Z => 
                           mult_21_C245_n1375);
   mult_21_C245_U954 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n923, Z => 
                           mult_21_C245_n1226);
   mult_21_C245_U952 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n922, Z => 
                           mult_21_C245_n1225);
   mult_21_C245_U950 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n921, Z => 
                           mult_21_C245_n1224);
   mult_21_C245_U948 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n920, Z => 
                           mult_21_C245_n1223);
   mult_21_C245_U946 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n919, Z => 
                           mult_21_C245_n1222);
   mult_21_C245_U944 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n918, Z => 
                           mult_21_C245_n1221);
   mult_21_C245_U942 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n917, Z => 
                           mult_21_C245_n1220);
   mult_21_C245_U940 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n916, Z => 
                           mult_21_C245_n1219);
   mult_21_C245_U938 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n915, Z => 
                           mult_21_C245_n1218);
   mult_21_C245_U936 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n914, Z => 
                           mult_21_C245_n1217);
   mult_21_C245_U934 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n913, Z => 
                           mult_21_C245_n1216);
   mult_21_C245_U932 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n912, Z => 
                           mult_21_C245_n1215);
   mult_21_C245_U930 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n911, Z => 
                           mult_21_C245_n1214);
   mult_21_C245_U928 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n910, Z => 
                           mult_21_C245_n1213);
   mult_21_C245_U926 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n909, Z => 
                           mult_21_C245_n1212);
   mult_21_C245_U924 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n908, Z => 
                           mult_21_C245_n1211);
   mult_21_C245_U922 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n907, Z => 
                           mult_21_C245_n1210);
   mult_21_C245_U920 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n906, Z => 
                           mult_21_C245_n1209);
   mult_21_C245_U918 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n905, Z => 
                           mult_21_C245_n1208);
   mult_21_C245_U916 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n904, Z => 
                           mult_21_C245_n1207);
   mult_21_C245_U914 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n903, Z => 
                           mult_21_C245_n1206);
   mult_21_C245_U912 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n902, Z => 
                           mult_21_C245_n1205);
   mult_21_C245_U910 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n901, Z => 
                           mult_21_C245_n1204);
   mult_21_C245_U908 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n900, Z => 
                           mult_21_C245_n1203);
   mult_21_C245_U906 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n899, Z => 
                           mult_21_C245_n1202);
   mult_21_C245_U904 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n898, Z => 
                           mult_21_C245_n1201);
   mult_21_C245_U902 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n897, Z => 
                           mult_21_C245_n1200);
   mult_21_C245_U900 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n896, Z => 
                           mult_21_C245_n1199);
   mult_21_C245_U898 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n895, Z => 
                           mult_21_C245_n1198);
   mult_21_C245_U896 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n894, Z => 
                           mult_21_C245_n1197);
   mult_21_C245_U894 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n893, Z => 
                           mult_21_C245_n1196);
   mult_21_C245_U892 : MUXB2DL port map( A0 => mult_21_C245_n1378, A1 => 
                           mult_21_C245_n1389, SL => mult_21_C245_n892, Z => 
                           mult_21_C245_n1195);
   mult_21_C245_U889 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n891, Z => 
                           mult_21_C245_n1194);
   mult_21_C245_U887 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n890, Z => 
                           mult_21_C245_n1193);
   mult_21_C245_U885 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n889, Z => 
                           mult_21_C245_n1192);
   mult_21_C245_U883 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n888, Z => 
                           mult_21_C245_n1191);
   mult_21_C245_U881 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n887, Z => 
                           mult_21_C245_n1190);
   mult_21_C245_U879 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n886, Z => 
                           mult_21_C245_n1189);
   mult_21_C245_U877 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n885, Z => 
                           mult_21_C245_n1188);
   mult_21_C245_U875 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n884, Z => 
                           mult_21_C245_n1187);
   mult_21_C245_U873 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n883, Z => 
                           mult_21_C245_n1186);
   mult_21_C245_U871 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n882, Z => 
                           mult_21_C245_n1185);
   mult_21_C245_U869 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n881, Z => 
                           mult_21_C245_n1184);
   mult_21_C245_U867 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n880, Z => 
                           mult_21_C245_n1183);
   mult_21_C245_U865 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n879, Z => 
                           mult_21_C245_n1182);
   mult_21_C245_U863 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n878, Z => 
                           mult_21_C245_n1181);
   mult_21_C245_U861 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n877, Z => 
                           mult_21_C245_n1180);
   mult_21_C245_U859 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n876, Z => 
                           mult_21_C245_n1179);
   mult_21_C245_U857 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n875, Z => 
                           mult_21_C245_n1178);
   mult_21_C245_U855 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n874, Z => 
                           mult_21_C245_n1177);
   mult_21_C245_U853 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n873, Z => 
                           mult_21_C245_n1176);
   mult_21_C245_U851 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n872, Z => 
                           mult_21_C245_n1175);
   mult_21_C245_U849 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n871, Z => 
                           mult_21_C245_n1174);
   mult_21_C245_U847 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n870, Z => 
                           mult_21_C245_n1173);
   mult_21_C245_U845 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n869, Z => 
                           mult_21_C245_n1172);
   mult_21_C245_U843 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n868, Z => 
                           mult_21_C245_n1171);
   mult_21_C245_U841 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n867, Z => 
                           mult_21_C245_n1170);
   mult_21_C245_U839 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n866, Z => 
                           mult_21_C245_n1169);
   mult_21_C245_U837 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n865, Z => 
                           mult_21_C245_n1168);
   mult_21_C245_U835 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n864, Z => 
                           mult_21_C245_n1167);
   mult_21_C245_U833 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n863, Z => 
                           mult_21_C245_n1166);
   mult_21_C245_U831 : MUXB2DL port map( A0 => mult_21_C245_n1379, A1 => 
                           mult_21_C245_n1390, SL => mult_21_C245_n862, Z => 
                           mult_21_C245_n1165);
   mult_21_C245_U828 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n861, Z => 
                           mult_21_C245_n1164);
   mult_21_C245_U826 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n860, Z => 
                           mult_21_C245_n1163);
   mult_21_C245_U824 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n859, Z => 
                           mult_21_C245_n1162);
   mult_21_C245_U822 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n858, Z => 
                           mult_21_C245_n1161);
   mult_21_C245_U820 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n857, Z => 
                           mult_21_C245_n1160);
   mult_21_C245_U818 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n856, Z => 
                           mult_21_C245_n1159);
   mult_21_C245_U816 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n855, Z => 
                           mult_21_C245_n1158);
   mult_21_C245_U814 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n854, Z => 
                           mult_21_C245_n1157);
   mult_21_C245_U812 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n853, Z => 
                           mult_21_C245_n1156);
   mult_21_C245_U810 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n852, Z => 
                           mult_21_C245_n1155);
   mult_21_C245_U808 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n851, Z => 
                           mult_21_C245_n1154);
   mult_21_C245_U806 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n850, Z => 
                           mult_21_C245_n1153);
   mult_21_C245_U804 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n849, Z => 
                           mult_21_C245_n1152);
   mult_21_C245_U802 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n848, Z => 
                           mult_21_C245_n1151);
   mult_21_C245_U800 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n847, Z => 
                           mult_21_C245_n1150);
   mult_21_C245_U798 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n846, Z => 
                           mult_21_C245_n1149);
   mult_21_C245_U796 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n845, Z => 
                           mult_21_C245_n1148);
   mult_21_C245_U794 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n844, Z => 
                           mult_21_C245_n1147);
   mult_21_C245_U792 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n843, Z => 
                           mult_21_C245_n1146);
   mult_21_C245_U790 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n842, Z => 
                           mult_21_C245_n1145);
   mult_21_C245_U788 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n841, Z => 
                           mult_21_C245_n1144);
   mult_21_C245_U786 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n840, Z => 
                           mult_21_C245_n1143);
   mult_21_C245_U784 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n839, Z => 
                           mult_21_C245_n1142);
   mult_21_C245_U782 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n838, Z => 
                           mult_21_C245_n1141);
   mult_21_C245_U780 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n837, Z => 
                           mult_21_C245_n1140);
   mult_21_C245_U778 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n836, Z => 
                           mult_21_C245_n1139);
   mult_21_C245_U776 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n835, Z => 
                           mult_21_C245_n1138);
   mult_21_C245_U774 : MUXB2DL port map( A0 => mult_21_C245_n1380, A1 => 
                           mult_21_C245_n1391, SL => mult_21_C245_n834, Z => 
                           mult_21_C245_n1137);
   mult_21_C245_U771 : MUXB2DL port map( A0 => mult_21_C245_n1381, A1 => 
                           mult_21_C245_n1393, SL => mult_21_C245_n833, Z => 
                           mult_21_C245_n1136);
   mult_21_C245_U769 : MUXB2DL port map( A0 => mult_21_C245_n1381, A1 => 
                           mult_21_C245_n1393, SL => mult_21_C245_n832, Z => 
                           mult_21_C245_n1135);
   mult_21_C245_U767 : MUXB2DL port map( A0 => mult_21_C245_n1381, A1 => 
                           mult_21_C245_n1393, SL => mult_21_C245_n831, Z => 
                           mult_21_C245_n1134);
   mult_21_C245_U765 : MUXB2DL port map( A0 => mult_21_C245_n1381, A1 => 
                           mult_21_C245_n1393, SL => mult_21_C245_n830, Z => 
                           mult_21_C245_n1133);
   mult_21_C245_U763 : MUXB2DL port map( A0 => mult_21_C245_n1381, A1 => 
                           mult_21_C245_n1393, SL => mult_21_C245_n829, Z => 
                           mult_21_C245_n1132);
   mult_21_C245_U761 : MUXB2DL port map( A0 => mult_21_C245_n1381, A1 => 
                           mult_21_C245_n1393, SL => mult_21_C245_n828, Z => 
                           mult_21_C245_n1131);
   mult_21_C245_U759 : MUXB2DL port map( A0 => mult_21_C245_n1381, A1 => 
                           mult_21_C245_n1393, SL => mult_21_C245_n827, Z => 
                           mult_21_C245_n1130);
   mult_21_C245_U757 : MUXB2DL port map( A0 => mult_21_C245_n1381, A1 => 
                           mult_21_C245_n1393, SL => mult_21_C245_n826, Z => 
                           mult_21_C245_n1129);
   mult_21_C245_U755 : MUXB2DL port map( A0 => mult_21_C245_n1381, A1 => 
                           mult_21_C245_n1393, SL => mult_21_C245_n825, Z => 
                           mult_21_C245_n1128);
   mult_21_C245_U753 : MUXB2DL port map( A0 => mult_21_C245_n1381, A1 => 
                           mult_21_C245_n1393, SL => mult_21_C245_n824, Z => 
                           mult_21_C245_n1127);
   mult_21_C245_U751 : MUXB2DL port map( A0 => mult_21_C245_n1381, A1 => 
                           mult_21_C245_n1393, SL => mult_21_C245_n823, Z => 
                           mult_21_C245_n1126);
   mult_21_C245_U749 : MUXB2DL port map( A0 => mult_21_C245_n1381, A1 => 
                           mult_21_C245_n1393, SL => mult_21_C245_n822, Z => 
                           mult_21_C245_n1125);
   mult_21_C245_U747 : MUXB2DL port map( A0 => mult_21_C245_n1381, A1 => 
                           mult_21_C245_n1393, SL => mult_21_C245_n821, Z => 
                           mult_21_C245_n1124);
   mult_21_C245_U745 : MUXB2DL port map( A0 => mult_21_C245_n1381, A1 => 
                           mult_21_C245_n1393, SL => mult_21_C245_n820, Z => 
                           mult_21_C245_n1123);
   mult_21_C245_U743 : MUXB2DL port map( A0 => mult_21_C245_n1381, A1 => 
                           mult_21_C245_n1393, SL => mult_21_C245_n819, Z => 
                           mult_21_C245_n1122);
   mult_21_C245_U741 : MUXB2DL port map( A0 => mult_21_C245_n1381, A1 => 
                           mult_21_C245_n1393, SL => mult_21_C245_n818, Z => 
                           mult_21_C245_n1121);
   mult_21_C245_U739 : MUXB2DL port map( A0 => mult_21_C245_n1381, A1 => 
                           mult_21_C245_n1393, SL => mult_21_C245_n817, Z => 
                           mult_21_C245_n1120);
   mult_21_C245_U737 : MUXB2DL port map( A0 => mult_21_C245_n1381, A1 => 
                           mult_21_C245_n1393, SL => mult_21_C245_n816, Z => 
                           mult_21_C245_n1119);
   mult_21_C245_U735 : MUXB2DL port map( A0 => mult_21_C245_n1381, A1 => 
                           mult_21_C245_n1393, SL => mult_21_C245_n815, Z => 
                           mult_21_C245_n1118);
   mult_21_C245_U733 : MUXB2DL port map( A0 => mult_21_C245_n1381, A1 => 
                           mult_21_C245_n1393, SL => mult_21_C245_n814, Z => 
                           mult_21_C245_n1117);
   mult_21_C245_U731 : MUXB2DL port map( A0 => mult_21_C245_n1381, A1 => 
                           mult_21_C245_n1393, SL => mult_21_C245_n813, Z => 
                           mult_21_C245_n1116);
   mult_21_C245_U729 : MUXB2DL port map( A0 => mult_21_C245_n1381, A1 => 
                           mult_21_C245_n1393, SL => mult_21_C245_n812, Z => 
                           mult_21_C245_n1115);
   mult_21_C245_U727 : MUXB2DL port map( A0 => mult_21_C245_n1381, A1 => 
                           mult_21_C245_n1393, SL => mult_21_C245_n811, Z => 
                           mult_21_C245_n1114);
   mult_21_C245_U725 : MUXB2DL port map( A0 => mult_21_C245_n1381, A1 => 
                           mult_21_C245_n1393, SL => mult_21_C245_n810, Z => 
                           mult_21_C245_n1113);
   mult_21_C245_U723 : MUXB2DL port map( A0 => mult_21_C245_n1381, A1 => 
                           mult_21_C245_n1393, SL => mult_21_C245_n809, Z => 
                           mult_21_C245_n1112);
   mult_21_C245_U721 : MUXB2DL port map( A0 => mult_21_C245_n1381, A1 => 
                           mult_21_C245_n1393, SL => mult_21_C245_n808, Z => 
                           mult_21_C245_n1111);
   mult_21_C245_U718 : MUXB2DL port map( A0 => mult_21_C245_n1382, A1 => 
                           mult_21_C245_n1395, SL => mult_21_C245_n807, Z => 
                           mult_21_C245_n1110);
   mult_21_C245_U716 : MUXB2DL port map( A0 => mult_21_C245_n1382, A1 => 
                           mult_21_C245_n1395, SL => mult_21_C245_n806, Z => 
                           mult_21_C245_n1109);
   mult_21_C245_U714 : MUXB2DL port map( A0 => mult_21_C245_n1382, A1 => 
                           mult_21_C245_n1395, SL => mult_21_C245_n805, Z => 
                           mult_21_C245_n1108);
   mult_21_C245_U712 : MUXB2DL port map( A0 => mult_21_C245_n1382, A1 => 
                           mult_21_C245_n1395, SL => mult_21_C245_n804, Z => 
                           mult_21_C245_n1107);
   mult_21_C245_U710 : MUXB2DL port map( A0 => mult_21_C245_n1382, A1 => 
                           mult_21_C245_n1395, SL => mult_21_C245_n803, Z => 
                           mult_21_C245_n1106);
   mult_21_C245_U708 : MUXB2DL port map( A0 => mult_21_C245_n1382, A1 => 
                           mult_21_C245_n1395, SL => mult_21_C245_n802, Z => 
                           mult_21_C245_n1105);
   mult_21_C245_U706 : MUXB2DL port map( A0 => mult_21_C245_n1382, A1 => 
                           mult_21_C245_n1395, SL => mult_21_C245_n801, Z => 
                           mult_21_C245_n1104);
   mult_21_C245_U704 : MUXB2DL port map( A0 => mult_21_C245_n1382, A1 => 
                           mult_21_C245_n1395, SL => mult_21_C245_n800, Z => 
                           mult_21_C245_n1103);
   mult_21_C245_U702 : MUXB2DL port map( A0 => mult_21_C245_n1382, A1 => 
                           mult_21_C245_n1395, SL => mult_21_C245_n799, Z => 
                           mult_21_C245_n1102);
   mult_21_C245_U700 : MUXB2DL port map( A0 => mult_21_C245_n1382, A1 => 
                           mult_21_C245_n1395, SL => mult_21_C245_n798, Z => 
                           mult_21_C245_n1101);
   mult_21_C245_U698 : MUXB2DL port map( A0 => mult_21_C245_n1382, A1 => 
                           mult_21_C245_n1395, SL => mult_21_C245_n797, Z => 
                           mult_21_C245_n1100);
   mult_21_C245_U696 : MUXB2DL port map( A0 => mult_21_C245_n1382, A1 => 
                           mult_21_C245_n1395, SL => mult_21_C245_n796, Z => 
                           mult_21_C245_n1099);
   mult_21_C245_U694 : MUXB2DL port map( A0 => mult_21_C245_n1382, A1 => 
                           mult_21_C245_n1395, SL => mult_21_C245_n795, Z => 
                           mult_21_C245_n1098);
   mult_21_C245_U692 : MUXB2DL port map( A0 => mult_21_C245_n1382, A1 => 
                           mult_21_C245_n1395, SL => mult_21_C245_n794, Z => 
                           mult_21_C245_n1097);
   mult_21_C245_U690 : MUXB2DL port map( A0 => mult_21_C245_n1382, A1 => 
                           mult_21_C245_n1395, SL => mult_21_C245_n793, Z => 
                           mult_21_C245_n1096);
   mult_21_C245_U688 : MUXB2DL port map( A0 => mult_21_C245_n1382, A1 => 
                           mult_21_C245_n1395, SL => mult_21_C245_n792, Z => 
                           mult_21_C245_n1095);
   mult_21_C245_U686 : MUXB2DL port map( A0 => mult_21_C245_n1382, A1 => 
                           mult_21_C245_n1395, SL => mult_21_C245_n791, Z => 
                           mult_21_C245_n1094);
   mult_21_C245_U684 : MUXB2DL port map( A0 => mult_21_C245_n1382, A1 => 
                           mult_21_C245_n1395, SL => mult_21_C245_n790, Z => 
                           mult_21_C245_n1093);
   mult_21_C245_U682 : MUXB2DL port map( A0 => mult_21_C245_n1382, A1 => 
                           mult_21_C245_n1395, SL => mult_21_C245_n789, Z => 
                           mult_21_C245_n1092);
   mult_21_C245_U680 : MUXB2DL port map( A0 => mult_21_C245_n1382, A1 => 
                           mult_21_C245_n1395, SL => mult_21_C245_n788, Z => 
                           mult_21_C245_n1091);
   mult_21_C245_U678 : MUXB2DL port map( A0 => mult_21_C245_n1382, A1 => 
                           mult_21_C245_n1395, SL => mult_21_C245_n787, Z => 
                           mult_21_C245_n1090);
   mult_21_C245_U676 : MUXB2DL port map( A0 => mult_21_C245_n1382, A1 => 
                           mult_21_C245_n1395, SL => mult_21_C245_n786, Z => 
                           mult_21_C245_n1089);
   mult_21_C245_U674 : MUXB2DL port map( A0 => mult_21_C245_n1382, A1 => 
                           mult_21_C245_n1395, SL => mult_21_C245_n785, Z => 
                           mult_21_C245_n1088);
   mult_21_C245_U672 : MUXB2DL port map( A0 => mult_21_C245_n1382, A1 => 
                           mult_21_C245_n1395, SL => mult_21_C245_n784, Z => 
                           mult_21_C245_n1087);
   mult_21_C245_U669 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n1397, SL => mult_21_C245_n783, Z => 
                           mult_21_C245_n1086);
   mult_21_C245_U667 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n1397, SL => mult_21_C245_n782, Z => 
                           mult_21_C245_n1085);
   mult_21_C245_U665 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n1397, SL => mult_21_C245_n781, Z => 
                           mult_21_C245_n1084);
   mult_21_C245_U663 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n1397, SL => mult_21_C245_n780, Z => 
                           mult_21_C245_n1083);
   mult_21_C245_U661 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n1397, SL => mult_21_C245_n779, Z => 
                           mult_21_C245_n1082);
   mult_21_C245_U659 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n1397, SL => mult_21_C245_n778, Z => 
                           mult_21_C245_n1081);
   mult_21_C245_U657 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n1397, SL => mult_21_C245_n777, Z => 
                           mult_21_C245_n1080);
   mult_21_C245_U655 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n1397, SL => mult_21_C245_n776, Z => 
                           mult_21_C245_n1079);
   mult_21_C245_U653 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n1397, SL => mult_21_C245_n775, Z => 
                           mult_21_C245_n1078);
   mult_21_C245_U651 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n1397, SL => mult_21_C245_n774, Z => 
                           mult_21_C245_n1077);
   mult_21_C245_U649 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n1397, SL => mult_21_C245_n773, Z => 
                           mult_21_C245_n1076);
   mult_21_C245_U647 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n1397, SL => mult_21_C245_n772, Z => 
                           mult_21_C245_n1075);
   mult_21_C245_U645 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n1397, SL => mult_21_C245_n771, Z => 
                           mult_21_C245_n1074);
   mult_21_C245_U643 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n1397, SL => mult_21_C245_n770, Z => 
                           mult_21_C245_n1073);
   mult_21_C245_U641 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n1397, SL => mult_21_C245_n769, Z => 
                           mult_21_C245_n1072);
   mult_21_C245_U639 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n1397, SL => mult_21_C245_n768, Z => 
                           mult_21_C245_n1071);
   mult_21_C245_U637 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n1397, SL => mult_21_C245_n767, Z => 
                           mult_21_C245_n1070);
   mult_21_C245_U635 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n1397, SL => mult_21_C245_n766, Z => 
                           mult_21_C245_n1069);
   mult_21_C245_U633 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n1397, SL => mult_21_C245_n765, Z => 
                           mult_21_C245_n1068);
   mult_21_C245_U631 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n1397, SL => mult_21_C245_n764, Z => 
                           mult_21_C245_n1067);
   mult_21_C245_U629 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n1397, SL => mult_21_C245_n763, Z => 
                           mult_21_C245_n1066);
   mult_21_C245_U627 : MUXB2DL port map( A0 => mult_21_C245_n42, A1 => 
                           mult_21_C245_n1397, SL => mult_21_C245_n762, Z => 
                           mult_21_C245_n1065);
   mult_21_C245_U624 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n1399, SL => mult_21_C245_n761, Z => 
                           mult_21_C245_n1064);
   mult_21_C245_U622 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n1399, SL => mult_21_C245_n760, Z => 
                           mult_21_C245_n1063);
   mult_21_C245_U620 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n1399, SL => mult_21_C245_n759, Z => 
                           mult_21_C245_n1062);
   mult_21_C245_U618 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n1399, SL => mult_21_C245_n758, Z => 
                           mult_21_C245_n1061);
   mult_21_C245_U616 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n1399, SL => mult_21_C245_n757, Z => 
                           mult_21_C245_n1060);
   mult_21_C245_U614 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n1399, SL => mult_21_C245_n756, Z => 
                           mult_21_C245_n1059);
   mult_21_C245_U612 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n1399, SL => mult_21_C245_n755, Z => 
                           mult_21_C245_n1058);
   mult_21_C245_U610 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n1399, SL => mult_21_C245_n754, Z => 
                           mult_21_C245_n1057);
   mult_21_C245_U608 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n1399, SL => mult_21_C245_n753, Z => 
                           mult_21_C245_n1056);
   mult_21_C245_U606 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n1399, SL => mult_21_C245_n752, Z => 
                           mult_21_C245_n1055);
   mult_21_C245_U604 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n1399, SL => mult_21_C245_n751, Z => 
                           mult_21_C245_n1054);
   mult_21_C245_U602 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n1399, SL => mult_21_C245_n750, Z => 
                           mult_21_C245_n1053);
   mult_21_C245_U600 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n1399, SL => mult_21_C245_n749, Z => 
                           mult_21_C245_n1052);
   mult_21_C245_U598 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n1399, SL => mult_21_C245_n748, Z => 
                           mult_21_C245_n1051);
   mult_21_C245_U596 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n1399, SL => mult_21_C245_n747, Z => 
                           mult_21_C245_n1050);
   mult_21_C245_U594 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n1399, SL => mult_21_C245_n746, Z => 
                           mult_21_C245_n1049);
   mult_21_C245_U592 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n1399, SL => mult_21_C245_n745, Z => 
                           mult_21_C245_n1048);
   mult_21_C245_U590 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n1399, SL => mult_21_C245_n744, Z => 
                           mult_21_C245_n1047);
   mult_21_C245_U588 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n1399, SL => mult_21_C245_n743, Z => 
                           mult_21_C245_n1046);
   mult_21_C245_U586 : MUXB2DL port map( A0 => mult_21_C245_n50, A1 => 
                           mult_21_C245_n1399, SL => mult_21_C245_n742, Z => 
                           mult_21_C245_n1045);
   mult_21_C245_U583 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n1401, SL => mult_21_C245_n741, Z => 
                           mult_21_C245_n1044);
   mult_21_C245_U581 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n1401, SL => mult_21_C245_n740, Z => 
                           mult_21_C245_n1043);
   mult_21_C245_U579 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n1401, SL => mult_21_C245_n739, Z => 
                           mult_21_C245_n1042);
   mult_21_C245_U577 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n1401, SL => mult_21_C245_n738, Z => 
                           mult_21_C245_n1041);
   mult_21_C245_U575 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n1401, SL => mult_21_C245_n737, Z => 
                           mult_21_C245_n1040);
   mult_21_C245_U573 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n1401, SL => mult_21_C245_n736, Z => 
                           mult_21_C245_n1039);
   mult_21_C245_U571 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n1401, SL => mult_21_C245_n735, Z => 
                           mult_21_C245_n1038);
   mult_21_C245_U569 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n1401, SL => mult_21_C245_n734, Z => 
                           mult_21_C245_n1037);
   mult_21_C245_U567 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n1401, SL => mult_21_C245_n733, Z => 
                           mult_21_C245_n1036);
   mult_21_C245_U565 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n1401, SL => mult_21_C245_n732, Z => 
                           mult_21_C245_n1035);
   mult_21_C245_U563 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n1401, SL => mult_21_C245_n731, Z => 
                           mult_21_C245_n1034);
   mult_21_C245_U561 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n1401, SL => mult_21_C245_n730, Z => 
                           mult_21_C245_n1033);
   mult_21_C245_U559 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n1401, SL => mult_21_C245_n729, Z => 
                           mult_21_C245_n1032);
   mult_21_C245_U557 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n1401, SL => mult_21_C245_n728, Z => 
                           mult_21_C245_n1031);
   mult_21_C245_U555 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n1401, SL => mult_21_C245_n727, Z => 
                           mult_21_C245_n1030);
   mult_21_C245_U553 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n1401, SL => mult_21_C245_n726, Z => 
                           mult_21_C245_n1029);
   mult_21_C245_U551 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n1401, SL => mult_21_C245_n725, Z => 
                           mult_21_C245_n1028);
   mult_21_C245_U549 : MUXB2DL port map( A0 => mult_21_C245_n58, A1 => 
                           mult_21_C245_n1401, SL => mult_21_C245_n724, Z => 
                           mult_21_C245_n1027);
   mult_21_C245_U546 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n1403, SL => mult_21_C245_n723, Z => 
                           mult_21_C245_n1026);
   mult_21_C245_U544 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n1403, SL => mult_21_C245_n722, Z => 
                           mult_21_C245_n1025);
   mult_21_C245_U542 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n1403, SL => mult_21_C245_n721, Z => 
                           mult_21_C245_n1024);
   mult_21_C245_U540 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n1403, SL => mult_21_C245_n720, Z => 
                           mult_21_C245_n1023);
   mult_21_C245_U538 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n1403, SL => mult_21_C245_n719, Z => 
                           mult_21_C245_n1022);
   mult_21_C245_U536 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n1403, SL => mult_21_C245_n718, Z => 
                           mult_21_C245_n1021);
   mult_21_C245_U534 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n1403, SL => mult_21_C245_n717, Z => 
                           mult_21_C245_n1020);
   mult_21_C245_U532 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n1403, SL => mult_21_C245_n716, Z => 
                           mult_21_C245_n1019);
   mult_21_C245_U530 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n1403, SL => mult_21_C245_n715, Z => 
                           mult_21_C245_n1018);
   mult_21_C245_U528 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n1403, SL => mult_21_C245_n714, Z => 
                           mult_21_C245_n1017);
   mult_21_C245_U526 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n1403, SL => mult_21_C245_n713, Z => 
                           mult_21_C245_n1016);
   mult_21_C245_U524 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n1403, SL => mult_21_C245_n712, Z => 
                           mult_21_C245_n1015);
   mult_21_C245_U522 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n1403, SL => mult_21_C245_n711, Z => 
                           mult_21_C245_n1014);
   mult_21_C245_U520 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n1403, SL => mult_21_C245_n710, Z => 
                           mult_21_C245_n1013);
   mult_21_C245_U518 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n1403, SL => mult_21_C245_n709, Z => 
                           mult_21_C245_n1012);
   mult_21_C245_U516 : MUXB2DL port map( A0 => mult_21_C245_n66, A1 => 
                           mult_21_C245_n1403, SL => mult_21_C245_n708, Z => 
                           mult_21_C245_n1011);
   mult_21_C245_U513 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n1405, SL => mult_21_C245_n707, Z => 
                           mult_21_C245_n1010);
   mult_21_C245_U511 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n1405, SL => mult_21_C245_n706, Z => 
                           mult_21_C245_n1009);
   mult_21_C245_U509 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n1405, SL => mult_21_C245_n705, Z => 
                           mult_21_C245_n1008);
   mult_21_C245_U507 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n1405, SL => mult_21_C245_n704, Z => 
                           mult_21_C245_n1007);
   mult_21_C245_U505 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n1405, SL => mult_21_C245_n703, Z => 
                           mult_21_C245_n1006);
   mult_21_C245_U503 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n1405, SL => mult_21_C245_n702, Z => 
                           mult_21_C245_n1005);
   mult_21_C245_U501 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n1405, SL => mult_21_C245_n701, Z => 
                           mult_21_C245_n1004);
   mult_21_C245_U499 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n1405, SL => mult_21_C245_n700, Z => 
                           mult_21_C245_n1003);
   mult_21_C245_U497 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n1405, SL => mult_21_C245_n699, Z => 
                           mult_21_C245_n1002);
   mult_21_C245_U495 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n1405, SL => mult_21_C245_n698, Z => 
                           mult_21_C245_n1001);
   mult_21_C245_U493 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n1405, SL => mult_21_C245_n697, Z => 
                           mult_21_C245_n1000);
   mult_21_C245_U491 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n1405, SL => mult_21_C245_n696, Z => 
                           mult_21_C245_n999);
   mult_21_C245_U489 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n1405, SL => mult_21_C245_n695, Z => 
                           mult_21_C245_n998);
   mult_21_C245_U487 : MUXB2DL port map( A0 => mult_21_C245_n73, A1 => 
                           mult_21_C245_n1405, SL => mult_21_C245_n694, Z => 
                           mult_21_C245_n997);
   mult_21_C245_U484 : MUXB2DL port map( A0 => mult_21_C245_n80, A1 => 
                           mult_21_C245_n1407, SL => mult_21_C245_n693, Z => 
                           mult_21_C245_n996);
   mult_21_C245_U482 : MUXB2DL port map( A0 => mult_21_C245_n80, A1 => 
                           mult_21_C245_n1407, SL => mult_21_C245_n692, Z => 
                           mult_21_C245_n995);
   mult_21_C245_U480 : MUXB2DL port map( A0 => mult_21_C245_n80, A1 => 
                           mult_21_C245_n1407, SL => mult_21_C245_n691, Z => 
                           mult_21_C245_n994);
   mult_21_C245_U478 : MUXB2DL port map( A0 => mult_21_C245_n80, A1 => 
                           mult_21_C245_n1407, SL => mult_21_C245_n690, Z => 
                           mult_21_C245_n993);
   mult_21_C245_U476 : MUXB2DL port map( A0 => mult_21_C245_n80, A1 => 
                           mult_21_C245_n1407, SL => mult_21_C245_n689, Z => 
                           mult_21_C245_n992);
   mult_21_C245_U474 : MUXB2DL port map( A0 => mult_21_C245_n80, A1 => 
                           mult_21_C245_n1407, SL => mult_21_C245_n688, Z => 
                           mult_21_C245_n991);
   mult_21_C245_U472 : MUXB2DL port map( A0 => mult_21_C245_n80, A1 => 
                           mult_21_C245_n1407, SL => mult_21_C245_n687, Z => 
                           mult_21_C245_n990);
   mult_21_C245_U470 : MUXB2DL port map( A0 => mult_21_C245_n80, A1 => 
                           mult_21_C245_n1407, SL => mult_21_C245_n686, Z => 
                           mult_21_C245_n989);
   mult_21_C245_U468 : MUXB2DL port map( A0 => mult_21_C245_n80, A1 => 
                           mult_21_C245_n1407, SL => mult_21_C245_n685, Z => 
                           mult_21_C245_n988);
   mult_21_C245_U466 : MUXB2DL port map( A0 => mult_21_C245_n80, A1 => 
                           mult_21_C245_n1407, SL => mult_21_C245_n684, Z => 
                           mult_21_C245_n987);
   mult_21_C245_U464 : MUXB2DL port map( A0 => mult_21_C245_n80, A1 => 
                           mult_21_C245_n1407, SL => mult_21_C245_n683, Z => 
                           mult_21_C245_n986);
   mult_21_C245_U462 : MUXB2DL port map( A0 => mult_21_C245_n80, A1 => 
                           mult_21_C245_n1407, SL => mult_21_C245_n682, Z => 
                           mult_21_C245_n985);
   mult_21_C245_U459 : MUXB2DL port map( A0 => mult_21_C245_n84, A1 => 
                           mult_21_C245_n1409, SL => mult_21_C245_n681, Z => 
                           mult_21_C245_n984);
   mult_21_C245_U457 : MUXB2DL port map( A0 => mult_21_C245_n84, A1 => 
                           mult_21_C245_n1409, SL => mult_21_C245_n680, Z => 
                           mult_21_C245_n983);
   mult_21_C245_U455 : MUXB2DL port map( A0 => mult_21_C245_n84, A1 => 
                           mult_21_C245_n1409, SL => mult_21_C245_n679, Z => 
                           mult_21_C245_n982);
   mult_21_C245_U453 : MUXB2DL port map( A0 => mult_21_C245_n84, A1 => 
                           mult_21_C245_n1409, SL => mult_21_C245_n678, Z => 
                           mult_21_C245_n981);
   mult_21_C245_U451 : MUXB2DL port map( A0 => mult_21_C245_n84, A1 => 
                           mult_21_C245_n1409, SL => mult_21_C245_n677, Z => 
                           mult_21_C245_n980);
   mult_21_C245_U449 : MUXB2DL port map( A0 => mult_21_C245_n84, A1 => 
                           mult_21_C245_n1409, SL => mult_21_C245_n676, Z => 
                           mult_21_C245_n979);
   mult_21_C245_U447 : MUXB2DL port map( A0 => mult_21_C245_n84, A1 => 
                           mult_21_C245_n1409, SL => mult_21_C245_n675, Z => 
                           mult_21_C245_n978);
   mult_21_C245_U445 : MUXB2DL port map( A0 => mult_21_C245_n84, A1 => 
                           mult_21_C245_n1409, SL => mult_21_C245_n674, Z => 
                           mult_21_C245_n977);
   mult_21_C245_U443 : MUXB2DL port map( A0 => mult_21_C245_n84, A1 => 
                           mult_21_C245_n1409, SL => mult_21_C245_n673, Z => 
                           mult_21_C245_n976);
   mult_21_C245_U441 : MUXB2DL port map( A0 => mult_21_C245_n84, A1 => 
                           mult_21_C245_n1409, SL => mult_21_C245_n672, Z => 
                           mult_21_C245_n975);
   mult_21_C245_U438 : MUXB2DL port map( A0 => mult_21_C245_n89, A1 => 
                           mult_21_C245_n1411, SL => mult_21_C245_n671, Z => 
                           mult_21_C245_n974);
   mult_21_C245_U436 : MUXB2DL port map( A0 => mult_21_C245_n89, A1 => 
                           mult_21_C245_n1411, SL => mult_21_C245_n670, Z => 
                           mult_21_C245_n973);
   mult_21_C245_U434 : MUXB2DL port map( A0 => mult_21_C245_n89, A1 => 
                           mult_21_C245_n1411, SL => mult_21_C245_n669, Z => 
                           mult_21_C245_n972);
   mult_21_C245_U432 : MUXB2DL port map( A0 => mult_21_C245_n89, A1 => 
                           mult_21_C245_n1411, SL => mult_21_C245_n668, Z => 
                           mult_21_C245_n971);
   mult_21_C245_U430 : MUXB2DL port map( A0 => mult_21_C245_n89, A1 => 
                           mult_21_C245_n1411, SL => mult_21_C245_n667, Z => 
                           mult_21_C245_n970);
   mult_21_C245_U428 : MUXB2DL port map( A0 => mult_21_C245_n89, A1 => 
                           mult_21_C245_n1411, SL => mult_21_C245_n666, Z => 
                           mult_21_C245_n969);
   mult_21_C245_U426 : MUXB2DL port map( A0 => mult_21_C245_n89, A1 => 
                           mult_21_C245_n1411, SL => mult_21_C245_n665, Z => 
                           mult_21_C245_n968);
   mult_21_C245_U424 : MUXB2DL port map( A0 => mult_21_C245_n89, A1 => 
                           mult_21_C245_n1411, SL => mult_21_C245_n664, Z => 
                           mult_21_C245_n967);
   mult_21_C245_U421 : MUXB2DL port map( A0 => mult_21_C245_n94, A1 => 
                           mult_21_C245_n1413, SL => mult_21_C245_n663, Z => 
                           mult_21_C245_n966);
   mult_21_C245_U419 : MUXB2DL port map( A0 => mult_21_C245_n94, A1 => 
                           mult_21_C245_n1413, SL => mult_21_C245_n662, Z => 
                           mult_21_C245_n965);
   mult_21_C245_U417 : MUXB2DL port map( A0 => mult_21_C245_n94, A1 => 
                           mult_21_C245_n1413, SL => mult_21_C245_n661, Z => 
                           mult_21_C245_n964);
   mult_21_C245_U415 : MUXB2DL port map( A0 => mult_21_C245_n94, A1 => 
                           mult_21_C245_n1413, SL => mult_21_C245_n660, Z => 
                           mult_21_C245_n963);
   mult_21_C245_U413 : MUXB2DL port map( A0 => mult_21_C245_n94, A1 => 
                           mult_21_C245_n1413, SL => mult_21_C245_n659, Z => 
                           mult_21_C245_n962);
   mult_21_C245_U411 : MUXB2DL port map( A0 => mult_21_C245_n94, A1 => 
                           mult_21_C245_n1413, SL => mult_21_C245_n658, Z => 
                           mult_21_C245_n961);
   mult_21_C245_U408 : MUXB2DL port map( A0 => mult_21_C245_n99, A1 => 
                           mult_21_C245_n1416, SL => mult_21_C245_n657, Z => 
                           mult_21_C245_n960);
   mult_21_C245_U406 : MUXB2DL port map( A0 => mult_21_C245_n99, A1 => 
                           mult_21_C245_n1416, SL => mult_21_C245_n656, Z => 
                           mult_21_C245_n959);
   mult_21_C245_U404 : MUXB2DL port map( A0 => mult_21_C245_n99, A1 => 
                           mult_21_C245_n1416, SL => mult_21_C245_n655, Z => 
                           mult_21_C245_n958);
   mult_21_C245_U402 : MUXB2DL port map( A0 => mult_21_C245_n99, A1 => 
                           mult_21_C245_n1416, SL => mult_21_C245_n654, Z => 
                           mult_21_C245_n957);
   mult_21_C245_U399 : MUXB2DL port map( A0 => mult_21_C245_n104, A1 => 
                           mult_21_C245_n1417, SL => mult_21_C245_n653, Z => 
                           mult_21_C245_n956);
   mult_21_C245_U397 : MUXB2DL port map( A0 => mult_21_C245_n104, A1 => 
                           mult_21_C245_n1417, SL => mult_21_C245_n652, Z => 
                           mult_21_C245_n955);
   mult_21_C245_U395 : ADHALFDL port map( A => mult_21_C245_n1224, B => 
                           mult_21_C245_n953, CO => mult_21_C245_n650, S => 
                           mult_21_C245_n651);
   mult_21_C245_U394 : ADHALFDL port map( A => mult_21_C245_n650, B => 
                           mult_21_C245_n1223, CO => mult_21_C245_n648, S => 
                           mult_21_C245_n649);
   mult_21_C245_U393 : ADHALFDL port map( A => mult_21_C245_n1222, B => 
                           mult_21_C245_n952, CO => mult_21_C245_n646, S => 
                           mult_21_C245_n647);
   mult_21_C245_U392 : ADFULD1 port map( A => mult_21_C245_n1192, B => 
                           mult_21_C245_n1164, CI => mult_21_C245_n647, CO => 
                           mult_21_C245_n644, S => mult_21_C245_n645);
   mult_21_C245_U391 : ADHALFDL port map( A => mult_21_C245_n646, B => 
                           mult_21_C245_n1221, CO => mult_21_C245_n642, S => 
                           mult_21_C245_n643);
   mult_21_C245_U390 : ADFULD1 port map( A => mult_21_C245_n1163, B => 
                           mult_21_C245_n1191, CI => mult_21_C245_n643, CO => 
                           mult_21_C245_n640, S => mult_21_C245_n641);
   mult_21_C245_U389 : ADHALFDL port map( A => mult_21_C245_n1220, B => 
                           mult_21_C245_n951, CO => mult_21_C245_n638, S => 
                           mult_21_C245_n639);
   mult_21_C245_U388 : ADFULD1 port map( A => mult_21_C245_n1190, B => 
                           mult_21_C245_n1136, CI => mult_21_C245_n1162, CO => 
                           mult_21_C245_n636, S => mult_21_C245_n637);
   mult_21_C245_U387 : ADFULD1 port map( A => mult_21_C245_n642, B => 
                           mult_21_C245_n639, CI => mult_21_C245_n637, CO => 
                           mult_21_C245_n634, S => mult_21_C245_n635);
   mult_21_C245_U386 : ADHALFDL port map( A => mult_21_C245_n638, B => 
                           mult_21_C245_n1219, CO => mult_21_C245_n632, S => 
                           mult_21_C245_n633);
   mult_21_C245_U385 : ADFULD1 port map( A => mult_21_C245_n1135, B => 
                           mult_21_C245_n1189, CI => mult_21_C245_n1161, CO => 
                           mult_21_C245_n630, S => mult_21_C245_n631);
   mult_21_C245_U384 : ADFULD1 port map( A => mult_21_C245_n636, B => 
                           mult_21_C245_n633, CI => mult_21_C245_n631, CO => 
                           mult_21_C245_n628, S => mult_21_C245_n629);
   mult_21_C245_U383 : ADHALFDL port map( A => mult_21_C245_n1218, B => 
                           mult_21_C245_n950, CO => mult_21_C245_n626, S => 
                           mult_21_C245_n627);
   mult_21_C245_U382 : ADFULD1 port map( A => mult_21_C245_n1188, B => 
                           mult_21_C245_n1110, CI => mult_21_C245_n1134, CO => 
                           mult_21_C245_n624, S => mult_21_C245_n625);
   mult_21_C245_U381 : ADFULD1 port map( A => mult_21_C245_n627, B => 
                           mult_21_C245_n1160, CI => mult_21_C245_n632, CO => 
                           mult_21_C245_n622, S => mult_21_C245_n623);
   mult_21_C245_U380 : ADFULD1 port map( A => mult_21_C245_n625, B => 
                           mult_21_C245_n630, CI => mult_21_C245_n623, CO => 
                           mult_21_C245_n620, S => mult_21_C245_n621);
   mult_21_C245_U379 : ADHALFDL port map( A => mult_21_C245_n626, B => 
                           mult_21_C245_n1217, CO => mult_21_C245_n618, S => 
                           mult_21_C245_n619);
   mult_21_C245_U378 : ADFULD1 port map( A => mult_21_C245_n1109, B => 
                           mult_21_C245_n1133, CI => mult_21_C245_n1159, CO => 
                           mult_21_C245_n616, S => mult_21_C245_n617);
   mult_21_C245_U377 : ADFULD1 port map( A => mult_21_C245_n619, B => 
                           mult_21_C245_n1187, CI => mult_21_C245_n624, CO => 
                           mult_21_C245_n614, S => mult_21_C245_n615);
   mult_21_C245_U376 : ADFULD1 port map( A => mult_21_C245_n617, B => 
                           mult_21_C245_n622, CI => mult_21_C245_n615, CO => 
                           mult_21_C245_n612, S => mult_21_C245_n613);
   mult_21_C245_U375 : ADHALFDL port map( A => mult_21_C245_n1216, B => 
                           mult_21_C245_n949, CO => mult_21_C245_n610, S => 
                           mult_21_C245_n611);
   mult_21_C245_U374 : ADFULD1 port map( A => mult_21_C245_n1132, B => 
                           mult_21_C245_n1086, CI => mult_21_C245_n1186, CO => 
                           mult_21_C245_n608, S => mult_21_C245_n609);
   mult_21_C245_U373 : ADFULD1 port map( A => mult_21_C245_n1108, B => 
                           mult_21_C245_n1158, CI => mult_21_C245_n611, CO => 
                           mult_21_C245_n606, S => mult_21_C245_n607);
   mult_21_C245_U372 : ADFULD1 port map( A => mult_21_C245_n616, B => 
                           mult_21_C245_n618, CI => mult_21_C245_n609, CO => 
                           mult_21_C245_n604, S => mult_21_C245_n605);
   mult_21_C245_U371 : ADFULD1 port map( A => mult_21_C245_n614, B => 
                           mult_21_C245_n607, CI => mult_21_C245_n605, CO => 
                           mult_21_C245_n602, S => mult_21_C245_n603);
   mult_21_C245_U370 : ADHALFDL port map( A => mult_21_C245_n610, B => 
                           mult_21_C245_n1215, CO => mult_21_C245_n600, S => 
                           mult_21_C245_n601);
   mult_21_C245_U369 : ADFULD1 port map( A => mult_21_C245_n1085, B => 
                           mult_21_C245_n1131, CI => mult_21_C245_n1185, CO => 
                           mult_21_C245_n598, S => mult_21_C245_n599);
   mult_21_C245_U368 : ADFULD1 port map( A => mult_21_C245_n1107, B => 
                           mult_21_C245_n1157, CI => mult_21_C245_n601, CO => 
                           mult_21_C245_n596, S => mult_21_C245_n597);
   mult_21_C245_U367 : ADFULD1 port map( A => mult_21_C245_n606, B => 
                           mult_21_C245_n608, CI => mult_21_C245_n599, CO => 
                           mult_21_C245_n594, S => mult_21_C245_n595);
   mult_21_C245_U366 : ADFULD1 port map( A => mult_21_C245_n604, B => 
                           mult_21_C245_n597, CI => mult_21_C245_n595, CO => 
                           mult_21_C245_n592, S => mult_21_C245_n593);
   mult_21_C245_U365 : ADHALFDL port map( A => mult_21_C245_n1214, B => 
                           mult_21_C245_n948, CO => mult_21_C245_n590, S => 
                           mult_21_C245_n591);
   mult_21_C245_U364 : ADFULD1 port map( A => mult_21_C245_n1130, B => 
                           mult_21_C245_n1064, CI => mult_21_C245_n1184, CO => 
                           mult_21_C245_n588, S => mult_21_C245_n589);
   mult_21_C245_U363 : ADFULD1 port map( A => mult_21_C245_n1084, B => 
                           mult_21_C245_n1156, CI => mult_21_C245_n591, CO => 
                           mult_21_C245_n586, S => mult_21_C245_n587);
   mult_21_C245_U362 : ADFULD1 port map( A => mult_21_C245_n600, B => 
                           mult_21_C245_n1106, CI => mult_21_C245_n598, CO => 
                           mult_21_C245_n584, S => mult_21_C245_n585);
   mult_21_C245_U361 : ADFULD1 port map( A => mult_21_C245_n587, B => 
                           mult_21_C245_n589, CI => mult_21_C245_n596, CO => 
                           mult_21_C245_n582, S => mult_21_C245_n583);
   mult_21_C245_U360 : ADFULD1 port map( A => mult_21_C245_n585, B => 
                           mult_21_C245_n594, CI => mult_21_C245_n583, CO => 
                           mult_21_C245_n580, S => mult_21_C245_n581);
   mult_21_C245_U359 : ADHALFDL port map( A => mult_21_C245_n590, B => 
                           mult_21_C245_n1213, CO => mult_21_C245_n578, S => 
                           mult_21_C245_n579);
   mult_21_C245_U358 : ADFULD1 port map( A => mult_21_C245_n1183, B => 
                           mult_21_C245_n1105, CI => mult_21_C245_n1155, CO => 
                           mult_21_C245_n576, S => mult_21_C245_n577);
   mult_21_C245_U357 : ADFULD1 port map( A => mult_21_C245_n1063, B => 
                           mult_21_C245_n1129, CI => mult_21_C245_n1083, CO => 
                           mult_21_C245_n574, S => mult_21_C245_n575);
   mult_21_C245_U356 : ADFULD1 port map( A => mult_21_C245_n588, B => 
                           mult_21_C245_n579, CI => mult_21_C245_n586, CO => 
                           mult_21_C245_n572, S => mult_21_C245_n573);
   mult_21_C245_U355 : ADFULD1 port map( A => mult_21_C245_n577, B => 
                           mult_21_C245_n575, CI => mult_21_C245_n584, CO => 
                           mult_21_C245_n570, S => mult_21_C245_n571);
   mult_21_C245_U354 : ADFULD1 port map( A => mult_21_C245_n582, B => 
                           mult_21_C245_n573, CI => mult_21_C245_n571, CO => 
                           mult_21_C245_n568, S => mult_21_C245_n569);
   mult_21_C245_U353 : ADHALFDL port map( A => mult_21_C245_n1212, B => 
                           mult_21_C245_n947, CO => mult_21_C245_n566, S => 
                           mult_21_C245_n567);
   mult_21_C245_U352 : ADFULD1 port map( A => mult_21_C245_n1104, B => 
                           mult_21_C245_n1044, CI => mult_21_C245_n1182, CO => 
                           mult_21_C245_n564, S => mult_21_C245_n565);
   mult_21_C245_U351 : ADFULD1 port map( A => mult_21_C245_n1154, B => 
                           mult_21_C245_n1082, CI => mult_21_C245_n567, CO => 
                           mult_21_C245_n562, S => mult_21_C245_n563);
   mult_21_C245_U350 : ADFULD1 port map( A => mult_21_C245_n1062, B => 
                           mult_21_C245_n1128, CI => mult_21_C245_n578, CO => 
                           mult_21_C245_n560, S => mult_21_C245_n561);
   mult_21_C245_U349 : ADFULD1 port map( A => mult_21_C245_n574, B => 
                           mult_21_C245_n576, CI => mult_21_C245_n565, CO => 
                           mult_21_C245_n558, S => mult_21_C245_n559);
   mult_21_C245_U348 : ADFULD1 port map( A => mult_21_C245_n561, B => 
                           mult_21_C245_n563, CI => mult_21_C245_n572, CO => 
                           mult_21_C245_n556, S => mult_21_C245_n557);
   mult_21_C245_U347 : ADFULD1 port map( A => mult_21_C245_n570, B => 
                           mult_21_C245_n559, CI => mult_21_C245_n557, CO => 
                           mult_21_C245_n554, S => mult_21_C245_n555);
   mult_21_C245_U346 : ADHALFDL port map( A => mult_21_C245_n566, B => 
                           mult_21_C245_n1211, CO => mult_21_C245_n552, S => 
                           mult_21_C245_n553);
   mult_21_C245_U345 : ADFULD1 port map( A => mult_21_C245_n1043, B => 
                           mult_21_C245_n1103, CI => mult_21_C245_n1061, CO => 
                           mult_21_C245_n550, S => mult_21_C245_n551);
   mult_21_C245_U344 : ADFULD1 port map( A => mult_21_C245_n1181, B => 
                           mult_21_C245_n1081, CI => mult_21_C245_n1127, CO => 
                           mult_21_C245_n548, S => mult_21_C245_n549);
   mult_21_C245_U343 : ADFULD1 port map( A => mult_21_C245_n553, B => 
                           mult_21_C245_n1153, CI => mult_21_C245_n564, CO => 
                           mult_21_C245_n546, S => mult_21_C245_n547);
   mult_21_C245_U342 : ADFULD1 port map( A => mult_21_C245_n560, B => 
                           mult_21_C245_n562, CI => mult_21_C245_n549, CO => 
                           mult_21_C245_n544, S => mult_21_C245_n545);
   mult_21_C245_U341 : ADFULD1 port map( A => mult_21_C245_n547, B => 
                           mult_21_C245_n551, CI => mult_21_C245_n558, CO => 
                           mult_21_C245_n542, S => mult_21_C245_n543);
   mult_21_C245_U340 : ADFULD1 port map( A => mult_21_C245_n556, B => 
                           mult_21_C245_n545, CI => mult_21_C245_n543, CO => 
                           mult_21_C245_n540, S => mult_21_C245_n541);
   mult_21_C245_U339 : ADHALFDL port map( A => mult_21_C245_n1210, B => 
                           mult_21_C245_n946, CO => mult_21_C245_n538, S => 
                           mult_21_C245_n539);
   mult_21_C245_U338 : ADFULD1 port map( A => mult_21_C245_n1102, B => 
                           mult_21_C245_n1026, CI => mult_21_C245_n1180, CO => 
                           mult_21_C245_n536, S => mult_21_C245_n537);
   mult_21_C245_U337 : ADFULD1 port map( A => mult_21_C245_n1042, B => 
                           mult_21_C245_n1060, CI => mult_21_C245_n539, CO => 
                           mult_21_C245_n534, S => mult_21_C245_n535);
   mult_21_C245_U336 : ADFULD1 port map( A => mult_21_C245_n1080, B => 
                           mult_21_C245_n1152, CI => mult_21_C245_n1126, CO => 
                           mult_21_C245_n532, S => mult_21_C245_n533);
   mult_21_C245_U335 : ADFULD1 port map( A => mult_21_C245_n550, B => 
                           mult_21_C245_n552, CI => mult_21_C245_n548, CO => 
                           mult_21_C245_n530, S => mult_21_C245_n531);
   mult_21_C245_U334 : ADFULD1 port map( A => mult_21_C245_n533, B => 
                           mult_21_C245_n537, CI => mult_21_C245_n535, CO => 
                           mult_21_C245_n528, S => mult_21_C245_n529);
   mult_21_C245_U333 : ADFULD1 port map( A => mult_21_C245_n544, B => 
                           mult_21_C245_n546, CI => mult_21_C245_n531, CO => 
                           mult_21_C245_n526, S => mult_21_C245_n527);
   mult_21_C245_U332 : ADFULD1 port map( A => mult_21_C245_n542, B => 
                           mult_21_C245_n529, CI => mult_21_C245_n527, CO => 
                           mult_21_C245_n524, S => mult_21_C245_n525);
   mult_21_C245_U331 : ADHALFDL port map( A => mult_21_C245_n538, B => 
                           mult_21_C245_n1209, CO => mult_21_C245_n522, S => 
                           mult_21_C245_n523);
   mult_21_C245_U330 : ADFULD1 port map( A => mult_21_C245_n1179, B => 
                           mult_21_C245_n1079, CI => mult_21_C245_n1151, CO => 
                           mult_21_C245_n520, S => mult_21_C245_n521);
   mult_21_C245_U329 : ADFULD1 port map( A => mult_21_C245_n1025, B => 
                           mult_21_C245_n1041, CI => mult_21_C245_n1059, CO => 
                           mult_21_C245_n518, S => mult_21_C245_n519);
   mult_21_C245_U328 : ADFULD1 port map( A => mult_21_C245_n1101, B => 
                           mult_21_C245_n1125, CI => mult_21_C245_n523, CO => 
                           mult_21_C245_n516, S => mult_21_C245_n517);
   mult_21_C245_U327 : ADFULD1 port map( A => mult_21_C245_n534, B => 
                           mult_21_C245_n536, CI => mult_21_C245_n532, CO => 
                           mult_21_C245_n514, S => mult_21_C245_n515);
   mult_21_C245_U326 : ADFULD1 port map( A => mult_21_C245_n521, B => 
                           mult_21_C245_n519, CI => mult_21_C245_n517, CO => 
                           mult_21_C245_n512, S => mult_21_C245_n513);
   mult_21_C245_U325 : ADFULD1 port map( A => mult_21_C245_n528, B => 
                           mult_21_C245_n530, CI => mult_21_C245_n515, CO => 
                           mult_21_C245_n510, S => mult_21_C245_n511);
   mult_21_C245_U324 : ADFULD1 port map( A => mult_21_C245_n526, B => 
                           mult_21_C245_n513, CI => mult_21_C245_n511, CO => 
                           mult_21_C245_n508, S => mult_21_C245_n509);
   mult_21_C245_U323 : ADHALFDL port map( A => mult_21_C245_n1208, B => 
                           mult_21_C245_n945, CO => mult_21_C245_n506, S => 
                           mult_21_C245_n507);
   mult_21_C245_U322 : ADFULD1 port map( A => mult_21_C245_n1078, B => 
                           mult_21_C245_n1010, CI => mult_21_C245_n1024, CO => 
                           mult_21_C245_n504, S => mult_21_C245_n505);
   mult_21_C245_U321 : ADFULD1 port map( A => mult_21_C245_n1178, B => 
                           mult_21_C245_n1100, CI => mult_21_C245_n507, CO => 
                           mult_21_C245_n502, S => mult_21_C245_n503);
   mult_21_C245_U320 : ADFULD1 port map( A => mult_21_C245_n1040, B => 
                           mult_21_C245_n1150, CI => mult_21_C245_n1058, CO => 
                           mult_21_C245_n500, S => mult_21_C245_n501);
   mult_21_C245_U319 : ADFULD1 port map( A => mult_21_C245_n522, B => 
                           mult_21_C245_n1124, CI => mult_21_C245_n520, CO => 
                           mult_21_C245_n498, S => mult_21_C245_n499);
   mult_21_C245_U318 : ADFULD1 port map( A => mult_21_C245_n505, B => 
                           mult_21_C245_n518, CI => mult_21_C245_n501, CO => 
                           mult_21_C245_n496, S => mult_21_C245_n497);
   mult_21_C245_U317 : ADFULD1 port map( A => mult_21_C245_n516, B => 
                           mult_21_C245_n503, CI => mult_21_C245_n514, CO => 
                           mult_21_C245_n494, S => mult_21_C245_n495);
   mult_21_C245_U316 : ADFULD1 port map( A => mult_21_C245_n497, B => 
                           mult_21_C245_n499, CI => mult_21_C245_n512, CO => 
                           mult_21_C245_n492, S => mult_21_C245_n493);
   mult_21_C245_U315 : ADFULD1 port map( A => mult_21_C245_n510, B => 
                           mult_21_C245_n495, CI => mult_21_C245_n493, CO => 
                           mult_21_C245_n490, S => mult_21_C245_n491);
   mult_21_C245_U314 : ADHALFDL port map( A => mult_21_C245_n506, B => 
                           mult_21_C245_n1207, CO => mult_21_C245_n488, S => 
                           mult_21_C245_n489);
   mult_21_C245_U313 : ADFULD1 port map( A => mult_21_C245_n1009, B => 
                           mult_21_C245_n1077, CI => mult_21_C245_n1023, CO => 
                           mult_21_C245_n486, S => mult_21_C245_n487);
   mult_21_C245_U312 : ADFULD1 port map( A => mult_21_C245_n1177, B => 
                           mult_21_C245_n1099, CI => mult_21_C245_n1039, CO => 
                           mult_21_C245_n484, S => mult_21_C245_n485);
   mult_21_C245_U311 : ADFULD1 port map( A => mult_21_C245_n1057, B => 
                           mult_21_C245_n1149, CI => mult_21_C245_n1123, CO => 
                           mult_21_C245_n482, S => mult_21_C245_n483);
   mult_21_C245_U310 : ADFULD1 port map( A => mult_21_C245_n504, B => 
                           mult_21_C245_n489, CI => mult_21_C245_n502, CO => 
                           mult_21_C245_n480, S => mult_21_C245_n481);
   mult_21_C245_U309 : ADFULD1 port map( A => mult_21_C245_n483, B => 
                           mult_21_C245_n500, CI => mult_21_C245_n485, CO => 
                           mult_21_C245_n478, S => mult_21_C245_n479);
   mult_21_C245_U308 : ADFULD1 port map( A => mult_21_C245_n498, B => 
                           mult_21_C245_n487, CI => mult_21_C245_n496, CO => 
                           mult_21_C245_n476, S => mult_21_C245_n477);
   mult_21_C245_U307 : ADFULD1 port map( A => mult_21_C245_n479, B => 
                           mult_21_C245_n481, CI => mult_21_C245_n494, CO => 
                           mult_21_C245_n474, S => mult_21_C245_n475);
   mult_21_C245_U306 : ADFULD1 port map( A => mult_21_C245_n492, B => 
                           mult_21_C245_n477, CI => mult_21_C245_n475, CO => 
                           mult_21_C245_n472, S => mult_21_C245_n473);
   mult_21_C245_U305 : ADHALFDL port map( A => mult_21_C245_n1206, B => 
                           mult_21_C245_n944, CO => mult_21_C245_n470, S => 
                           mult_21_C245_n471);
   mult_21_C245_U304 : ADFULD1 port map( A => mult_21_C245_n1076, B => 
                           mult_21_C245_n996, CI => mult_21_C245_n1176, CO => 
                           mult_21_C245_n468, S => mult_21_C245_n469);
   mult_21_C245_U303 : ADFULD1 port map( A => mult_21_C245_n1008, B => 
                           mult_21_C245_n1038, CI => mult_21_C245_n471, CO => 
                           mult_21_C245_n466, S => mult_21_C245_n467);
   mult_21_C245_U302 : ADFULD1 port map( A => mult_21_C245_n1022, B => 
                           mult_21_C245_n1148, CI => mult_21_C245_n1056, CO => 
                           mult_21_C245_n464, S => mult_21_C245_n465);
   mult_21_C245_U301 : ADFULD1 port map( A => mult_21_C245_n1098, B => 
                           mult_21_C245_n1122, CI => mult_21_C245_n488, CO => 
                           mult_21_C245_n462, S => mult_21_C245_n463);
   mult_21_C245_U300 : ADFULD1 port map( A => mult_21_C245_n482, B => 
                           mult_21_C245_n486, CI => mult_21_C245_n484, CO => 
                           mult_21_C245_n460, S => mult_21_C245_n461);
   mult_21_C245_U299 : ADFULD1 port map( A => mult_21_C245_n465, B => 
                           mult_21_C245_n469, CI => mult_21_C245_n467, CO => 
                           mult_21_C245_n458, S => mult_21_C245_n459);
   mult_21_C245_U298 : ADFULD1 port map( A => mult_21_C245_n480, B => 
                           mult_21_C245_n463, CI => mult_21_C245_n478, CO => 
                           mult_21_C245_n456, S => mult_21_C245_n457);
   mult_21_C245_U297 : ADFULD1 port map( A => mult_21_C245_n459, B => 
                           mult_21_C245_n461, CI => mult_21_C245_n476, CO => 
                           mult_21_C245_n454, S => mult_21_C245_n455);
   mult_21_C245_U296 : ADFULD1 port map( A => mult_21_C245_n474, B => 
                           mult_21_C245_n457, CI => mult_21_C245_n455, CO => 
                           mult_21_C245_n452, S => mult_21_C245_n453);
   mult_21_C245_U295 : ADHALFDL port map( A => mult_21_C245_n470, B => 
                           mult_21_C245_n1205, CO => mult_21_C245_n450, S => 
                           mult_21_C245_n451);
   mult_21_C245_U294 : ADFULD1 port map( A => mult_21_C245_n1175, B => 
                           mult_21_C245_n1055, CI => mult_21_C245_n1147, CO => 
                           mult_21_C245_n448, S => mult_21_C245_n449);
   mult_21_C245_U293 : ADFULD1 port map( A => mult_21_C245_n1121, B => 
                           mult_21_C245_n1021, CI => mult_21_C245_n1097, CO => 
                           mult_21_C245_n446, S => mult_21_C245_n447);
   mult_21_C245_U292 : ADFULD1 port map( A => mult_21_C245_n995, B => 
                           mult_21_C245_n1075, CI => mult_21_C245_n1007, CO => 
                           mult_21_C245_n444, S => mult_21_C245_n445);
   mult_21_C245_U291 : ADFULD1 port map( A => mult_21_C245_n451, B => 
                           mult_21_C245_n1037, CI => mult_21_C245_n468, CO => 
                           mult_21_C245_n442, S => mult_21_C245_n443);
   mult_21_C245_U290 : ADFULD1 port map( A => mult_21_C245_n464, B => 
                           mult_21_C245_n466, CI => mult_21_C245_n462, CO => 
                           mult_21_C245_n440, S => mult_21_C245_n441);
   mult_21_C245_U289 : ADFULD1 port map( A => mult_21_C245_n449, B => 
                           mult_21_C245_n445, CI => mult_21_C245_n447, CO => 
                           mult_21_C245_n438, S => mult_21_C245_n439);
   mult_21_C245_U288 : ADFULD1 port map( A => mult_21_C245_n443, B => 
                           mult_21_C245_n460, CI => mult_21_C245_n458, CO => 
                           mult_21_C245_n436, S => mult_21_C245_n437);
   mult_21_C245_U287 : ADFULD1 port map( A => mult_21_C245_n439, B => 
                           mult_21_C245_n441, CI => mult_21_C245_n456, CO => 
                           mult_21_C245_n434, S => mult_21_C245_n435);
   mult_21_C245_U286 : ADFULD1 port map( A => mult_21_C245_n454, B => 
                           mult_21_C245_n437, CI => mult_21_C245_n435, CO => 
                           mult_21_C245_n432, S => mult_21_C245_n433);
   mult_21_C245_U285 : ADHALFDL port map( A => mult_21_C245_n1204, B => 
                           mult_21_C245_n943, CO => mult_21_C245_n430, S => 
                           mult_21_C245_n431);
   mult_21_C245_U284 : ADFULD1 port map( A => mult_21_C245_n1054, B => 
                           mult_21_C245_n984, CI => mult_21_C245_n994, CO => 
                           mult_21_C245_n428, S => mult_21_C245_n429);
   mult_21_C245_U283 : ADFULD1 port map( A => mult_21_C245_n1174, B => 
                           mult_21_C245_n1036, CI => mult_21_C245_n431, CO => 
                           mult_21_C245_n426, S => mult_21_C245_n427);
   mult_21_C245_U282 : ADFULD1 port map( A => mult_21_C245_n1006, B => 
                           mult_21_C245_n1146, CI => mult_21_C245_n1020, CO => 
                           mult_21_C245_n424, S => mult_21_C245_n425);
   mult_21_C245_U281 : ADFULD1 port map( A => mult_21_C245_n1074, B => 
                           mult_21_C245_n1120, CI => mult_21_C245_n1096, CO => 
                           mult_21_C245_n422, S => mult_21_C245_n423);
   mult_21_C245_U280 : ADFULD1 port map( A => mult_21_C245_n448, B => 
                           mult_21_C245_n450, CI => mult_21_C245_n446, CO => 
                           mult_21_C245_n420, S => mult_21_C245_n421);
   mult_21_C245_U279 : ADFULD1 port map( A => mult_21_C245_n429, B => 
                           mult_21_C245_n444, CI => mult_21_C245_n423, CO => 
                           mult_21_C245_n418, S => mult_21_C245_n419);
   mult_21_C245_U278 : ADFULD1 port map( A => mult_21_C245_n427, B => 
                           mult_21_C245_n425, CI => mult_21_C245_n442, CO => 
                           mult_21_C245_n416, S => mult_21_C245_n417);
   mult_21_C245_U277 : ADFULD1 port map( A => mult_21_C245_n421, B => 
                           mult_21_C245_n440, CI => mult_21_C245_n438, CO => 
                           mult_21_C245_n414, S => mult_21_C245_n415);
   mult_21_C245_U276 : ADFULD1 port map( A => mult_21_C245_n417, B => 
                           mult_21_C245_n419, CI => mult_21_C245_n436, CO => 
                           mult_21_C245_n412, S => mult_21_C245_n413);
   mult_21_C245_U275 : ADFULD1 port map( A => mult_21_C245_n434, B => 
                           mult_21_C245_n415, CI => mult_21_C245_n413, CO => 
                           mult_21_C245_n410, S => mult_21_C245_n411);
   mult_21_C245_U274 : ADHALFDL port map( A => mult_21_C245_n430, B => 
                           mult_21_C245_n1203, CO => mult_21_C245_n408, S => 
                           mult_21_C245_n409);
   mult_21_C245_U273 : ADFULD1 port map( A => mult_21_C245_n983, B => 
                           mult_21_C245_n1053, CI => mult_21_C245_n993, CO => 
                           mult_21_C245_n406, S => mult_21_C245_n407);
   mult_21_C245_U272 : ADFULD1 port map( A => mult_21_C245_n1173, B => 
                           mult_21_C245_n1035, CI => mult_21_C245_n1145, CO => 
                           mult_21_C245_n404, S => mult_21_C245_n405);
   mult_21_C245_U271 : ADFULD1 port map( A => mult_21_C245_n1005, B => 
                           mult_21_C245_n1119, CI => mult_21_C245_n1019, CO => 
                           mult_21_C245_n402, S => mult_21_C245_n403);
   mult_21_C245_U270 : ADFULD1 port map( A => mult_21_C245_n1073, B => 
                           mult_21_C245_n1095, CI => mult_21_C245_n409, CO => 
                           mult_21_C245_n400, S => mult_21_C245_n401);
   mult_21_C245_U269 : ADFULD1 port map( A => mult_21_C245_n426, B => 
                           mult_21_C245_n428, CI => mult_21_C245_n422, CO => 
                           mult_21_C245_n398, S => mult_21_C245_n399);
   mult_21_C245_U268 : ADFULD1 port map( A => mult_21_C245_n403, B => 
                           mult_21_C245_n424, CI => mult_21_C245_n405, CO => 
                           mult_21_C245_n396, S => mult_21_C245_n397);
   mult_21_C245_U267 : ADFULD1 port map( A => mult_21_C245_n401, B => 
                           mult_21_C245_n407, CI => mult_21_C245_n420, CO => 
                           mult_21_C245_n394, S => mult_21_C245_n395);
   mult_21_C245_U266 : ADFULD1 port map( A => mult_21_C245_n399, B => 
                           mult_21_C245_n418, CI => mult_21_C245_n416, CO => 
                           mult_21_C245_n392, S => mult_21_C245_n393);
   mult_21_C245_U265 : ADFULD1 port map( A => mult_21_C245_n395, B => 
                           mult_21_C245_n397, CI => mult_21_C245_n414, CO => 
                           mult_21_C245_n390, S => mult_21_C245_n391);
   mult_21_C245_U264 : ADFULD1 port map( A => mult_21_C245_n412, B => 
                           mult_21_C245_n393, CI => mult_21_C245_n391, CO => 
                           mult_21_C245_n388, S => mult_21_C245_n389);
   mult_21_C245_U263 : ADHALFDL port map( A => mult_21_C245_n1202, B => 
                           mult_21_C245_n942, CO => mult_21_C245_n386, S => 
                           mult_21_C245_n387);
   mult_21_C245_U262 : ADFULD1 port map( A => mult_21_C245_n1052, B => 
                           mult_21_C245_n974, CI => mult_21_C245_n1172, CO => 
                           mult_21_C245_n384, S => mult_21_C245_n385);
   mult_21_C245_U261 : ADFULD1 port map( A => mult_21_C245_n982, B => 
                           mult_21_C245_n1018, CI => mult_21_C245_n387, CO => 
                           mult_21_C245_n382, S => mult_21_C245_n383);
   mult_21_C245_U260 : ADFULD1 port map( A => mult_21_C245_n992, B => 
                           mult_21_C245_n1144, CI => mult_21_C245_n1118, CO => 
                           mult_21_C245_n380, S => mult_21_C245_n381);
   mult_21_C245_U259 : ADFULD1 port map( A => mult_21_C245_n1004, B => 
                           mult_21_C245_n1094, CI => mult_21_C245_n1034, CO => 
                           mult_21_C245_n378, S => mult_21_C245_n379);
   mult_21_C245_U258 : ADFULD1 port map( A => mult_21_C245_n408, B => 
                           mult_21_C245_n1072, CI => mult_21_C245_n406, CO => 
                           mult_21_C245_n376, S => mult_21_C245_n377);
   mult_21_C245_U257 : ADFULD1 port map( A => mult_21_C245_n402, B => 
                           mult_21_C245_n404, CI => mult_21_C245_n385, CO => 
                           mult_21_C245_n374, S => mult_21_C245_n375);
   mult_21_C245_U256 : ADFULD1 port map( A => mult_21_C245_n383, B => 
                           mult_21_C245_n379, CI => mult_21_C245_n381, CO => 
                           mult_21_C245_n372, S => mult_21_C245_n373);
   mult_21_C245_U255 : ADFULD1 port map( A => mult_21_C245_n398, B => 
                           mult_21_C245_n400, CI => mult_21_C245_n377, CO => 
                           mult_21_C245_n370, S => mult_21_C245_n371);
   mult_21_C245_U254 : ADFULD1 port map( A => mult_21_C245_n375, B => 
                           mult_21_C245_n396, CI => mult_21_C245_n373, CO => 
                           mult_21_C245_n368, S => mult_21_C245_n369);
   mult_21_C245_U253 : ADFULD1 port map( A => mult_21_C245_n371, B => 
                           mult_21_C245_n394, CI => mult_21_C245_n392, CO => 
                           mult_21_C245_n366, S => mult_21_C245_n367);
   mult_21_C245_U252 : ADFULD1 port map( A => mult_21_C245_n390, B => 
                           mult_21_C245_n369, CI => mult_21_C245_n367, CO => 
                           mult_21_C245_n364, S => mult_21_C245_n365);
   mult_21_C245_U251 : ADHALFDL port map( A => mult_21_C245_n386, B => 
                           mult_21_C245_n1201, CO => mult_21_C245_n362, S => 
                           mult_21_C245_n363);
   mult_21_C245_U250 : ADFULD1 port map( A => mult_21_C245_n1171, B => 
                           mult_21_C245_n1051, CI => mult_21_C245_n1143, CO => 
                           mult_21_C245_n360, S => mult_21_C245_n361);
   mult_21_C245_U249 : ADFULD1 port map( A => mult_21_C245_n973, B => 
                           mult_21_C245_n1003, CI => mult_21_C245_n981, CO => 
                           mult_21_C245_n358, S => mult_21_C245_n359);
   mult_21_C245_U248 : ADFULD1 port map( A => mult_21_C245_n991, B => 
                           mult_21_C245_n1117, CI => mult_21_C245_n1017, CO => 
                           mult_21_C245_n356, S => mult_21_C245_n357);
   mult_21_C245_U247 : ADFULD1 port map( A => mult_21_C245_n1033, B => 
                           mult_21_C245_n1093, CI => mult_21_C245_n1071, CO => 
                           mult_21_C245_n354, S => mult_21_C245_n355);
   mult_21_C245_U246 : ADFULD1 port map( A => mult_21_C245_n384, B => 
                           mult_21_C245_n363, CI => mult_21_C245_n382, CO => 
                           mult_21_C245_n352, S => mult_21_C245_n353);
   mult_21_C245_U245 : ADFULD1 port map( A => mult_21_C245_n378, B => 
                           mult_21_C245_n380, CI => mult_21_C245_n355, CO => 
                           mult_21_C245_n350, S => mult_21_C245_n351);
   mult_21_C245_U244 : ADFULD1 port map( A => mult_21_C245_n361, B => 
                           mult_21_C245_n357, CI => mult_21_C245_n359, CO => 
                           mult_21_C245_n348, S => mult_21_C245_n349);
   mult_21_C245_U243 : ADFULD1 port map( A => mult_21_C245_n374, B => 
                           mult_21_C245_n376, CI => mult_21_C245_n353, CO => 
                           mult_21_C245_n346, S => mult_21_C245_n347);
   mult_21_C245_U242 : ADFULD1 port map( A => mult_21_C245_n351, B => 
                           mult_21_C245_n372, CI => mult_21_C245_n349, CO => 
                           mult_21_C245_n344, S => mult_21_C245_n345);
   mult_21_C245_U241 : ADFULD1 port map( A => mult_21_C245_n347, B => 
                           mult_21_C245_n370, CI => mult_21_C245_n368, CO => 
                           mult_21_C245_n342, S => mult_21_C245_n343);
   mult_21_C245_U240 : ADFULD1 port map( A => mult_21_C245_n366, B => 
                           mult_21_C245_n345, CI => mult_21_C245_n343, CO => 
                           mult_21_C245_n340, S => mult_21_C245_n341);
   mult_21_C245_U239 : ADHALFDL port map( A => mult_21_C245_n1200, B => 
                           mult_21_C245_n941, CO => mult_21_C245_n338, S => 
                           mult_21_C245_n339);
   mult_21_C245_U238 : ADFULD1 port map( A => mult_21_C245_n1050, B => 
                           mult_21_C245_n966, CI => mult_21_C245_n972, CO => 
                           mult_21_C245_n336, S => mult_21_C245_n337);
   mult_21_C245_U237 : ADFULD1 port map( A => mult_21_C245_n980, B => 
                           mult_21_C245_n1032, CI => mult_21_C245_n339, CO => 
                           mult_21_C245_n334, S => mult_21_C245_n335);
   mult_21_C245_U236 : ADFULD1 port map( A => mult_21_C245_n990, B => 
                           mult_21_C245_n1170, CI => mult_21_C245_n1002, CO => 
                           mult_21_C245_n332, S => mult_21_C245_n333);
   mult_21_C245_U235 : ADFULD1 port map( A => mult_21_C245_n1016, B => 
                           mult_21_C245_n1142, CI => mult_21_C245_n1070, CO => 
                           mult_21_C245_n330, S => mult_21_C245_n331);
   mult_21_C245_U234 : ADFULD1 port map( A => mult_21_C245_n1092, B => 
                           mult_21_C245_n1116, CI => mult_21_C245_n362, CO => 
                           mult_21_C245_n328, S => mult_21_C245_n329);
   mult_21_C245_U233 : ADFULD1 port map( A => mult_21_C245_n354, B => 
                           mult_21_C245_n360, CI => mult_21_C245_n356, CO => 
                           mult_21_C245_n326, S => mult_21_C245_n327);
   mult_21_C245_U232 : ADFULD1 port map( A => mult_21_C245_n337, B => 
                           mult_21_C245_n358, CI => mult_21_C245_n331, CO => 
                           mult_21_C245_n324, S => mult_21_C245_n325);
   mult_21_C245_U231 : ADFULD1 port map( A => mult_21_C245_n333, B => 
                           mult_21_C245_n335, CI => mult_21_C245_n329, CO => 
                           mult_21_C245_n322, S => mult_21_C245_n323);
   mult_21_C245_U230 : ADFULD1 port map( A => mult_21_C245_n350, B => 
                           mult_21_C245_n352, CI => mult_21_C245_n348, CO => 
                           mult_21_C245_n320, S => mult_21_C245_n321);
   mult_21_C245_U229 : ADFULD1 port map( A => mult_21_C245_n325, B => 
                           mult_21_C245_n327, CI => mult_21_C245_n323, CO => 
                           mult_21_C245_n318, S => mult_21_C245_n319);
   mult_21_C245_U228 : ADFULD1 port map( A => mult_21_C245_n344, B => 
                           mult_21_C245_n346, CI => mult_21_C245_n321, CO => 
                           mult_21_C245_n316, S => mult_21_C245_n317);
   mult_21_C245_U227 : ADFULD1 port map( A => mult_21_C245_n342, B => 
                           mult_21_C245_n319, CI => mult_21_C245_n317, CO => 
                           mult_21_C245_n314, S => mult_21_C245_n315);
   mult_21_C245_U226 : ADHALFDL port map( A => mult_21_C245_n338, B => 
                           mult_21_C245_n1199, CO => mult_21_C245_n312, S => 
                           mult_21_C245_n313);
   mult_21_C245_U225 : ADFULD1 port map( A => mult_21_C245_n965, B => 
                           mult_21_C245_n1031, CI => mult_21_C245_n971, CO => 
                           mult_21_C245_n310, S => mult_21_C245_n311);
   mult_21_C245_U224 : ADFULD1 port map( A => mult_21_C245_n979, B => 
                           mult_21_C245_n1049, CI => mult_21_C245_n1169, CO => 
                           mult_21_C245_n308, S => mult_21_C245_n309);
   mult_21_C245_U223 : ADFULD1 port map( A => mult_21_C245_n1141, B => 
                           mult_21_C245_n1001, CI => mult_21_C245_n989, CO => 
                           mult_21_C245_n306, S => mult_21_C245_n307);
   mult_21_C245_U222 : ADFULD1 port map( A => mult_21_C245_n1015, B => 
                           mult_21_C245_n1115, CI => mult_21_C245_n1069, CO => 
                           mult_21_C245_n304, S => mult_21_C245_n305);
   mult_21_C245_U221 : ADFULD1 port map( A => mult_21_C245_n313, B => 
                           mult_21_C245_n1091, CI => mult_21_C245_n336, CO => 
                           mult_21_C245_n302, S => mult_21_C245_n303);
   mult_21_C245_U220 : ADFULD1 port map( A => mult_21_C245_n332, B => 
                           mult_21_C245_n330, CI => mult_21_C245_n334, CO => 
                           mult_21_C245_n300, S => mult_21_C245_n301);
   mult_21_C245_U219 : ADFULD1 port map( A => mult_21_C245_n305, B => 
                           mult_21_C245_n328, CI => mult_21_C245_n311, CO => 
                           mult_21_C245_n298, S => mult_21_C245_n299);
   mult_21_C245_U218 : ADFULD1 port map( A => mult_21_C245_n307, B => 
                           mult_21_C245_n309, CI => mult_21_C245_n326, CO => 
                           mult_21_C245_n296, S => mult_21_C245_n297);
   mult_21_C245_U217 : ADFULD1 port map( A => mult_21_C245_n324, B => 
                           mult_21_C245_n303, CI => mult_21_C245_n301, CO => 
                           mult_21_C245_n294, S => mult_21_C245_n295);
   mult_21_C245_U216 : ADFULD1 port map( A => mult_21_C245_n299, B => 
                           mult_21_C245_n322, CI => mult_21_C245_n320, CO => 
                           mult_21_C245_n292, S => mult_21_C245_n293);
   mult_21_C245_U215 : ADFULD1 port map( A => mult_21_C245_n318, B => 
                           mult_21_C245_n297, CI => mult_21_C245_n295, CO => 
                           mult_21_C245_n290, S => mult_21_C245_n291);
   mult_21_C245_U214 : ADFULD1 port map( A => mult_21_C245_n316, B => 
                           mult_21_C245_n293, CI => mult_21_C245_n291, CO => 
                           mult_21_C245_n288, S => mult_21_C245_n289);
   mult_21_C245_U213 : ADHALFDL port map( A => mult_21_C245_n1198, B => 
                           mult_21_C245_n940, CO => mult_21_C245_n286, S => 
                           mult_21_C245_n287);
   mult_21_C245_U212 : ADFULD1 port map( A => mult_21_C245_n1030, B => 
                           mult_21_C245_n960, CI => mult_21_C245_n1168, CO => 
                           mult_21_C245_n284, S => mult_21_C245_n285);
   mult_21_C245_U211 : ADFULD1 port map( A => mult_21_C245_n1140, B => 
                           mult_21_C245_n1000, CI => mult_21_C245_n287, CO => 
                           mult_21_C245_n282, S => mult_21_C245_n283);
   mult_21_C245_U210 : ADFULD1 port map( A => mult_21_C245_n964, B => 
                           mult_21_C245_n1114, CI => mult_21_C245_n970, CO => 
                           mult_21_C245_n280, S => mult_21_C245_n281);
   mult_21_C245_U209 : ADFULD1 port map( A => mult_21_C245_n978, B => 
                           mult_21_C245_n1090, CI => mult_21_C245_n988, CO => 
                           mult_21_C245_n278, S => mult_21_C245_n279);
   mult_21_C245_U208 : ADFULD1 port map( A => mult_21_C245_n1014, B => 
                           mult_21_C245_n1068, CI => mult_21_C245_n1048, CO => 
                           mult_21_C245_n276, S => mult_21_C245_n277);
   mult_21_C245_U207 : ADFULD1 port map( A => mult_21_C245_n304, B => 
                           mult_21_C245_n312, CI => mult_21_C245_n306, CO => 
                           mult_21_C245_n274, S => mult_21_C245_n275);
   mult_21_C245_U206 : ADFULD1 port map( A => mult_21_C245_n310, B => 
                           mult_21_C245_n308, CI => mult_21_C245_n285, CO => 
                           mult_21_C245_n272, S => mult_21_C245_n273);
   mult_21_C245_U205 : ADFULD1 port map( A => mult_21_C245_n283, B => 
                           mult_21_C245_n277, CI => mult_21_C245_n279, CO => 
                           mult_21_C245_n270, S => mult_21_C245_n271);
   mult_21_C245_U204 : ADFULD1 port map( A => mult_21_C245_n302, B => 
                           mult_21_C245_n281, CI => mult_21_C245_n300, CO => 
                           mult_21_C245_n268, S => mult_21_C245_n269);
   mult_21_C245_U203 : ADFULD1 port map( A => mult_21_C245_n275, B => 
                           mult_21_C245_n298, CI => mult_21_C245_n273, CO => 
                           mult_21_C245_n266, S => mult_21_C245_n267);
   mult_21_C245_U202 : ADFULD1 port map( A => mult_21_C245_n296, B => 
                           mult_21_C245_n271, CI => mult_21_C245_n269, CO => 
                           mult_21_C245_n264, S => mult_21_C245_n265);
   mult_21_C245_U201 : ADFULD1 port map( A => mult_21_C245_n267, B => 
                           mult_21_C245_n294, CI => mult_21_C245_n292, CO => 
                           mult_21_C245_n262, S => mult_21_C245_n263);
   mult_21_C245_U200 : ADFULD1 port map( A => mult_21_C245_n290, B => 
                           mult_21_C245_n265, CI => mult_21_C245_n263, CO => 
                           mult_21_C245_n260, S => mult_21_C245_n261);
   mult_21_C245_U199 : ADHALFDL port map( A => mult_21_C245_n286, B => 
                           mult_21_C245_n1197, CO => mult_21_C245_n258, S => 
                           mult_21_C245_n259);
   mult_21_C245_U198 : ADFULD1 port map( A => mult_21_C245_n1167, B => 
                           mult_21_C245_n1029, CI => mult_21_C245_n1139, CO => 
                           mult_21_C245_n256, S => mult_21_C245_n257);
   mult_21_C245_U197 : ADFULD1 port map( A => mult_21_C245_n1113, B => 
                           mult_21_C245_n987, CI => mult_21_C245_n1089, CO => 
                           mult_21_C245_n254, S => mult_21_C245_n255);
   mult_21_C245_U196 : ADFULD1 port map( A => mult_21_C245_n959, B => 
                           mult_21_C245_n969, CI => mult_21_C245_n963, CO => 
                           mult_21_C245_n252, S => mult_21_C245_n253);
   mult_21_C245_U195 : ADFULD1 port map( A => mult_21_C245_n977, B => 
                           mult_21_C245_n1067, CI => mult_21_C245_n999, CO => 
                           mult_21_C245_n250, S => mult_21_C245_n251);
   mult_21_C245_U194 : ADFULD1 port map( A => mult_21_C245_n1047, B => 
                           mult_21_C245_n1013, CI => mult_21_C245_n259, CO => 
                           mult_21_C245_n248, S => mult_21_C245_n249);
   mult_21_C245_U193 : ADFULD1 port map( A => mult_21_C245_n278, B => 
                           mult_21_C245_n284, CI => mult_21_C245_n282, CO => 
                           mult_21_C245_n246, S => mult_21_C245_n247);
   mult_21_C245_U192 : ADFULD1 port map( A => mult_21_C245_n280, B => 
                           mult_21_C245_n276, CI => mult_21_C245_n251, CO => 
                           mult_21_C245_n244, S => mult_21_C245_n245);
   mult_21_C245_U191 : ADFULD1 port map( A => mult_21_C245_n253, B => 
                           mult_21_C245_n255, CI => mult_21_C245_n257, CO => 
                           mult_21_C245_n242, S => mult_21_C245_n243);
   mult_21_C245_U190 : ADFULD1 port map( A => mult_21_C245_n274, B => 
                           mult_21_C245_n249, CI => mult_21_C245_n272, CO => 
                           mult_21_C245_n240, S => mult_21_C245_n241);
   mult_21_C245_U189 : ADFULD1 port map( A => mult_21_C245_n270, B => 
                           mult_21_C245_n247, CI => mult_21_C245_n245, CO => 
                           mult_21_C245_n238, S => mult_21_C245_n239);
   mult_21_C245_U188 : ADFULD1 port map( A => mult_21_C245_n268, B => 
                           mult_21_C245_n243, CI => mult_21_C245_n241, CO => 
                           mult_21_C245_n236, S => mult_21_C245_n237);
   mult_21_C245_U187 : ADFULD1 port map( A => mult_21_C245_n239, B => 
                           mult_21_C245_n266, CI => mult_21_C245_n264, CO => 
                           mult_21_C245_n234, S => mult_21_C245_n235);
   mult_21_C245_U186 : ADFULD1 port map( A => mult_21_C245_n262, B => 
                           mult_21_C245_n237, CI => mult_21_C245_n235, CO => 
                           mult_21_C245_n232, S => mult_21_C245_n233);
   mult_21_C245_U185 : ADHALFDL port map( A => mult_21_C245_n1196, B => 
                           mult_21_C245_n939, CO => mult_21_C245_n230, S => 
                           mult_21_C245_n231);
   mult_21_C245_U184 : ADFULD1 port map( A => mult_21_C245_n1028, B => 
                           mult_21_C245_n956, CI => mult_21_C245_n958, CO => 
                           mult_21_C245_n228, S => mult_21_C245_n229);
   mult_21_C245_U183 : ADFULD1 port map( A => mult_21_C245_n1166, B => 
                           mult_21_C245_n1012, CI => mult_21_C245_n231, CO => 
                           mult_21_C245_n226, S => mult_21_C245_n227);
   mult_21_C245_U182 : ADFULD1 port map( A => mult_21_C245_n962, B => 
                           mult_21_C245_n1138, CI => mult_21_C245_n968, CO => 
                           mult_21_C245_n224, S => mult_21_C245_n225);
   mult_21_C245_U181 : ADFULD1 port map( A => mult_21_C245_n986, B => 
                           mult_21_C245_n976, CI => mult_21_C245_n998, CO => 
                           mult_21_C245_n222, S => mult_21_C245_n223);
   mult_21_C245_U180 : ADFULD1 port map( A => mult_21_C245_n1046, B => 
                           mult_21_C245_n1112, CI => mult_21_C245_n1066, CO => 
                           mult_21_C245_n220, S => mult_21_C245_n221);
   mult_21_C245_U179 : ADFULD1 port map( A => mult_21_C245_n258, B => 
                           mult_21_C245_n1088, CI => mult_21_C245_n250, CO => 
                           mult_21_C245_n218, S => mult_21_C245_n219);
   mult_21_C245_U178 : ADFULD1 port map( A => mult_21_C245_n256, B => 
                           mult_21_C245_n252, CI => mult_21_C245_n254, CO => 
                           mult_21_C245_n216, S => mult_21_C245_n217);
   mult_21_C245_U177 : ADFULD1 port map( A => mult_21_C245_n221, B => 
                           mult_21_C245_n229, CI => mult_21_C245_n227, CO => 
                           mult_21_C245_n214, S => mult_21_C245_n215);
   mult_21_C245_U176 : ADFULD1 port map( A => mult_21_C245_n225, B => 
                           mult_21_C245_n223, CI => mult_21_C245_n248, CO => 
                           mult_21_C245_n212, S => mult_21_C245_n213);
   mult_21_C245_U175 : ADFULD1 port map( A => mult_21_C245_n244, B => 
                           mult_21_C245_n246, CI => mult_21_C245_n219, CO => 
                           mult_21_C245_n210, S => mult_21_C245_n211);
   mult_21_C245_U174 : ADFULD1 port map( A => mult_21_C245_n217, B => 
                           mult_21_C245_n242, CI => mult_21_C245_n215, CO => 
                           mult_21_C245_n208, S => mult_21_C245_n209);
   mult_21_C245_U173 : ADFULD1 port map( A => mult_21_C245_n240, B => 
                           mult_21_C245_n213, CI => mult_21_C245_n238, CO => 
                           mult_21_C245_n206, S => mult_21_C245_n207);
   mult_21_C245_U172 : ADFULD1 port map( A => mult_21_C245_n209, B => 
                           mult_21_C245_n211, CI => mult_21_C245_n236, CO => 
                           mult_21_C245_n204, S => mult_21_C245_n205);
   mult_21_C245_U171 : ADFULD1 port map( A => mult_21_C245_n234, B => 
                           mult_21_C245_n207, CI => mult_21_C245_n205, CO => 
                           mult_21_C245_n202, S => mult_21_C245_n203);
   mult_21_C245_U155 : ADHALFDL port map( A => mult_21_C245_n1226, B => N2978, 
                           CO => mult_21_C245_n186, S => N3297);
   mult_21_C245_U154 : ADHALFDL port map( A => mult_21_C245_n186, B => 
                           mult_21_C245_n1225, CO => mult_21_C245_n185, S => 
                           N3298);
   mult_21_C245_U153 : ADFULD1 port map( A => mult_21_C245_n651, B => 
                           mult_21_C245_n1194, CI => mult_21_C245_n185, CO => 
                           mult_21_C245_n184, S => N3299);
   mult_21_C245_U152 : ADFULD1 port map( A => mult_21_C245_n649, B => 
                           mult_21_C245_n1193, CI => mult_21_C245_n184, CO => 
                           mult_21_C245_n183, S => N3300);
   mult_21_C245_U151 : ADFULD1 port map( A => mult_21_C245_n645, B => 
                           mult_21_C245_n648, CI => mult_21_C245_n183, CO => 
                           mult_21_C245_n182, S => N3301);
   mult_21_C245_U150 : ADFULD1 port map( A => mult_21_C245_n641, B => 
                           mult_21_C245_n644, CI => mult_21_C245_n182, CO => 
                           mult_21_C245_n181, S => N3302);
   mult_21_C245_U149 : ADFULD1 port map( A => mult_21_C245_n635, B => 
                           mult_21_C245_n640, CI => mult_21_C245_n181, CO => 
                           mult_21_C245_n180, S => N3303);
   mult_21_C245_U148 : ADFULD1 port map( A => mult_21_C245_n629, B => 
                           mult_21_C245_n634, CI => mult_21_C245_n180, CO => 
                           mult_21_C245_n179, S => N3304);
   mult_21_C245_U147 : ADFULD1 port map( A => mult_21_C245_n621, B => 
                           mult_21_C245_n628, CI => mult_21_C245_n179, CO => 
                           mult_21_C245_n178, S => N3305);
   mult_21_C245_U146 : ADFULD1 port map( A => mult_21_C245_n613, B => 
                           mult_21_C245_n620, CI => mult_21_C245_n178, CO => 
                           mult_21_C245_n177, S => N3306);
   mult_21_C245_U145 : ADFULD1 port map( A => mult_21_C245_n603, B => 
                           mult_21_C245_n612, CI => mult_21_C245_n177, CO => 
                           mult_21_C245_n176, S => N3307);
   mult_21_C245_U144 : ADFULD1 port map( A => mult_21_C245_n593, B => 
                           mult_21_C245_n602, CI => mult_21_C245_n176, CO => 
                           mult_21_C245_n175, S => N3308);
   mult_21_C245_U143 : ADFULD1 port map( A => mult_21_C245_n581, B => 
                           mult_21_C245_n592, CI => mult_21_C245_n175, CO => 
                           mult_21_C245_n174, S => N3309);
   mult_21_C245_U142 : ADFULD1 port map( A => mult_21_C245_n569, B => 
                           mult_21_C245_n580, CI => mult_21_C245_n174, CO => 
                           mult_21_C245_n173, S => N3310);
   mult_21_C245_U141 : ADFULD1 port map( A => mult_21_C245_n555, B => 
                           mult_21_C245_n568, CI => mult_21_C245_n173, CO => 
                           mult_21_C245_n172, S => N3311);
   mult_21_C245_U140 : ADFULD1 port map( A => mult_21_C245_n541, B => 
                           mult_21_C245_n554, CI => mult_21_C245_n172, CO => 
                           mult_21_C245_n171, S => N3312);
   mult_21_C245_U139 : ADFULD1 port map( A => mult_21_C245_n525, B => 
                           mult_21_C245_n540, CI => mult_21_C245_n171, CO => 
                           mult_21_C245_n170, S => N3313);
   mult_21_C245_U138 : ADFULD1 port map( A => mult_21_C245_n509, B => 
                           mult_21_C245_n524, CI => mult_21_C245_n170, CO => 
                           mult_21_C245_n169, S => N3314);
   mult_21_C245_U137 : ADFULD1 port map( A => mult_21_C245_n491, B => 
                           mult_21_C245_n508, CI => mult_21_C245_n169, CO => 
                           mult_21_C245_n168, S => N3315);
   mult_21_C245_U136 : ADFULD1 port map( A => mult_21_C245_n473, B => 
                           mult_21_C245_n490, CI => mult_21_C245_n168, CO => 
                           mult_21_C245_n167, S => N3316);
   mult_21_C245_U135 : ADFULD1 port map( A => mult_21_C245_n453, B => 
                           mult_21_C245_n472, CI => mult_21_C245_n167, CO => 
                           mult_21_C245_n166, S => N3317);
   mult_21_C245_U134 : ADFULD1 port map( A => mult_21_C245_n433, B => 
                           mult_21_C245_n452, CI => mult_21_C245_n166, CO => 
                           mult_21_C245_n165, S => N3318);
   mult_21_C245_U133 : ADFULD1 port map( A => mult_21_C245_n411, B => 
                           mult_21_C245_n432, CI => mult_21_C245_n165, CO => 
                           mult_21_C245_n164, S => N3319);
   mult_21_C245_U132 : ADFULD1 port map( A => mult_21_C245_n389, B => 
                           mult_21_C245_n410, CI => mult_21_C245_n164, CO => 
                           mult_21_C245_n163, S => N3320);
   mult_21_C245_U131 : ADFULD1 port map( A => mult_21_C245_n365, B => 
                           mult_21_C245_n388, CI => mult_21_C245_n163, CO => 
                           mult_21_C245_n162, S => N3321);
   mult_21_C245_U130 : ADFULD1 port map( A => mult_21_C245_n341, B => 
                           mult_21_C245_n364, CI => mult_21_C245_n162, CO => 
                           mult_21_C245_n161, S => N3322);
   mult_21_C245_U129 : ADFULD1 port map( A => mult_21_C245_n315, B => 
                           mult_21_C245_n340, CI => mult_21_C245_n161, CO => 
                           mult_21_C245_n160, S => N3323);
   mult_21_C245_U128 : ADFULD1 port map( A => mult_21_C245_n289, B => 
                           mult_21_C245_n314, CI => mult_21_C245_n160, CO => 
                           mult_21_C245_n159, S => N3324);
   mult_21_C245_U127 : ADFULD1 port map( A => mult_21_C245_n261, B => 
                           mult_21_C245_n288, CI => mult_21_C245_n159, CO => 
                           mult_21_C245_n158, S => N3325);
   mult_21_C245_U126 : ADFULD1 port map( A => mult_21_C245_n233, B => 
                           mult_21_C245_n260, CI => mult_21_C245_n158, CO => 
                           mult_21_C245_n157, S => N3326);
   mult_21_C245_U125 : ADFULD1 port map( A => mult_21_C245_n203, B => 
                           mult_21_C245_n232, CI => mult_21_C245_n157, CO => 
                           mult_21_C245_n156, S => N3327);
   mult_21_C247_U1402 : AOI21D1 port map( A1 => N3036, A2 => N3037, B => 
                           mult_21_C247_n1427, Z => mult_21_C247_n940);
   mult_21_C247_U1401 : OAI21D1 port map( A1 => N3039, A2 => N3038, B => 
                           mult_21_C247_n1428, Z => mult_21_C247_n104);
   mult_21_C247_U1400 : AOI21D1 port map( A1 => N3038, A2 => N3039, B => 
                           mult_21_C247_n1428, Z => mult_21_C247_n939);
   mult_21_C247_U1399 : AOI21D1 port map( A1 => N3010, A2 => N3011, B => 
                           mult_21_C247_n1401, Z => mult_21_C247_n953);
   mult_21_C247_U1398 : AOI21D1 port map( A1 => N3012, A2 => N3013, B => 
                           mult_21_C247_n1403, Z => mult_21_C247_n952);
   mult_21_C247_U1397 : AOI21D1 port map( A1 => N3014, A2 => N3015, B => 
                           mult_21_C247_n1405, Z => mult_21_C247_n951);
   mult_21_C247_U1396 : AOI21D1 port map( A1 => N3016, A2 => N3017, B => 
                           mult_21_C247_n1407, Z => mult_21_C247_n950);
   mult_21_C247_U1395 : AOI21D1 port map( A1 => N3018, A2 => N3019, B => 
                           mult_21_C247_n1409, Z => mult_21_C247_n949);
   mult_21_C247_U1394 : AOI21D1 port map( A1 => N3020, A2 => N3021, B => 
                           mult_21_C247_n1411, Z => mult_21_C247_n948);
   mult_21_C247_U1393 : AOI21D1 port map( A1 => N3022, A2 => N3023, B => 
                           mult_21_C247_n1413, Z => mult_21_C247_n947);
   mult_21_C247_U1392 : EXOR2D1 port map( A1 => N3039, A2 => N3038, Z => 
                           mult_21_C247_n1457);
   mult_21_C247_U1391 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C247_n1457, Z => mult_21_C247_n652);
   mult_21_C247_U1390 : NAN2D1 port map( A1 => N3201, A2 => mult_21_C247_n1457,
                           Z => mult_21_C247_n653);
   mult_21_C247_U1389 : EXOR2D1 port map( A1 => N3037, A2 => N3036, Z => 
                           mult_21_C247_n1456);
   mult_21_C247_U1388 : MUXB2DL port map( A0 => N3203, A1 => mult_21_C247_n1390
                           , SL => mult_21_C247_n1456, Z => mult_21_C247_n654);
   mult_21_C247_U1387 : MUXB2DL port map( A0 => mult_21_C247_n1394, A1 => 
                           mult_21_C247_n1392, SL => mult_21_C247_n1456, Z => 
                           mult_21_C247_n655);
   mult_21_C247_U1386 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C247_n1456, Z => mult_21_C247_n656);
   mult_21_C247_U1385 : NAN2D1 port map( A1 => N3201, A2 => mult_21_C247_n1456,
                           Z => mult_21_C247_n657);
   mult_21_C247_U1384 : EXOR2D1 port map( A1 => N3035, A2 => N3034, Z => 
                           mult_21_C247_n1455);
   mult_21_C247_U1383 : MUXB2DL port map( A0 => mult_21_C247_n1387, A1 => 
                           mult_21_C247_n1385, SL => mult_21_C247_n1455, Z => 
                           mult_21_C247_n658);
   mult_21_C247_U1382 : MUXB2DL port map( A0 => mult_21_C247_n1389, A1 => N3205
                           , SL => mult_21_C247_n1455, Z => mult_21_C247_n659);
   mult_21_C247_U1381 : MUXB2DL port map( A0 => N3203, A1 => mult_21_C247_n1390
                           , SL => mult_21_C247_n1455, Z => mult_21_C247_n660);
   mult_21_C247_U1380 : MUXB2DL port map( A0 => mult_21_C247_n1394, A1 => N3203
                           , SL => mult_21_C247_n1455, Z => mult_21_C247_n661);
   mult_21_C247_U1379 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C247_n1455, Z => mult_21_C247_n662);
   mult_21_C247_U1378 : NAN2D1 port map( A1 => N3201, A2 => mult_21_C247_n1455,
                           Z => mult_21_C247_n663);
   mult_21_C247_U1377 : EXOR2D1 port map( A1 => N3033, A2 => N3032, Z => 
                           mult_21_C247_n1454);
   mult_21_C247_U1376 : MUXB2DL port map( A0 => N3207, A1 => N3208, SL => 
                           mult_21_C247_n1454, Z => mult_21_C247_n664);
   mult_21_C247_U1375 : MUXB2DL port map( A0 => N3206, A1 => N3207, SL => 
                           mult_21_C247_n1454, Z => mult_21_C247_n665);
   mult_21_C247_U1374 : MUXB2DL port map( A0 => mult_21_C247_n1387, A1 => N3206
                           , SL => mult_21_C247_n1454, Z => mult_21_C247_n666);
   mult_21_C247_U1373 : MUXB2DL port map( A0 => mult_21_C247_n1389, A1 => N3205
                           , SL => mult_21_C247_n1454, Z => mult_21_C247_n667);
   mult_21_C247_U1372 : MUXB2DL port map( A0 => N3203, A1 => mult_21_C247_n1390
                           , SL => mult_21_C247_n1454, Z => mult_21_C247_n668);
   mult_21_C247_U1371 : MUXB2DL port map( A0 => mult_21_C247_n1394, A1 => N3203
                           , SL => mult_21_C247_n1454, Z => mult_21_C247_n669);
   mult_21_C247_U1370 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C247_n1454, Z => mult_21_C247_n670);
   mult_21_C247_U1369 : NAN2D1 port map( A1 => N3201, A2 => mult_21_C247_n1454,
                           Z => mult_21_C247_n671);
   mult_21_C247_U1368 : MUXB2DL port map( A0 => N3209, A1 => N3210, SL => 
                           mult_21_C247_n1453, Z => mult_21_C247_n672);
   mult_21_C247_U1367 : MUXB2DL port map( A0 => N3208, A1 => N3209, SL => 
                           mult_21_C247_n1453, Z => mult_21_C247_n673);
   mult_21_C247_U1366 : MUXB2DL port map( A0 => N3207, A1 => N3208, SL => 
                           mult_21_C247_n1453, Z => mult_21_C247_n674);
   mult_21_C247_U1365 : MUXB2DL port map( A0 => N3206, A1 => N3207, SL => 
                           mult_21_C247_n1453, Z => mult_21_C247_n675);
   mult_21_C247_U1364 : MUXB2DL port map( A0 => N3205, A1 => mult_21_C247_n1385
                           , SL => mult_21_C247_n1453, Z => mult_21_C247_n676);
   mult_21_C247_U1363 : MUXB2DL port map( A0 => mult_21_C247_n1389, A1 => N3205
                           , SL => mult_21_C247_n1453, Z => mult_21_C247_n677);
   mult_21_C247_U1362 : MUXB2DL port map( A0 => N3203, A1 => mult_21_C247_n1390
                           , SL => mult_21_C247_n1453, Z => mult_21_C247_n678);
   mult_21_C247_U1361 : MUXB2DL port map( A0 => mult_21_C247_n1394, A1 => N3203
                           , SL => mult_21_C247_n1453, Z => mult_21_C247_n679);
   mult_21_C247_U1360 : AOI21D1 port map( A1 => N3024, A2 => N3025, B => 
                           mult_21_C247_n1415, Z => mult_21_C247_n946);
   mult_21_C247_U1359 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C247_n1453, Z => mult_21_C247_n680);
   mult_21_C247_U1358 : NAN2D1 port map( A1 => mult_21_C247_n1396, A2 => 
                           mult_21_C247_n1453, Z => mult_21_C247_n681);
   mult_21_C247_U1357 : MUXB2DL port map( A0 => N3211, A1 => N3212, SL => 
                           mult_21_C247_n1452, Z => mult_21_C247_n682);
   mult_21_C247_U1356 : MUXB2DL port map( A0 => N3210, A1 => N3211, SL => 
                           mult_21_C247_n1452, Z => mult_21_C247_n683);
   mult_21_C247_U1355 : MUXB2DL port map( A0 => N3209, A1 => N3210, SL => 
                           mult_21_C247_n1452, Z => mult_21_C247_n684);
   mult_21_C247_U1354 : MUXB2DL port map( A0 => N3208, A1 => N3209, SL => 
                           mult_21_C247_n1452, Z => mult_21_C247_n685);
   mult_21_C247_U1353 : MUXB2DL port map( A0 => N3207, A1 => N3208, SL => 
                           mult_21_C247_n1452, Z => mult_21_C247_n686);
   mult_21_C247_U1352 : MUXB2DL port map( A0 => N3206, A1 => N3207, SL => 
                           mult_21_C247_n1452, Z => mult_21_C247_n687);
   mult_21_C247_U1351 : MUXB2DL port map( A0 => mult_21_C247_n1387, A1 => 
                           mult_21_C247_n1385, SL => mult_21_C247_n1452, Z => 
                           mult_21_C247_n688);
   mult_21_C247_U1350 : MUXB2DL port map( A0 => mult_21_C247_n1389, A1 => N3205
                           , SL => mult_21_C247_n1452, Z => mult_21_C247_n689);
   mult_21_C247_U1349 : MUXB2DL port map( A0 => N3203, A1 => mult_21_C247_n1390
                           , SL => mult_21_C247_n1452, Z => mult_21_C247_n690);
   mult_21_C247_U1348 : MUXB2DL port map( A0 => mult_21_C247_n1394, A1 => N3203
                           , SL => mult_21_C247_n1452, Z => mult_21_C247_n691);
   mult_21_C247_U1347 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C247_n1452, Z => mult_21_C247_n692);
   mult_21_C247_U1346 : NAN2D1 port map( A1 => mult_21_C247_n1396, A2 => 
                           mult_21_C247_n1452, Z => mult_21_C247_n693);
   mult_21_C247_U1345 : MUXB2DL port map( A0 => N3213, A1 => N3214, SL => 
                           mult_21_C247_n1451, Z => mult_21_C247_n694);
   mult_21_C247_U1344 : MUXB2DL port map( A0 => N3212, A1 => N3213, SL => 
                           mult_21_C247_n1451, Z => mult_21_C247_n695);
   mult_21_C247_U1343 : MUXB2DL port map( A0 => N3211, A1 => N3212, SL => 
                           mult_21_C247_n1451, Z => mult_21_C247_n696);
   mult_21_C247_U1342 : MUXB2DL port map( A0 => N3210, A1 => N3211, SL => 
                           mult_21_C247_n1451, Z => mult_21_C247_n697);
   mult_21_C247_U1341 : MUXB2DL port map( A0 => N3209, A1 => N3210, SL => 
                           mult_21_C247_n1451, Z => mult_21_C247_n698);
   mult_21_C247_U1340 : MUXB2DL port map( A0 => N3208, A1 => N3209, SL => 
                           mult_21_C247_n1451, Z => mult_21_C247_n699);
   mult_21_C247_U1339 : MUXB2DL port map( A0 => N3207, A1 => N3208, SL => 
                           mult_21_C247_n1451, Z => mult_21_C247_n700);
   mult_21_C247_U1338 : MUXB2DL port map( A0 => N3206, A1 => N3207, SL => 
                           mult_21_C247_n1451, Z => mult_21_C247_n701);
   mult_21_C247_U1337 : MUXB2DL port map( A0 => mult_21_C247_n1387, A1 => 
                           mult_21_C247_n1385, SL => mult_21_C247_n1451, Z => 
                           mult_21_C247_n702);
   mult_21_C247_U1336 : MUXB2DL port map( A0 => mult_21_C247_n1389, A1 => N3205
                           , SL => mult_21_C247_n1451, Z => mult_21_C247_n703);
   mult_21_C247_U1335 : MUXB2DL port map( A0 => N3203, A1 => mult_21_C247_n1390
                           , SL => mult_21_C247_n1451, Z => mult_21_C247_n704);
   mult_21_C247_U1334 : MUXB2DL port map( A0 => mult_21_C247_n1394, A1 => 
                           mult_21_C247_n1392, SL => mult_21_C247_n1451, Z => 
                           mult_21_C247_n705);
   mult_21_C247_U1333 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C247_n1451, Z => mult_21_C247_n706);
   mult_21_C247_U1332 : NAN2D1 port map( A1 => mult_21_C247_n1396, A2 => 
                           mult_21_C247_n1451, Z => mult_21_C247_n707);
   mult_21_C247_U1331 : MUXB2DL port map( A0 => N3215, A1 => N3216, SL => 
                           mult_21_C247_n1450, Z => mult_21_C247_n708);
   mult_21_C247_U1330 : MUXB2DL port map( A0 => N3214, A1 => N3215, SL => 
                           mult_21_C247_n1450, Z => mult_21_C247_n709);
   mult_21_C247_U1329 : MUXB2DL port map( A0 => N3213, A1 => N3214, SL => 
                           mult_21_C247_n1450, Z => mult_21_C247_n710);
   mult_21_C247_U1328 : MUXB2DL port map( A0 => N3212, A1 => N3213, SL => 
                           mult_21_C247_n1450, Z => mult_21_C247_n711);
   mult_21_C247_U1327 : MUXB2DL port map( A0 => N3211, A1 => N3212, SL => 
                           mult_21_C247_n1450, Z => mult_21_C247_n712);
   mult_21_C247_U1326 : MUXB2DL port map( A0 => N3210, A1 => N3211, SL => 
                           mult_21_C247_n1450, Z => mult_21_C247_n713);
   mult_21_C247_U1325 : MUXB2DL port map( A0 => N3209, A1 => N3210, SL => 
                           mult_21_C247_n1450, Z => mult_21_C247_n714);
   mult_21_C247_U1324 : MUXB2DL port map( A0 => N3208, A1 => N3209, SL => 
                           mult_21_C247_n1450, Z => mult_21_C247_n715);
   mult_21_C247_U1323 : MUXB2DL port map( A0 => N3207, A1 => N3208, SL => 
                           mult_21_C247_n1450, Z => mult_21_C247_n716);
   mult_21_C247_U1322 : MUXB2DL port map( A0 => N3206, A1 => N3207, SL => 
                           mult_21_C247_n1450, Z => mult_21_C247_n717);
   mult_21_C247_U1321 : MUXB2DL port map( A0 => mult_21_C247_n1387, A1 => 
                           mult_21_C247_n1385, SL => mult_21_C247_n1450, Z => 
                           mult_21_C247_n718);
   mult_21_C247_U1320 : MUXB2DL port map( A0 => mult_21_C247_n1389, A1 => N3205
                           , SL => mult_21_C247_n1450, Z => mult_21_C247_n719);
   mult_21_C247_U1319 : MUXB2DL port map( A0 => N3203, A1 => mult_21_C247_n1390
                           , SL => mult_21_C247_n1450, Z => mult_21_C247_n720);
   mult_21_C247_U1318 : MUXB2DL port map( A0 => mult_21_C247_n1394, A1 => 
                           mult_21_C247_n1392, SL => mult_21_C247_n1450, Z => 
                           mult_21_C247_n721);
   mult_21_C247_U1317 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C247_n1450, Z => mult_21_C247_n722);
   mult_21_C247_U1316 : NAN2D1 port map( A1 => mult_21_C247_n1396, A2 => 
                           mult_21_C247_n1450, Z => mult_21_C247_n723);
   mult_21_C247_U1315 : MUXB2DL port map( A0 => N3217, A1 => N3218, SL => 
                           mult_21_C247_n1449, Z => mult_21_C247_n724);
   mult_21_C247_U1314 : MUXB2DL port map( A0 => N3216, A1 => N3217, SL => 
                           mult_21_C247_n1449, Z => mult_21_C247_n725);
   mult_21_C247_U1313 : MUXB2DL port map( A0 => N3215, A1 => N3216, SL => 
                           mult_21_C247_n1449, Z => mult_21_C247_n726);
   mult_21_C247_U1312 : MUXB2DL port map( A0 => N3214, A1 => N3215, SL => 
                           mult_21_C247_n1449, Z => mult_21_C247_n727);
   mult_21_C247_U1311 : MUXB2DL port map( A0 => N3213, A1 => N3214, SL => 
                           mult_21_C247_n1449, Z => mult_21_C247_n728);
   mult_21_C247_U1310 : MUXB2DL port map( A0 => N3212, A1 => N3213, SL => 
                           mult_21_C247_n1449, Z => mult_21_C247_n729);
   mult_21_C247_U1309 : MUXB2DL port map( A0 => N3211, A1 => N3212, SL => 
                           mult_21_C247_n1449, Z => mult_21_C247_n730);
   mult_21_C247_U1308 : MUXB2DL port map( A0 => N3210, A1 => N3211, SL => 
                           mult_21_C247_n1449, Z => mult_21_C247_n731);
   mult_21_C247_U1307 : MUXB2DL port map( A0 => N3209, A1 => N3210, SL => 
                           mult_21_C247_n1449, Z => mult_21_C247_n732);
   mult_21_C247_U1306 : MUXB2DL port map( A0 => N3208, A1 => N3209, SL => 
                           mult_21_C247_n1449, Z => mult_21_C247_n733);
   mult_21_C247_U1305 : MUXB2DL port map( A0 => N3207, A1 => N3208, SL => 
                           mult_21_C247_n1449, Z => mult_21_C247_n734);
   mult_21_C247_U1304 : MUXB2DL port map( A0 => N3206, A1 => N3207, SL => 
                           mult_21_C247_n1449, Z => mult_21_C247_n735);
   mult_21_C247_U1303 : MUXB2DL port map( A0 => mult_21_C247_n1387, A1 => 
                           mult_21_C247_n1385, SL => mult_21_C247_n1449, Z => 
                           mult_21_C247_n736);
   mult_21_C247_U1302 : MUXB2DL port map( A0 => mult_21_C247_n1389, A1 => N3205
                           , SL => mult_21_C247_n1449, Z => mult_21_C247_n737);
   mult_21_C247_U1301 : MUXB2DL port map( A0 => N3203, A1 => mult_21_C247_n1390
                           , SL => mult_21_C247_n1449, Z => mult_21_C247_n738);
   mult_21_C247_U1300 : MUXB2DL port map( A0 => mult_21_C247_n1394, A1 => 
                           mult_21_C247_n1392, SL => mult_21_C247_n1449, Z => 
                           mult_21_C247_n739);
   mult_21_C247_U1299 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C247_n1449, Z => mult_21_C247_n740);
   mult_21_C247_U1298 : NAN2D1 port map( A1 => mult_21_C247_n1396, A2 => 
                           mult_21_C247_n1449, Z => mult_21_C247_n741);
   mult_21_C247_U1297 : MUXB2DL port map( A0 => N3219, A1 => N3220, SL => 
                           mult_21_C247_n1448, Z => mult_21_C247_n742);
   mult_21_C247_U1296 : MUXB2DL port map( A0 => N3218, A1 => N3219, SL => 
                           mult_21_C247_n1448, Z => mult_21_C247_n743);
   mult_21_C247_U1295 : MUXB2DL port map( A0 => N3217, A1 => N3218, SL => 
                           mult_21_C247_n1448, Z => mult_21_C247_n744);
   mult_21_C247_U1294 : MUXB2DL port map( A0 => N3216, A1 => N3217, SL => 
                           mult_21_C247_n1448, Z => mult_21_C247_n745);
   mult_21_C247_U1293 : MUXB2DL port map( A0 => N3215, A1 => N3216, SL => 
                           mult_21_C247_n1448, Z => mult_21_C247_n746);
   mult_21_C247_U1292 : MUXB2DL port map( A0 => N3214, A1 => N3215, SL => 
                           mult_21_C247_n1448, Z => mult_21_C247_n747);
   mult_21_C247_U1291 : MUXB2DL port map( A0 => N3213, A1 => N3214, SL => 
                           mult_21_C247_n1448, Z => mult_21_C247_n748);
   mult_21_C247_U1290 : MUXB2DL port map( A0 => N3212, A1 => N3213, SL => 
                           mult_21_C247_n1448, Z => mult_21_C247_n749);
   mult_21_C247_U1289 : AOI21D1 port map( A1 => N3026, A2 => N3027, B => 
                           mult_21_C247_n1417, Z => mult_21_C247_n945);
   mult_21_C247_U1288 : MUXB2DL port map( A0 => N3211, A1 => N3212, SL => 
                           mult_21_C247_n1448, Z => mult_21_C247_n750);
   mult_21_C247_U1287 : MUXB2DL port map( A0 => N3210, A1 => N3211, SL => 
                           mult_21_C247_n1448, Z => mult_21_C247_n751);
   mult_21_C247_U1286 : MUXB2DL port map( A0 => N3209, A1 => N3210, SL => 
                           mult_21_C247_n1448, Z => mult_21_C247_n752);
   mult_21_C247_U1285 : MUXB2DL port map( A0 => N3208, A1 => N3209, SL => 
                           mult_21_C247_n1448, Z => mult_21_C247_n753);
   mult_21_C247_U1284 : MUXB2DL port map( A0 => N3207, A1 => N3208, SL => 
                           mult_21_C247_n1448, Z => mult_21_C247_n754);
   mult_21_C247_U1283 : MUXB2DL port map( A0 => N3206, A1 => N3207, SL => 
                           mult_21_C247_n1448, Z => mult_21_C247_n755);
   mult_21_C247_U1282 : MUXB2DL port map( A0 => mult_21_C247_n1387, A1 => 
                           mult_21_C247_n1385, SL => mult_21_C247_n1448, Z => 
                           mult_21_C247_n756);
   mult_21_C247_U1281 : MUXB2DL port map( A0 => mult_21_C247_n1389, A1 => N3205
                           , SL => mult_21_C247_n1448, Z => mult_21_C247_n757);
   mult_21_C247_U1280 : MUXB2DL port map( A0 => N3203, A1 => mult_21_C247_n1390
                           , SL => mult_21_C247_n1448, Z => mult_21_C247_n758);
   mult_21_C247_U1279 : MUXB2DL port map( A0 => N3202, A1 => mult_21_C247_n1392
                           , SL => mult_21_C247_n1448, Z => mult_21_C247_n759);
   mult_21_C247_U1278 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C247_n1448, Z => mult_21_C247_n760);
   mult_21_C247_U1277 : NAN2D1 port map( A1 => mult_21_C247_n1396, A2 => 
                           mult_21_C247_n1448, Z => mult_21_C247_n761);
   mult_21_C247_U1276 : MUXB2DL port map( A0 => N3221, A1 => N3222, SL => 
                           mult_21_C247_n1447, Z => mult_21_C247_n762);
   mult_21_C247_U1275 : MUXB2DL port map( A0 => N3220, A1 => N3221, SL => 
                           mult_21_C247_n1447, Z => mult_21_C247_n763);
   mult_21_C247_U1274 : MUXB2DL port map( A0 => N3219, A1 => N3220, SL => 
                           mult_21_C247_n1447, Z => mult_21_C247_n764);
   mult_21_C247_U1273 : MUXB2DL port map( A0 => N3218, A1 => N3219, SL => 
                           mult_21_C247_n1447, Z => mult_21_C247_n765);
   mult_21_C247_U1272 : MUXB2DL port map( A0 => N3217, A1 => N3218, SL => 
                           mult_21_C247_n1447, Z => mult_21_C247_n766);
   mult_21_C247_U1271 : MUXB2DL port map( A0 => N3216, A1 => N3217, SL => 
                           mult_21_C247_n1447, Z => mult_21_C247_n767);
   mult_21_C247_U1270 : MUXB2DL port map( A0 => N3215, A1 => N3216, SL => 
                           mult_21_C247_n1447, Z => mult_21_C247_n768);
   mult_21_C247_U1269 : MUXB2DL port map( A0 => N3214, A1 => N3215, SL => 
                           mult_21_C247_n1447, Z => mult_21_C247_n769);
   mult_21_C247_U1268 : MUXB2DL port map( A0 => N3213, A1 => N3214, SL => 
                           mult_21_C247_n1447, Z => mult_21_C247_n770);
   mult_21_C247_U1267 : MUXB2DL port map( A0 => N3212, A1 => N3213, SL => 
                           mult_21_C247_n1447, Z => mult_21_C247_n771);
   mult_21_C247_U1266 : MUXB2DL port map( A0 => N3211, A1 => N3212, SL => 
                           mult_21_C247_n1447, Z => mult_21_C247_n772);
   mult_21_C247_U1265 : MUXB2DL port map( A0 => N3210, A1 => N3211, SL => 
                           mult_21_C247_n1447, Z => mult_21_C247_n773);
   mult_21_C247_U1264 : MUXB2DL port map( A0 => N3209, A1 => N3210, SL => 
                           mult_21_C247_n1447, Z => mult_21_C247_n774);
   mult_21_C247_U1263 : MUXB2DL port map( A0 => N3208, A1 => N3209, SL => 
                           mult_21_C247_n1447, Z => mult_21_C247_n775);
   mult_21_C247_U1262 : MUXB2DL port map( A0 => N3207, A1 => N3208, SL => 
                           mult_21_C247_n1447, Z => mult_21_C247_n776);
   mult_21_C247_U1261 : MUXB2DL port map( A0 => N3206, A1 => N3207, SL => 
                           mult_21_C247_n1447, Z => mult_21_C247_n777);
   mult_21_C247_U1260 : MUXB2DL port map( A0 => mult_21_C247_n1387, A1 => 
                           mult_21_C247_n1385, SL => mult_21_C247_n1447, Z => 
                           mult_21_C247_n778);
   mult_21_C247_U1259 : MUXB2DL port map( A0 => mult_21_C247_n1390, A1 => N3205
                           , SL => mult_21_C247_n1447, Z => mult_21_C247_n779);
   mult_21_C247_U1258 : MUXB2DL port map( A0 => mult_21_C247_n1392, A1 => 
                           mult_21_C247_n1390, SL => mult_21_C247_n1447, Z => 
                           mult_21_C247_n780);
   mult_21_C247_U1257 : MUXB2DL port map( A0 => mult_21_C247_n1394, A1 => 
                           mult_21_C247_n1392, SL => mult_21_C247_n1447, Z => 
                           mult_21_C247_n781);
   mult_21_C247_U1256 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C247_n1447, Z => mult_21_C247_n782);
   mult_21_C247_U1255 : NAN2D1 port map( A1 => mult_21_C247_n1396, A2 => 
                           mult_21_C247_n1447, Z => mult_21_C247_n783);
   mult_21_C247_U1254 : MUXB2DL port map( A0 => N3223, A1 => N3224, SL => 
                           mult_21_C247_n1377, Z => mult_21_C247_n784);
   mult_21_C247_U1253 : MUXB2DL port map( A0 => N3222, A1 => N3223, SL => 
                           mult_21_C247_n1377, Z => mult_21_C247_n785);
   mult_21_C247_U1252 : MUXB2DL port map( A0 => N3221, A1 => N3222, SL => 
                           mult_21_C247_n1377, Z => mult_21_C247_n786);
   mult_21_C247_U1251 : MUXB2DL port map( A0 => N3220, A1 => N3221, SL => 
                           mult_21_C247_n1377, Z => mult_21_C247_n787);
   mult_21_C247_U1250 : MUXB2DL port map( A0 => N3219, A1 => N3220, SL => 
                           mult_21_C247_n1377, Z => mult_21_C247_n788);
   mult_21_C247_U1249 : MUXB2DL port map( A0 => N3218, A1 => N3219, SL => 
                           mult_21_C247_n1377, Z => mult_21_C247_n789);
   mult_21_C247_U1248 : MUXB2DL port map( A0 => N3217, A1 => N3218, SL => 
                           mult_21_C247_n1377, Z => mult_21_C247_n790);
   mult_21_C247_U1247 : MUXB2DL port map( A0 => N3216, A1 => N3217, SL => 
                           mult_21_C247_n1377, Z => mult_21_C247_n791);
   mult_21_C247_U1246 : MUXB2DL port map( A0 => N3215, A1 => N3216, SL => 
                           mult_21_C247_n1377, Z => mult_21_C247_n792);
   mult_21_C247_U1245 : MUXB2DL port map( A0 => N3214, A1 => N3215, SL => 
                           mult_21_C247_n1377, Z => mult_21_C247_n793);
   mult_21_C247_U1244 : MUXB2DL port map( A0 => N3213, A1 => N3214, SL => 
                           mult_21_C247_n1377, Z => mult_21_C247_n794);
   mult_21_C247_U1243 : MUXB2DL port map( A0 => N3212, A1 => N3213, SL => 
                           mult_21_C247_n1377, Z => mult_21_C247_n795);
   mult_21_C247_U1242 : MUXB2DL port map( A0 => N3211, A1 => N3212, SL => 
                           mult_21_C247_n1377, Z => mult_21_C247_n796);
   mult_21_C247_U1241 : MUXB2DL port map( A0 => N3210, A1 => N3211, SL => 
                           mult_21_C247_n1377, Z => mult_21_C247_n797);
   mult_21_C247_U1240 : MUXB2DL port map( A0 => N3209, A1 => N3210, SL => 
                           mult_21_C247_n1377, Z => mult_21_C247_n798);
   mult_21_C247_U1239 : MUXB2DL port map( A0 => N3208, A1 => N3209, SL => 
                           mult_21_C247_n1377, Z => mult_21_C247_n799);
   mult_21_C247_U1238 : MUXB2DL port map( A0 => N3207, A1 => N3208, SL => 
                           mult_21_C247_n1377, Z => mult_21_C247_n800);
   mult_21_C247_U1237 : MUXB2DL port map( A0 => N3206, A1 => N3207, SL => 
                           mult_21_C247_n1377, Z => mult_21_C247_n801);
   mult_21_C247_U1236 : MUXB2DL port map( A0 => mult_21_C247_n1387, A1 => 
                           mult_21_C247_n1385, SL => mult_21_C247_n1377, Z => 
                           mult_21_C247_n802);
   mult_21_C247_U1235 : MUXB2DL port map( A0 => mult_21_C247_n1389, A1 => 
                           mult_21_C247_n1387, SL => mult_21_C247_n1377, Z => 
                           mult_21_C247_n803);
   mult_21_C247_U1234 : MUXB2DL port map( A0 => N3203, A1 => mult_21_C247_n1390
                           , SL => mult_21_C247_n1377, Z => mult_21_C247_n804);
   mult_21_C247_U1233 : MUXB2DL port map( A0 => N3202, A1 => mult_21_C247_n1392
                           , SL => mult_21_C247_n1377, Z => mult_21_C247_n805);
   mult_21_C247_U1232 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C247_n1377, Z => mult_21_C247_n806);
   mult_21_C247_U1231 : NAN2D1 port map( A1 => mult_21_C247_n1396, A2 => 
                           mult_21_C247_n1377, Z => mult_21_C247_n807);
   mult_21_C247_U1230 : MUXB2DL port map( A0 => N3225, A1 => N3226, SL => 
                           mult_21_C247_n1376, Z => mult_21_C247_n808);
   mult_21_C247_U1229 : MUXB2DL port map( A0 => N3224, A1 => N3225, SL => 
                           mult_21_C247_n1376, Z => mult_21_C247_n809);
   mult_21_C247_U1228 : AOI21D1 port map( A1 => N3028, A2 => N3029, B => 
                           mult_21_C247_n1419, Z => mult_21_C247_n944);
   mult_21_C247_U1227 : MUXB2DL port map( A0 => N3223, A1 => N3224, SL => 
                           mult_21_C247_n1376, Z => mult_21_C247_n810);
   mult_21_C247_U1226 : MUXB2DL port map( A0 => N3222, A1 => N3223, SL => 
                           mult_21_C247_n1376, Z => mult_21_C247_n811);
   mult_21_C247_U1225 : MUXB2DL port map( A0 => N3221, A1 => N3222, SL => 
                           mult_21_C247_n1376, Z => mult_21_C247_n812);
   mult_21_C247_U1224 : MUXB2DL port map( A0 => N3220, A1 => N3221, SL => 
                           mult_21_C247_n1376, Z => mult_21_C247_n813);
   mult_21_C247_U1223 : MUXB2DL port map( A0 => N3219, A1 => N3220, SL => 
                           mult_21_C247_n1376, Z => mult_21_C247_n814);
   mult_21_C247_U1222 : MUXB2DL port map( A0 => N3218, A1 => N3219, SL => 
                           mult_21_C247_n1376, Z => mult_21_C247_n815);
   mult_21_C247_U1221 : MUXB2DL port map( A0 => N3217, A1 => N3218, SL => 
                           mult_21_C247_n1376, Z => mult_21_C247_n816);
   mult_21_C247_U1220 : MUXB2DL port map( A0 => N3216, A1 => N3217, SL => 
                           mult_21_C247_n1376, Z => mult_21_C247_n817);
   mult_21_C247_U1219 : MUXB2DL port map( A0 => N3215, A1 => N3216, SL => 
                           mult_21_C247_n1376, Z => mult_21_C247_n818);
   mult_21_C247_U1218 : MUXB2DL port map( A0 => N3214, A1 => N3215, SL => 
                           mult_21_C247_n1376, Z => mult_21_C247_n819);
   mult_21_C247_U1217 : MUXB2DL port map( A0 => N3213, A1 => N3214, SL => 
                           mult_21_C247_n1376, Z => mult_21_C247_n820);
   mult_21_C247_U1216 : MUXB2DL port map( A0 => N3212, A1 => N3213, SL => 
                           mult_21_C247_n1376, Z => mult_21_C247_n821);
   mult_21_C247_U1215 : MUXB2DL port map( A0 => N3211, A1 => N3212, SL => 
                           mult_21_C247_n1376, Z => mult_21_C247_n822);
   mult_21_C247_U1214 : MUXB2DL port map( A0 => N3210, A1 => N3211, SL => 
                           mult_21_C247_n1376, Z => mult_21_C247_n823);
   mult_21_C247_U1213 : MUXB2DL port map( A0 => N3209, A1 => N3210, SL => 
                           mult_21_C247_n1376, Z => mult_21_C247_n824);
   mult_21_C247_U1212 : MUXB2DL port map( A0 => N3208, A1 => N3209, SL => 
                           mult_21_C247_n1376, Z => mult_21_C247_n825);
   mult_21_C247_U1211 : MUXB2DL port map( A0 => N3207, A1 => N3208, SL => 
                           mult_21_C247_n1376, Z => mult_21_C247_n826);
   mult_21_C247_U1210 : MUXB2DL port map( A0 => N3206, A1 => N3207, SL => 
                           mult_21_C247_n1376, Z => mult_21_C247_n827);
   mult_21_C247_U1209 : MUXB2DL port map( A0 => mult_21_C247_n1387, A1 => 
                           mult_21_C247_n1385, SL => mult_21_C247_n1376, Z => 
                           mult_21_C247_n828);
   mult_21_C247_U1208 : MUXB2DL port map( A0 => mult_21_C247_n1389, A1 => 
                           mult_21_C247_n1387, SL => mult_21_C247_n1376, Z => 
                           mult_21_C247_n829);
   mult_21_C247_U1207 : MUXB2DL port map( A0 => mult_21_C247_n1392, A1 => 
                           mult_21_C247_n1390, SL => mult_21_C247_n1376, Z => 
                           mult_21_C247_n830);
   mult_21_C247_U1206 : MUXB2DL port map( A0 => mult_21_C247_n1394, A1 => 
                           mult_21_C247_n1392, SL => mult_21_C247_n1376, Z => 
                           mult_21_C247_n831);
   mult_21_C247_U1205 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C247_n1376, Z => mult_21_C247_n832);
   mult_21_C247_U1204 : NAN2D1 port map( A1 => mult_21_C247_n1396, A2 => 
                           mult_21_C247_n1376, Z => mult_21_C247_n833);
   mult_21_C247_U1203 : MUXB2DL port map( A0 => N3227, A1 => N3228, SL => 
                           mult_21_C247_n1375, Z => mult_21_C247_n834);
   mult_21_C247_U1202 : MUXB2DL port map( A0 => N3226, A1 => N3227, SL => 
                           mult_21_C247_n1375, Z => mult_21_C247_n835);
   mult_21_C247_U1201 : MUXB2DL port map( A0 => N3225, A1 => N3226, SL => 
                           mult_21_C247_n1375, Z => mult_21_C247_n836);
   mult_21_C247_U1200 : MUXB2DL port map( A0 => N3224, A1 => N3225, SL => 
                           mult_21_C247_n1375, Z => mult_21_C247_n837);
   mult_21_C247_U1199 : MUXB2DL port map( A0 => N3223, A1 => N3224, SL => 
                           mult_21_C247_n1375, Z => mult_21_C247_n838);
   mult_21_C247_U1198 : MUXB2DL port map( A0 => N3222, A1 => N3223, SL => 
                           mult_21_C247_n1375, Z => mult_21_C247_n839);
   mult_21_C247_U1197 : MUXB2DL port map( A0 => N3221, A1 => N3222, SL => 
                           mult_21_C247_n1375, Z => mult_21_C247_n840);
   mult_21_C247_U1196 : MUXB2DL port map( A0 => N3220, A1 => N3221, SL => 
                           mult_21_C247_n1375, Z => mult_21_C247_n841);
   mult_21_C247_U1195 : MUXB2DL port map( A0 => N3219, A1 => N3220, SL => 
                           mult_21_C247_n1375, Z => mult_21_C247_n842);
   mult_21_C247_U1194 : MUXB2DL port map( A0 => N3218, A1 => N3219, SL => 
                           mult_21_C247_n1375, Z => mult_21_C247_n843);
   mult_21_C247_U1193 : MUXB2DL port map( A0 => N3217, A1 => N3218, SL => 
                           mult_21_C247_n1375, Z => mult_21_C247_n844);
   mult_21_C247_U1192 : MUXB2DL port map( A0 => N3216, A1 => N3217, SL => 
                           mult_21_C247_n1375, Z => mult_21_C247_n845);
   mult_21_C247_U1191 : MUXB2DL port map( A0 => N3215, A1 => N3216, SL => 
                           mult_21_C247_n1375, Z => mult_21_C247_n846);
   mult_21_C247_U1190 : MUXB2DL port map( A0 => N3214, A1 => N3215, SL => 
                           mult_21_C247_n1375, Z => mult_21_C247_n847);
   mult_21_C247_U1189 : MUXB2DL port map( A0 => N3213, A1 => N3214, SL => 
                           mult_21_C247_n1375, Z => mult_21_C247_n848);
   mult_21_C247_U1188 : MUXB2DL port map( A0 => N3212, A1 => N3213, SL => 
                           mult_21_C247_n1375, Z => mult_21_C247_n849);
   mult_21_C247_U1187 : MUXB2DL port map( A0 => N3211, A1 => N3212, SL => 
                           mult_21_C247_n1375, Z => mult_21_C247_n850);
   mult_21_C247_U1186 : MUXB2DL port map( A0 => N3210, A1 => N3211, SL => 
                           mult_21_C247_n1375, Z => mult_21_C247_n851);
   mult_21_C247_U1185 : MUXB2DL port map( A0 => N3209, A1 => N3210, SL => 
                           mult_21_C247_n1375, Z => mult_21_C247_n852);
   mult_21_C247_U1184 : MUXB2DL port map( A0 => N3208, A1 => N3209, SL => 
                           mult_21_C247_n1375, Z => mult_21_C247_n853);
   mult_21_C247_U1183 : MUXB2DL port map( A0 => N3207, A1 => N3208, SL => 
                           mult_21_C247_n1375, Z => mult_21_C247_n854);
   mult_21_C247_U1182 : MUXB2DL port map( A0 => N3206, A1 => N3207, SL => 
                           mult_21_C247_n1375, Z => mult_21_C247_n855);
   mult_21_C247_U1181 : MUXB2DL port map( A0 => mult_21_C247_n1387, A1 => 
                           mult_21_C247_n1385, SL => mult_21_C247_n1375, Z => 
                           mult_21_C247_n856);
   mult_21_C247_U1180 : MUXB2DL port map( A0 => mult_21_C247_n1389, A1 => 
                           mult_21_C247_n1387, SL => mult_21_C247_n1375, Z => 
                           mult_21_C247_n857);
   mult_21_C247_U1179 : MUXB2DL port map( A0 => N3203, A1 => mult_21_C247_n1390
                           , SL => mult_21_C247_n1375, Z => mult_21_C247_n858);
   mult_21_C247_U1178 : MUXB2DL port map( A0 => mult_21_C247_n1394, A1 => 
                           mult_21_C247_n1392, SL => mult_21_C247_n1375, Z => 
                           mult_21_C247_n859);
   mult_21_C247_U1177 : AOI21D1 port map( A1 => N3030, A2 => N3031, B => 
                           mult_21_C247_n1421, Z => mult_21_C247_n943);
   mult_21_C247_U1176 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C247_n1375, Z => mult_21_C247_n860);
   mult_21_C247_U1175 : NAN2D1 port map( A1 => mult_21_C247_n1396, A2 => 
                           mult_21_C247_n1375, Z => mult_21_C247_n861);
   mult_21_C247_U1174 : MUXB2DL port map( A0 => N3228, A1 => N3229, SL => 
                           mult_21_C247_n1384, Z => mult_21_C247_n863);
   mult_21_C247_U1173 : MUXB2DL port map( A0 => N3227, A1 => N3228, SL => 
                           mult_21_C247_n1384, Z => mult_21_C247_n864);
   mult_21_C247_U1172 : MUXB2DL port map( A0 => N3226, A1 => N3227, SL => 
                           mult_21_C247_n1384, Z => mult_21_C247_n865);
   mult_21_C247_U1171 : MUXB2DL port map( A0 => N3225, A1 => N3226, SL => 
                           mult_21_C247_n1384, Z => mult_21_C247_n866);
   mult_21_C247_U1170 : MUXB2DL port map( A0 => N3224, A1 => N3225, SL => 
                           mult_21_C247_n1384, Z => mult_21_C247_n867);
   mult_21_C247_U1169 : MUXB2DL port map( A0 => N3223, A1 => N3224, SL => 
                           mult_21_C247_n1384, Z => mult_21_C247_n868);
   mult_21_C247_U1168 : MUXB2DL port map( A0 => N3222, A1 => N3223, SL => 
                           mult_21_C247_n1384, Z => mult_21_C247_n869);
   mult_21_C247_U1167 : MUXB2DL port map( A0 => N3221, A1 => N3222, SL => 
                           mult_21_C247_n1384, Z => mult_21_C247_n870);
   mult_21_C247_U1166 : MUXB2DL port map( A0 => N3220, A1 => N3221, SL => 
                           mult_21_C247_n1384, Z => mult_21_C247_n871);
   mult_21_C247_U1165 : MUXB2DL port map( A0 => N3219, A1 => N3220, SL => 
                           mult_21_C247_n1384, Z => mult_21_C247_n872);
   mult_21_C247_U1164 : MUXB2DL port map( A0 => N3218, A1 => N3219, SL => 
                           mult_21_C247_n1384, Z => mult_21_C247_n873);
   mult_21_C247_U1163 : MUXB2DL port map( A0 => N3217, A1 => N3218, SL => 
                           mult_21_C247_n1384, Z => mult_21_C247_n874);
   mult_21_C247_U1162 : MUXB2DL port map( A0 => N3216, A1 => N3217, SL => 
                           mult_21_C247_n1384, Z => mult_21_C247_n875);
   mult_21_C247_U1161 : MUXB2DL port map( A0 => N3215, A1 => N3216, SL => 
                           mult_21_C247_n1384, Z => mult_21_C247_n876);
   mult_21_C247_U1160 : MUXB2DL port map( A0 => N3214, A1 => N3215, SL => 
                           mult_21_C247_n1384, Z => mult_21_C247_n877);
   mult_21_C247_U1159 : MUXB2DL port map( A0 => N3213, A1 => N3214, SL => 
                           mult_21_C247_n1384, Z => mult_21_C247_n878);
   mult_21_C247_U1158 : MUXB2DL port map( A0 => N3212, A1 => N3213, SL => 
                           mult_21_C247_n1384, Z => mult_21_C247_n879);
   mult_21_C247_U1157 : MUXB2DL port map( A0 => N3211, A1 => N3212, SL => 
                           mult_21_C247_n1384, Z => mult_21_C247_n880);
   mult_21_C247_U1156 : MUXB2DL port map( A0 => N3210, A1 => N3211, SL => 
                           mult_21_C247_n1384, Z => mult_21_C247_n881);
   mult_21_C247_U1155 : MUXB2DL port map( A0 => N3209, A1 => N3210, SL => 
                           mult_21_C247_n1384, Z => mult_21_C247_n882);
   mult_21_C247_U1154 : MUXB2DL port map( A0 => N3208, A1 => N3209, SL => 
                           mult_21_C247_n1384, Z => mult_21_C247_n883);
   mult_21_C247_U1153 : MUXB2DL port map( A0 => N3207, A1 => N3208, SL => 
                           mult_21_C247_n1384, Z => mult_21_C247_n884);
   mult_21_C247_U1152 : MUXB2DL port map( A0 => N3206, A1 => N3207, SL => 
                           mult_21_C247_n1384, Z => mult_21_C247_n885);
   mult_21_C247_U1151 : MUXB2DL port map( A0 => mult_21_C247_n1387, A1 => 
                           mult_21_C247_n1385, SL => mult_21_C247_n1384, Z => 
                           mult_21_C247_n886);
   mult_21_C247_U1150 : MUXB2DL port map( A0 => mult_21_C247_n1389, A1 => 
                           mult_21_C247_n1387, SL => mult_21_C247_n1384, Z => 
                           mult_21_C247_n887);
   mult_21_C247_U1149 : MUXB2DL port map( A0 => N3203, A1 => mult_21_C247_n1390
                           , SL => mult_21_C247_n1384, Z => mult_21_C247_n888);
   mult_21_C247_U1148 : MUXB2DL port map( A0 => mult_21_C247_n1394, A1 => 
                           mult_21_C247_n1392, SL => mult_21_C247_n1384, Z => 
                           mult_21_C247_n889);
   mult_21_C247_U1147 : OAI21D1 port map( A1 => N3033, A2 => N3032, B => 
                           mult_21_C247_n1423, Z => mult_21_C247_n89);
   mult_21_C247_U1146 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C247_n1384, Z => mult_21_C247_n890);
   mult_21_C247_U1145 : NAN2D1 port map( A1 => mult_21_C247_n1396, A2 => 
                           mult_21_C247_n1384, Z => mult_21_C247_n891);
   mult_21_C247_U1144 : MUXB2DL port map( A0 => N3231, A1 => N3232, SL => N3009
                           , Z => mult_21_C247_n892);
   mult_21_C247_U1143 : MUXB2DL port map( A0 => N3230, A1 => N3231, SL => N3009
                           , Z => mult_21_C247_n893);
   mult_21_C247_U1142 : MUXB2DL port map( A0 => N3229, A1 => N3230, SL => N3009
                           , Z => mult_21_C247_n894);
   mult_21_C247_U1141 : MUXB2DL port map( A0 => N3228, A1 => N3229, SL => N3009
                           , Z => mult_21_C247_n895);
   mult_21_C247_U1140 : MUXB2DL port map( A0 => N3227, A1 => N3228, SL => N3009
                           , Z => mult_21_C247_n896);
   mult_21_C247_U1139 : MUXB2DL port map( A0 => N3226, A1 => N3227, SL => N3009
                           , Z => mult_21_C247_n897);
   mult_21_C247_U1138 : MUXB2DL port map( A0 => N3225, A1 => N3226, SL => N3009
                           , Z => mult_21_C247_n898);
   mult_21_C247_U1137 : MUXB2DL port map( A0 => N3224, A1 => N3225, SL => N3009
                           , Z => mult_21_C247_n899);
   mult_21_C247_U1136 : MUXB2DL port map( A0 => N3223, A1 => N3224, SL => N3009
                           , Z => mult_21_C247_n900);
   mult_21_C247_U1135 : MUXB2DL port map( A0 => N3222, A1 => N3223, SL => N3009
                           , Z => mult_21_C247_n901);
   mult_21_C247_U1134 : MUXB2DL port map( A0 => N3221, A1 => N3222, SL => N3009
                           , Z => mult_21_C247_n902);
   mult_21_C247_U1133 : MUXB2DL port map( A0 => N3220, A1 => N3221, SL => N3009
                           , Z => mult_21_C247_n903);
   mult_21_C247_U1132 : MUXB2DL port map( A0 => N3219, A1 => N3220, SL => N3009
                           , Z => mult_21_C247_n904);
   mult_21_C247_U1131 : MUXB2DL port map( A0 => N3218, A1 => N3219, SL => N3009
                           , Z => mult_21_C247_n905);
   mult_21_C247_U1130 : MUXB2DL port map( A0 => N3217, A1 => N3218, SL => N3009
                           , Z => mult_21_C247_n906);
   mult_21_C247_U1129 : MUXB2DL port map( A0 => N3216, A1 => N3217, SL => N3009
                           , Z => mult_21_C247_n907);
   mult_21_C247_U1128 : MUXB2DL port map( A0 => N3215, A1 => N3216, SL => N3009
                           , Z => mult_21_C247_n908);
   mult_21_C247_U1127 : MUXB2DL port map( A0 => N3214, A1 => N3215, SL => N3009
                           , Z => mult_21_C247_n909);
   mult_21_C247_U1126 : AOI21D1 port map( A1 => N3032, A2 => N3033, B => 
                           mult_21_C247_n1423, Z => mult_21_C247_n942);
   mult_21_C247_U1125 : MUXB2DL port map( A0 => N3213, A1 => N3214, SL => N3009
                           , Z => mult_21_C247_n910);
   mult_21_C247_U1124 : MUXB2DL port map( A0 => N3212, A1 => N3213, SL => N3009
                           , Z => mult_21_C247_n911);
   mult_21_C247_U1123 : MUXB2DL port map( A0 => N3211, A1 => N3212, SL => N3009
                           , Z => mult_21_C247_n912);
   mult_21_C247_U1122 : MUXB2DL port map( A0 => N3210, A1 => N3211, SL => N3009
                           , Z => mult_21_C247_n913);
   mult_21_C247_U1121 : MUXB2DL port map( A0 => N3209, A1 => N3210, SL => N3009
                           , Z => mult_21_C247_n914);
   mult_21_C247_U1120 : MUXB2DL port map( A0 => N3208, A1 => N3209, SL => N3009
                           , Z => mult_21_C247_n915);
   mult_21_C247_U1119 : MUXB2DL port map( A0 => N3207, A1 => N3208, SL => N3009
                           , Z => mult_21_C247_n916);
   mult_21_C247_U1118 : MUXB2DL port map( A0 => N3206, A1 => N3207, SL => N3009
                           , Z => mult_21_C247_n917);
   mult_21_C247_U1117 : MUXB2DL port map( A0 => mult_21_C247_n1387, A1 => 
                           mult_21_C247_n1385, SL => N3009, Z => 
                           mult_21_C247_n918);
   mult_21_C247_U1116 : MUXB2DL port map( A0 => mult_21_C247_n1389, A1 => N3205
                           , SL => N3009, Z => mult_21_C247_n919);
   mult_21_C247_U1115 : MUXB2DL port map( A0 => mult_21_C247_n1392, A1 => 
                           mult_21_C247_n1390, SL => N3009, Z => 
                           mult_21_C247_n920);
   mult_21_C247_U1114 : MUXB2DL port map( A0 => mult_21_C247_n1394, A1 => 
                           mult_21_C247_n1392, SL => N3009, Z => 
                           mult_21_C247_n921);
   mult_21_C247_U1113 : MUXB2DL port map( A0 => mult_21_C247_n1396, A1 => N3202
                           , SL => N3009, Z => mult_21_C247_n922);
   mult_21_C247_U1112 : NAN2D1 port map( A1 => mult_21_C247_n1396, A2 => N3009,
                           Z => mult_21_C247_n923);
   mult_21_C247_U1111 : OAI21D1 port map( A1 => N3035, A2 => N3034, B => 
                           mult_21_C247_n1424, Z => mult_21_C247_n94);
   mult_21_C247_U1110 : AOI21D1 port map( A1 => N3034, A2 => N3035, B => 
                           mult_21_C247_n1424, Z => mult_21_C247_n941);
   mult_21_C247_U1109 : OAI21D1 port map( A1 => N3037, A2 => N3036, B => 
                           mult_21_C247_n1427, Z => mult_21_C247_n99);
   mult_21_C247_U1108 : EXOR2D1 port map( A1 => mult_21_C247_n230, A2 => 
                           mult_21_C247_n228, Z => mult_21_C247_n1446);
   mult_21_C247_U1107 : EXOR3D1 port map( A1 => mult_21_C247_n226, A2 => 
                           mult_21_C247_n224, A3 => mult_21_C247_n1446, Z => 
                           mult_21_C247_n1441);
   mult_21_C247_U1106 : EXOR2D1 port map( A1 => mult_21_C247_n222, A2 => 
                           mult_21_C247_n220, Z => mult_21_C247_n1445);
   mult_21_C247_U1105 : EXOR3D1 port map( A1 => mult_21_C247_n216, A2 => 
                           mult_21_C247_n1195, A3 => mult_21_C247_n1445, Z => 
                           mult_21_C247_n1442);
   mult_21_C247_U1104 : EXOR3D1 port map( A1 => mult_21_C247_n1165, A2 => 
                           mult_21_C247_n1137, A3 => mult_21_C247_n1045, Z => 
                           mult_21_C247_n1444);
   mult_21_C247_U1103 : EXOR3D1 port map( A1 => mult_21_C247_n1027, A2 => 
                           mult_21_C247_n1011, A3 => mult_21_C247_n1444, Z => 
                           mult_21_C247_n1443);
   mult_21_C247_U1102 : EXOR3D1 port map( A1 => mult_21_C247_n1441, A2 => 
                           mult_21_C247_n1442, A3 => mult_21_C247_n1443, Z => 
                           mult_21_C247_n1433);
   mult_21_C247_U1101 : EXOR2D1 port map( A1 => mult_21_C247_n985, A2 => 
                           mult_21_C247_n967, Z => mult_21_C247_n1440);
   mult_21_C247_U1100 : EXOR3D1 port map( A1 => mult_21_C247_n961, A2 => 
                           mult_21_C247_n218, A3 => mult_21_C247_n1440, Z => 
                           mult_21_C247_n1437);
   mult_21_C247_U1099 : EXNOR2D1 port map( A1 => mult_21_C247_n210, A2 => 
                           mult_21_C247_n1111, Z => mult_21_C247_n1439);
   mult_21_C247_U1098 : EXOR3D1 port map( A1 => mult_21_C247_n1087, A2 => 
                           mult_21_C247_n1065, A3 => mult_21_C247_n1439, Z => 
                           mult_21_C247_n1438);
   mult_21_C247_U1097 : EXOR3D1 port map( A1 => mult_21_C247_n1437, A2 => 
                           mult_21_C247_n204, A3 => mult_21_C247_n1438, Z => 
                           mult_21_C247_n1434);
   mult_21_C247_U1096 : EXNOR2D1 port map( A1 => mult_21_C247_n997, A2 => 
                           mult_21_C247_n975, Z => mult_21_C247_n1436);
   mult_21_C247_U1095 : EXOR3D1 port map( A1 => mult_21_C247_n957, A2 => 
                           mult_21_C247_n955, A3 => mult_21_C247_n1436, Z => 
                           mult_21_C247_n1435);
   mult_21_C247_U1094 : EXOR3D1 port map( A1 => mult_21_C247_n1433, A2 => 
                           mult_21_C247_n1434, A3 => mult_21_C247_n1435, Z => 
                           mult_21_C247_n1429);
   mult_21_C247_U1093 : EXOR2D1 port map( A1 => mult_21_C247_n202, A2 => 
                           mult_21_C247_n156, Z => mult_21_C247_n1430);
   mult_21_C247_U1092 : EXOR2D1 port map( A1 => mult_21_C247_n214, A2 => 
                           mult_21_C247_n212, Z => mult_21_C247_n1432);
   mult_21_C247_U1091 : EXOR3D1 port map( A1 => mult_21_C247_n208, A2 => 
                           mult_21_C247_n206, A3 => mult_21_C247_n1432, Z => 
                           mult_21_C247_n1431);
   mult_21_C247_U1090 : EXOR3D1 port map( A1 => mult_21_C247_n1429, A2 => 
                           mult_21_C247_n1430, A3 => mult_21_C247_n1431, Z => 
                           N3360);
   mult_21_C247_U1089 : INVD1 port map( A => N3040, Z => mult_21_C247_n1428);
   mult_21_C247_U1088 : MUXB2DL port map( A0 => N3230, A1 => N3229, SL => 
                           mult_21_C247_n1383, Z => mult_21_C247_n862);
   mult_21_C247_U1087 : INVD1 port map( A => N3038, Z => mult_21_C247_n1427);
   mult_21_C247_U1086 : INVD1 port map( A => N3036, Z => mult_21_C247_n1424);
   mult_21_C247_U1085 : INVD1 port map( A => N3034, Z => mult_21_C247_n1423);
   mult_21_C247_U1084 : OAI21D1 port map( A1 => N3031, A2 => N3030, B => 
                           mult_21_C247_n1421, Z => mult_21_C247_n84);
   mult_21_C247_U1083 : INVD1 port map( A => N3032, Z => mult_21_C247_n1421);
   mult_21_C247_U1082 : EXOR2D1 port map( A1 => N3031, A2 => N3030, Z => 
                           mult_21_C247_n1453);
   mult_21_C247_U1081 : OAI21D1 port map( A1 => N3029, A2 => N3028, B => 
                           mult_21_C247_n1419, Z => mult_21_C247_n80);
   mult_21_C247_U1080 : INVD1 port map( A => N3030, Z => mult_21_C247_n1419);
   mult_21_C247_U1079 : EXOR2D1 port map( A1 => N3029, A2 => N3028, Z => 
                           mult_21_C247_n1452);
   mult_21_C247_U1078 : OAI21D1 port map( A1 => N3027, A2 => N3026, B => 
                           mult_21_C247_n1417, Z => mult_21_C247_n73);
   mult_21_C247_U1077 : INVD1 port map( A => N3028, Z => mult_21_C247_n1417);
   mult_21_C247_U1076 : EXOR2D1 port map( A1 => N3027, A2 => N3026, Z => 
                           mult_21_C247_n1451);
   mult_21_C247_U1075 : OAI21D1 port map( A1 => N3025, A2 => N3024, B => 
                           mult_21_C247_n1415, Z => mult_21_C247_n66);
   mult_21_C247_U1074 : INVD1 port map( A => N3026, Z => mult_21_C247_n1415);
   mult_21_C247_U1073 : EXOR2D1 port map( A1 => N3025, A2 => N3024, Z => 
                           mult_21_C247_n1450);
   mult_21_C247_U1072 : OAI21D1 port map( A1 => N3023, A2 => N3022, B => 
                           mult_21_C247_n1413, Z => mult_21_C247_n58);
   mult_21_C247_U1071 : INVD1 port map( A => N3024, Z => mult_21_C247_n1413);
   mult_21_C247_U1070 : EXOR2D1 port map( A1 => N3023, A2 => N3022, Z => 
                           mult_21_C247_n1449);
   mult_21_C247_U1069 : OAI21D1 port map( A1 => N3021, A2 => N3020, B => 
                           mult_21_C247_n1411, Z => mult_21_C247_n50);
   mult_21_C247_U1068 : INVD1 port map( A => N3022, Z => mult_21_C247_n1411);
   mult_21_C247_U1067 : EXOR2D1 port map( A1 => N3021, A2 => N3020, Z => 
                           mult_21_C247_n1448);
   mult_21_C247_U1066 : OAI21D1 port map( A1 => N3018, A2 => N3019, B => 
                           mult_21_C247_n1409, Z => mult_21_C247_n42);
   mult_21_C247_U1065 : INVD1 port map( A => N3020, Z => mult_21_C247_n1409);
   mult_21_C247_U1064 : EXOR2D1 port map( A1 => N3019, A2 => N3018, Z => 
                           mult_21_C247_n1447);
   mult_21_C247_U1063 : INVD1 port map( A => N3018, Z => mult_21_C247_n1407);
   mult_21_C247_U1062 : INVD1 port map( A => N3016, Z => mult_21_C247_n1405);
   mult_21_C247_U1061 : INVD1 port map( A => N3206, Z => mult_21_C247_n1386);
   mult_21_C247_U1060 : INVD1 port map( A => N3014, Z => mult_21_C247_n1403);
   mult_21_C247_U1059 : INVD1 port map( A => N3012, Z => mult_21_C247_n1401);
   mult_21_C247_U1058 : INVD1 port map( A => N3205, Z => mult_21_C247_n1388);
   mult_21_C247_U1057 : INVD1 port map( A => N3204, Z => mult_21_C247_n1391);
   mult_21_C247_U1056 : INVD1 port map( A => N3201, Z => mult_21_C247_n1397);
   mult_21_C247_U1055 : INVD1 port map( A => N3202, Z => mult_21_C247_n1395);
   mult_21_C247_U1054 : INVD1 port map( A => N3203, Z => mult_21_C247_n1393);
   mult_21_C247_U1053 : EXNOR2D1 port map( A1 => N3011, A2 => N3010, Z => 
                           mult_21_C247_n1383);
   mult_21_C247_U1052 : INVD1 port map( A => N3010, Z => mult_21_C247_n1398);
   mult_21_C247_U1051 : INVD1 port map( A => mult_21_C247_n939, Z => 
                           mult_21_C247_n1426);
   mult_21_C247_U1050 : INVD1 port map( A => mult_21_C247_n940, Z => 
                           mult_21_C247_n1425);
   mult_21_C247_U1049 : INVD1 port map( A => mult_21_C247_n941, Z => 
                           mult_21_C247_n1422);
   mult_21_C247_U1048 : INVD1 port map( A => mult_21_C247_n942, Z => 
                           mult_21_C247_n1420);
   mult_21_C247_U1047 : INVD1 port map( A => mult_21_C247_n943, Z => 
                           mult_21_C247_n1418);
   mult_21_C247_U1046 : INVD1 port map( A => mult_21_C247_n944, Z => 
                           mult_21_C247_n1416);
   mult_21_C247_U1045 : INVD1 port map( A => mult_21_C247_n945, Z => 
                           mult_21_C247_n1414);
   mult_21_C247_U1044 : INVD1 port map( A => mult_21_C247_n946, Z => 
                           mult_21_C247_n1412);
   mult_21_C247_U1043 : INVD1 port map( A => mult_21_C247_n947, Z => 
                           mult_21_C247_n1410);
   mult_21_C247_U1042 : INVD1 port map( A => mult_21_C247_n948, Z => 
                           mult_21_C247_n1408);
   mult_21_C247_U1041 : INVD1 port map( A => mult_21_C247_n949, Z => 
                           mult_21_C247_n1406);
   mult_21_C247_U1040 : INVD1 port map( A => mult_21_C247_n950, Z => 
                           mult_21_C247_n1404);
   mult_21_C247_U1039 : INVD1 port map( A => mult_21_C247_n951, Z => 
                           mult_21_C247_n1402);
   mult_21_C247_U1038 : INVD1 port map( A => mult_21_C247_n952, Z => 
                           mult_21_C247_n1400);
   mult_21_C247_U1037 : INVD1 port map( A => mult_21_C247_n1388, Z => 
                           mult_21_C247_n1387);
   mult_21_C247_U1036 : INVD1 port map( A => mult_21_C247_n1386, Z => 
                           mult_21_C247_n1385);
   mult_21_C247_U1035 : INVD1 port map( A => mult_21_C247_n953, Z => 
                           mult_21_C247_n1399);
   mult_21_C247_U1034 : INVD1 port map( A => mult_21_C247_n1391, Z => 
                           mult_21_C247_n1390);
   mult_21_C247_U1033 : INVD1 port map( A => mult_21_C247_n1391, Z => 
                           mult_21_C247_n1389);
   mult_21_C247_U1032 : INVD1 port map( A => mult_21_C247_n1397, Z => 
                           mult_21_C247_n1396);
   mult_21_C247_U1031 : INVD1 port map( A => mult_21_C247_n1395, Z => 
                           mult_21_C247_n1394);
   mult_21_C247_U1030 : INVD1 port map( A => mult_21_C247_n1393, Z => 
                           mult_21_C247_n1392);
   mult_21_C247_U1029 : INVD1 port map( A => mult_21_C247_n1383, Z => 
                           mult_21_C247_n1384);
   mult_21_C247_U1028 : OAI21D1 port map( A1 => N3017, A2 => N3016, B => 
                           mult_21_C247_n1407, Z => mult_21_C247_n1382);
   mult_21_C247_U1027 : OAI21D1 port map( A1 => N3015, A2 => N3014, B => 
                           mult_21_C247_n1405, Z => mult_21_C247_n1381);
   mult_21_C247_U1026 : OAI21D1 port map( A1 => N3013, A2 => N3012, B => 
                           mult_21_C247_n1403, Z => mult_21_C247_n1380);
   mult_21_C247_U1025 : OAI21D1 port map( A1 => N3011, A2 => N3010, B => 
                           mult_21_C247_n1401, Z => mult_21_C247_n1379);
   mult_21_C247_U1024 : NAN2D1 port map( A1 => N3009, A2 => mult_21_C247_n1398,
                           Z => mult_21_C247_n1378);
   mult_21_C247_U1023 : EXOR2D1 port map( A1 => N3017, A2 => N3016, Z => 
                           mult_21_C247_n1377);
   mult_21_C247_U1022 : EXOR2D1 port map( A1 => N3015, A2 => N3014, Z => 
                           mult_21_C247_n1376);
   mult_21_C247_U1021 : EXOR2D1 port map( A1 => N3013, A2 => N3012, Z => 
                           mult_21_C247_n1375);
   mult_21_C247_U954 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n923, Z => 
                           mult_21_C247_n1226);
   mult_21_C247_U952 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n922, Z => 
                           mult_21_C247_n1225);
   mult_21_C247_U950 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n921, Z => 
                           mult_21_C247_n1224);
   mult_21_C247_U948 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n920, Z => 
                           mult_21_C247_n1223);
   mult_21_C247_U946 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n919, Z => 
                           mult_21_C247_n1222);
   mult_21_C247_U944 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n918, Z => 
                           mult_21_C247_n1221);
   mult_21_C247_U942 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n917, Z => 
                           mult_21_C247_n1220);
   mult_21_C247_U940 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n916, Z => 
                           mult_21_C247_n1219);
   mult_21_C247_U938 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n915, Z => 
                           mult_21_C247_n1218);
   mult_21_C247_U936 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n914, Z => 
                           mult_21_C247_n1217);
   mult_21_C247_U934 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n913, Z => 
                           mult_21_C247_n1216);
   mult_21_C247_U932 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n912, Z => 
                           mult_21_C247_n1215);
   mult_21_C247_U930 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n911, Z => 
                           mult_21_C247_n1214);
   mult_21_C247_U928 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n910, Z => 
                           mult_21_C247_n1213);
   mult_21_C247_U926 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n909, Z => 
                           mult_21_C247_n1212);
   mult_21_C247_U924 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n908, Z => 
                           mult_21_C247_n1211);
   mult_21_C247_U922 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n907, Z => 
                           mult_21_C247_n1210);
   mult_21_C247_U920 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n906, Z => 
                           mult_21_C247_n1209);
   mult_21_C247_U918 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n905, Z => 
                           mult_21_C247_n1208);
   mult_21_C247_U916 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n904, Z => 
                           mult_21_C247_n1207);
   mult_21_C247_U914 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n903, Z => 
                           mult_21_C247_n1206);
   mult_21_C247_U912 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n902, Z => 
                           mult_21_C247_n1205);
   mult_21_C247_U910 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n901, Z => 
                           mult_21_C247_n1204);
   mult_21_C247_U908 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n900, Z => 
                           mult_21_C247_n1203);
   mult_21_C247_U906 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n899, Z => 
                           mult_21_C247_n1202);
   mult_21_C247_U904 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n898, Z => 
                           mult_21_C247_n1201);
   mult_21_C247_U902 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n897, Z => 
                           mult_21_C247_n1200);
   mult_21_C247_U900 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n896, Z => 
                           mult_21_C247_n1199);
   mult_21_C247_U898 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n895, Z => 
                           mult_21_C247_n1198);
   mult_21_C247_U896 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n894, Z => 
                           mult_21_C247_n1197);
   mult_21_C247_U894 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n893, Z => 
                           mult_21_C247_n1196);
   mult_21_C247_U892 : MUXB2DL port map( A0 => mult_21_C247_n1378, A1 => 
                           mult_21_C247_n1398, SL => mult_21_C247_n892, Z => 
                           mult_21_C247_n1195);
   mult_21_C247_U889 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n891, Z => 
                           mult_21_C247_n1194);
   mult_21_C247_U887 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n890, Z => 
                           mult_21_C247_n1193);
   mult_21_C247_U885 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n889, Z => 
                           mult_21_C247_n1192);
   mult_21_C247_U883 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n888, Z => 
                           mult_21_C247_n1191);
   mult_21_C247_U881 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n887, Z => 
                           mult_21_C247_n1190);
   mult_21_C247_U879 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n886, Z => 
                           mult_21_C247_n1189);
   mult_21_C247_U877 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n885, Z => 
                           mult_21_C247_n1188);
   mult_21_C247_U875 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n884, Z => 
                           mult_21_C247_n1187);
   mult_21_C247_U873 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n883, Z => 
                           mult_21_C247_n1186);
   mult_21_C247_U871 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n882, Z => 
                           mult_21_C247_n1185);
   mult_21_C247_U869 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n881, Z => 
                           mult_21_C247_n1184);
   mult_21_C247_U867 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n880, Z => 
                           mult_21_C247_n1183);
   mult_21_C247_U865 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n879, Z => 
                           mult_21_C247_n1182);
   mult_21_C247_U863 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n878, Z => 
                           mult_21_C247_n1181);
   mult_21_C247_U861 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n877, Z => 
                           mult_21_C247_n1180);
   mult_21_C247_U859 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n876, Z => 
                           mult_21_C247_n1179);
   mult_21_C247_U857 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n875, Z => 
                           mult_21_C247_n1178);
   mult_21_C247_U855 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n874, Z => 
                           mult_21_C247_n1177);
   mult_21_C247_U853 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n873, Z => 
                           mult_21_C247_n1176);
   mult_21_C247_U851 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n872, Z => 
                           mult_21_C247_n1175);
   mult_21_C247_U849 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n871, Z => 
                           mult_21_C247_n1174);
   mult_21_C247_U847 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n870, Z => 
                           mult_21_C247_n1173);
   mult_21_C247_U845 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n869, Z => 
                           mult_21_C247_n1172);
   mult_21_C247_U843 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n868, Z => 
                           mult_21_C247_n1171);
   mult_21_C247_U841 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n867, Z => 
                           mult_21_C247_n1170);
   mult_21_C247_U839 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n866, Z => 
                           mult_21_C247_n1169);
   mult_21_C247_U837 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n865, Z => 
                           mult_21_C247_n1168);
   mult_21_C247_U835 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n864, Z => 
                           mult_21_C247_n1167);
   mult_21_C247_U833 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n863, Z => 
                           mult_21_C247_n1166);
   mult_21_C247_U831 : MUXB2DL port map( A0 => mult_21_C247_n1379, A1 => 
                           mult_21_C247_n1399, SL => mult_21_C247_n862, Z => 
                           mult_21_C247_n1165);
   mult_21_C247_U828 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n861, Z => 
                           mult_21_C247_n1164);
   mult_21_C247_U826 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n860, Z => 
                           mult_21_C247_n1163);
   mult_21_C247_U824 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n859, Z => 
                           mult_21_C247_n1162);
   mult_21_C247_U822 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n858, Z => 
                           mult_21_C247_n1161);
   mult_21_C247_U820 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n857, Z => 
                           mult_21_C247_n1160);
   mult_21_C247_U818 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n856, Z => 
                           mult_21_C247_n1159);
   mult_21_C247_U816 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n855, Z => 
                           mult_21_C247_n1158);
   mult_21_C247_U814 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n854, Z => 
                           mult_21_C247_n1157);
   mult_21_C247_U812 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n853, Z => 
                           mult_21_C247_n1156);
   mult_21_C247_U810 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n852, Z => 
                           mult_21_C247_n1155);
   mult_21_C247_U808 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n851, Z => 
                           mult_21_C247_n1154);
   mult_21_C247_U806 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n850, Z => 
                           mult_21_C247_n1153);
   mult_21_C247_U804 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n849, Z => 
                           mult_21_C247_n1152);
   mult_21_C247_U802 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n848, Z => 
                           mult_21_C247_n1151);
   mult_21_C247_U800 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n847, Z => 
                           mult_21_C247_n1150);
   mult_21_C247_U798 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n846, Z => 
                           mult_21_C247_n1149);
   mult_21_C247_U796 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n845, Z => 
                           mult_21_C247_n1148);
   mult_21_C247_U794 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n844, Z => 
                           mult_21_C247_n1147);
   mult_21_C247_U792 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n843, Z => 
                           mult_21_C247_n1146);
   mult_21_C247_U790 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n842, Z => 
                           mult_21_C247_n1145);
   mult_21_C247_U788 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n841, Z => 
                           mult_21_C247_n1144);
   mult_21_C247_U786 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n840, Z => 
                           mult_21_C247_n1143);
   mult_21_C247_U784 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n839, Z => 
                           mult_21_C247_n1142);
   mult_21_C247_U782 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n838, Z => 
                           mult_21_C247_n1141);
   mult_21_C247_U780 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n837, Z => 
                           mult_21_C247_n1140);
   mult_21_C247_U778 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n836, Z => 
                           mult_21_C247_n1139);
   mult_21_C247_U776 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n835, Z => 
                           mult_21_C247_n1138);
   mult_21_C247_U774 : MUXB2DL port map( A0 => mult_21_C247_n1380, A1 => 
                           mult_21_C247_n1400, SL => mult_21_C247_n834, Z => 
                           mult_21_C247_n1137);
   mult_21_C247_U771 : MUXB2DL port map( A0 => mult_21_C247_n1381, A1 => 
                           mult_21_C247_n1402, SL => mult_21_C247_n833, Z => 
                           mult_21_C247_n1136);
   mult_21_C247_U769 : MUXB2DL port map( A0 => mult_21_C247_n1381, A1 => 
                           mult_21_C247_n1402, SL => mult_21_C247_n832, Z => 
                           mult_21_C247_n1135);
   mult_21_C247_U767 : MUXB2DL port map( A0 => mult_21_C247_n1381, A1 => 
                           mult_21_C247_n1402, SL => mult_21_C247_n831, Z => 
                           mult_21_C247_n1134);
   mult_21_C247_U765 : MUXB2DL port map( A0 => mult_21_C247_n1381, A1 => 
                           mult_21_C247_n1402, SL => mult_21_C247_n830, Z => 
                           mult_21_C247_n1133);
   mult_21_C247_U763 : MUXB2DL port map( A0 => mult_21_C247_n1381, A1 => 
                           mult_21_C247_n1402, SL => mult_21_C247_n829, Z => 
                           mult_21_C247_n1132);
   mult_21_C247_U761 : MUXB2DL port map( A0 => mult_21_C247_n1381, A1 => 
                           mult_21_C247_n1402, SL => mult_21_C247_n828, Z => 
                           mult_21_C247_n1131);
   mult_21_C247_U759 : MUXB2DL port map( A0 => mult_21_C247_n1381, A1 => 
                           mult_21_C247_n1402, SL => mult_21_C247_n827, Z => 
                           mult_21_C247_n1130);
   mult_21_C247_U757 : MUXB2DL port map( A0 => mult_21_C247_n1381, A1 => 
                           mult_21_C247_n1402, SL => mult_21_C247_n826, Z => 
                           mult_21_C247_n1129);
   mult_21_C247_U755 : MUXB2DL port map( A0 => mult_21_C247_n1381, A1 => 
                           mult_21_C247_n1402, SL => mult_21_C247_n825, Z => 
                           mult_21_C247_n1128);
   mult_21_C247_U753 : MUXB2DL port map( A0 => mult_21_C247_n1381, A1 => 
                           mult_21_C247_n1402, SL => mult_21_C247_n824, Z => 
                           mult_21_C247_n1127);
   mult_21_C247_U751 : MUXB2DL port map( A0 => mult_21_C247_n1381, A1 => 
                           mult_21_C247_n1402, SL => mult_21_C247_n823, Z => 
                           mult_21_C247_n1126);
   mult_21_C247_U749 : MUXB2DL port map( A0 => mult_21_C247_n1381, A1 => 
                           mult_21_C247_n1402, SL => mult_21_C247_n822, Z => 
                           mult_21_C247_n1125);
   mult_21_C247_U747 : MUXB2DL port map( A0 => mult_21_C247_n1381, A1 => 
                           mult_21_C247_n1402, SL => mult_21_C247_n821, Z => 
                           mult_21_C247_n1124);
   mult_21_C247_U745 : MUXB2DL port map( A0 => mult_21_C247_n1381, A1 => 
                           mult_21_C247_n1402, SL => mult_21_C247_n820, Z => 
                           mult_21_C247_n1123);
   mult_21_C247_U743 : MUXB2DL port map( A0 => mult_21_C247_n1381, A1 => 
                           mult_21_C247_n1402, SL => mult_21_C247_n819, Z => 
                           mult_21_C247_n1122);
   mult_21_C247_U741 : MUXB2DL port map( A0 => mult_21_C247_n1381, A1 => 
                           mult_21_C247_n1402, SL => mult_21_C247_n818, Z => 
                           mult_21_C247_n1121);
   mult_21_C247_U739 : MUXB2DL port map( A0 => mult_21_C247_n1381, A1 => 
                           mult_21_C247_n1402, SL => mult_21_C247_n817, Z => 
                           mult_21_C247_n1120);
   mult_21_C247_U737 : MUXB2DL port map( A0 => mult_21_C247_n1381, A1 => 
                           mult_21_C247_n1402, SL => mult_21_C247_n816, Z => 
                           mult_21_C247_n1119);
   mult_21_C247_U735 : MUXB2DL port map( A0 => mult_21_C247_n1381, A1 => 
                           mult_21_C247_n1402, SL => mult_21_C247_n815, Z => 
                           mult_21_C247_n1118);
   mult_21_C247_U733 : MUXB2DL port map( A0 => mult_21_C247_n1381, A1 => 
                           mult_21_C247_n1402, SL => mult_21_C247_n814, Z => 
                           mult_21_C247_n1117);
   mult_21_C247_U731 : MUXB2DL port map( A0 => mult_21_C247_n1381, A1 => 
                           mult_21_C247_n1402, SL => mult_21_C247_n813, Z => 
                           mult_21_C247_n1116);
   mult_21_C247_U729 : MUXB2DL port map( A0 => mult_21_C247_n1381, A1 => 
                           mult_21_C247_n1402, SL => mult_21_C247_n812, Z => 
                           mult_21_C247_n1115);
   mult_21_C247_U727 : MUXB2DL port map( A0 => mult_21_C247_n1381, A1 => 
                           mult_21_C247_n1402, SL => mult_21_C247_n811, Z => 
                           mult_21_C247_n1114);
   mult_21_C247_U725 : MUXB2DL port map( A0 => mult_21_C247_n1381, A1 => 
                           mult_21_C247_n1402, SL => mult_21_C247_n810, Z => 
                           mult_21_C247_n1113);
   mult_21_C247_U723 : MUXB2DL port map( A0 => mult_21_C247_n1381, A1 => 
                           mult_21_C247_n1402, SL => mult_21_C247_n809, Z => 
                           mult_21_C247_n1112);
   mult_21_C247_U721 : MUXB2DL port map( A0 => mult_21_C247_n1381, A1 => 
                           mult_21_C247_n1402, SL => mult_21_C247_n808, Z => 
                           mult_21_C247_n1111);
   mult_21_C247_U718 : MUXB2DL port map( A0 => mult_21_C247_n1382, A1 => 
                           mult_21_C247_n1404, SL => mult_21_C247_n807, Z => 
                           mult_21_C247_n1110);
   mult_21_C247_U716 : MUXB2DL port map( A0 => mult_21_C247_n1382, A1 => 
                           mult_21_C247_n1404, SL => mult_21_C247_n806, Z => 
                           mult_21_C247_n1109);
   mult_21_C247_U714 : MUXB2DL port map( A0 => mult_21_C247_n1382, A1 => 
                           mult_21_C247_n1404, SL => mult_21_C247_n805, Z => 
                           mult_21_C247_n1108);
   mult_21_C247_U712 : MUXB2DL port map( A0 => mult_21_C247_n1382, A1 => 
                           mult_21_C247_n1404, SL => mult_21_C247_n804, Z => 
                           mult_21_C247_n1107);
   mult_21_C247_U710 : MUXB2DL port map( A0 => mult_21_C247_n1382, A1 => 
                           mult_21_C247_n1404, SL => mult_21_C247_n803, Z => 
                           mult_21_C247_n1106);
   mult_21_C247_U708 : MUXB2DL port map( A0 => mult_21_C247_n1382, A1 => 
                           mult_21_C247_n1404, SL => mult_21_C247_n802, Z => 
                           mult_21_C247_n1105);
   mult_21_C247_U706 : MUXB2DL port map( A0 => mult_21_C247_n1382, A1 => 
                           mult_21_C247_n1404, SL => mult_21_C247_n801, Z => 
                           mult_21_C247_n1104);
   mult_21_C247_U704 : MUXB2DL port map( A0 => mult_21_C247_n1382, A1 => 
                           mult_21_C247_n1404, SL => mult_21_C247_n800, Z => 
                           mult_21_C247_n1103);
   mult_21_C247_U702 : MUXB2DL port map( A0 => mult_21_C247_n1382, A1 => 
                           mult_21_C247_n1404, SL => mult_21_C247_n799, Z => 
                           mult_21_C247_n1102);
   mult_21_C247_U700 : MUXB2DL port map( A0 => mult_21_C247_n1382, A1 => 
                           mult_21_C247_n1404, SL => mult_21_C247_n798, Z => 
                           mult_21_C247_n1101);
   mult_21_C247_U698 : MUXB2DL port map( A0 => mult_21_C247_n1382, A1 => 
                           mult_21_C247_n1404, SL => mult_21_C247_n797, Z => 
                           mult_21_C247_n1100);
   mult_21_C247_U696 : MUXB2DL port map( A0 => mult_21_C247_n1382, A1 => 
                           mult_21_C247_n1404, SL => mult_21_C247_n796, Z => 
                           mult_21_C247_n1099);
   mult_21_C247_U694 : MUXB2DL port map( A0 => mult_21_C247_n1382, A1 => 
                           mult_21_C247_n1404, SL => mult_21_C247_n795, Z => 
                           mult_21_C247_n1098);
   mult_21_C247_U692 : MUXB2DL port map( A0 => mult_21_C247_n1382, A1 => 
                           mult_21_C247_n1404, SL => mult_21_C247_n794, Z => 
                           mult_21_C247_n1097);
   mult_21_C247_U690 : MUXB2DL port map( A0 => mult_21_C247_n1382, A1 => 
                           mult_21_C247_n1404, SL => mult_21_C247_n793, Z => 
                           mult_21_C247_n1096);
   mult_21_C247_U688 : MUXB2DL port map( A0 => mult_21_C247_n1382, A1 => 
                           mult_21_C247_n1404, SL => mult_21_C247_n792, Z => 
                           mult_21_C247_n1095);
   mult_21_C247_U686 : MUXB2DL port map( A0 => mult_21_C247_n1382, A1 => 
                           mult_21_C247_n1404, SL => mult_21_C247_n791, Z => 
                           mult_21_C247_n1094);
   mult_21_C247_U684 : MUXB2DL port map( A0 => mult_21_C247_n1382, A1 => 
                           mult_21_C247_n1404, SL => mult_21_C247_n790, Z => 
                           mult_21_C247_n1093);
   mult_21_C247_U682 : MUXB2DL port map( A0 => mult_21_C247_n1382, A1 => 
                           mult_21_C247_n1404, SL => mult_21_C247_n789, Z => 
                           mult_21_C247_n1092);
   mult_21_C247_U680 : MUXB2DL port map( A0 => mult_21_C247_n1382, A1 => 
                           mult_21_C247_n1404, SL => mult_21_C247_n788, Z => 
                           mult_21_C247_n1091);
   mult_21_C247_U678 : MUXB2DL port map( A0 => mult_21_C247_n1382, A1 => 
                           mult_21_C247_n1404, SL => mult_21_C247_n787, Z => 
                           mult_21_C247_n1090);
   mult_21_C247_U676 : MUXB2DL port map( A0 => mult_21_C247_n1382, A1 => 
                           mult_21_C247_n1404, SL => mult_21_C247_n786, Z => 
                           mult_21_C247_n1089);
   mult_21_C247_U674 : MUXB2DL port map( A0 => mult_21_C247_n1382, A1 => 
                           mult_21_C247_n1404, SL => mult_21_C247_n785, Z => 
                           mult_21_C247_n1088);
   mult_21_C247_U672 : MUXB2DL port map( A0 => mult_21_C247_n1382, A1 => 
                           mult_21_C247_n1404, SL => mult_21_C247_n784, Z => 
                           mult_21_C247_n1087);
   mult_21_C247_U669 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n1406, SL => mult_21_C247_n783, Z => 
                           mult_21_C247_n1086);
   mult_21_C247_U667 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n1406, SL => mult_21_C247_n782, Z => 
                           mult_21_C247_n1085);
   mult_21_C247_U665 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n1406, SL => mult_21_C247_n781, Z => 
                           mult_21_C247_n1084);
   mult_21_C247_U663 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n1406, SL => mult_21_C247_n780, Z => 
                           mult_21_C247_n1083);
   mult_21_C247_U661 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n1406, SL => mult_21_C247_n779, Z => 
                           mult_21_C247_n1082);
   mult_21_C247_U659 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n1406, SL => mult_21_C247_n778, Z => 
                           mult_21_C247_n1081);
   mult_21_C247_U657 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n1406, SL => mult_21_C247_n777, Z => 
                           mult_21_C247_n1080);
   mult_21_C247_U655 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n1406, SL => mult_21_C247_n776, Z => 
                           mult_21_C247_n1079);
   mult_21_C247_U653 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n1406, SL => mult_21_C247_n775, Z => 
                           mult_21_C247_n1078);
   mult_21_C247_U651 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n1406, SL => mult_21_C247_n774, Z => 
                           mult_21_C247_n1077);
   mult_21_C247_U649 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n1406, SL => mult_21_C247_n773, Z => 
                           mult_21_C247_n1076);
   mult_21_C247_U647 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n1406, SL => mult_21_C247_n772, Z => 
                           mult_21_C247_n1075);
   mult_21_C247_U645 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n1406, SL => mult_21_C247_n771, Z => 
                           mult_21_C247_n1074);
   mult_21_C247_U643 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n1406, SL => mult_21_C247_n770, Z => 
                           mult_21_C247_n1073);
   mult_21_C247_U641 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n1406, SL => mult_21_C247_n769, Z => 
                           mult_21_C247_n1072);
   mult_21_C247_U639 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n1406, SL => mult_21_C247_n768, Z => 
                           mult_21_C247_n1071);
   mult_21_C247_U637 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n1406, SL => mult_21_C247_n767, Z => 
                           mult_21_C247_n1070);
   mult_21_C247_U635 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n1406, SL => mult_21_C247_n766, Z => 
                           mult_21_C247_n1069);
   mult_21_C247_U633 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n1406, SL => mult_21_C247_n765, Z => 
                           mult_21_C247_n1068);
   mult_21_C247_U631 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n1406, SL => mult_21_C247_n764, Z => 
                           mult_21_C247_n1067);
   mult_21_C247_U629 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n1406, SL => mult_21_C247_n763, Z => 
                           mult_21_C247_n1066);
   mult_21_C247_U627 : MUXB2DL port map( A0 => mult_21_C247_n42, A1 => 
                           mult_21_C247_n1406, SL => mult_21_C247_n762, Z => 
                           mult_21_C247_n1065);
   mult_21_C247_U624 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n1408, SL => mult_21_C247_n761, Z => 
                           mult_21_C247_n1064);
   mult_21_C247_U622 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n1408, SL => mult_21_C247_n760, Z => 
                           mult_21_C247_n1063);
   mult_21_C247_U620 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n1408, SL => mult_21_C247_n759, Z => 
                           mult_21_C247_n1062);
   mult_21_C247_U618 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n1408, SL => mult_21_C247_n758, Z => 
                           mult_21_C247_n1061);
   mult_21_C247_U616 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n1408, SL => mult_21_C247_n757, Z => 
                           mult_21_C247_n1060);
   mult_21_C247_U614 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n1408, SL => mult_21_C247_n756, Z => 
                           mult_21_C247_n1059);
   mult_21_C247_U612 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n1408, SL => mult_21_C247_n755, Z => 
                           mult_21_C247_n1058);
   mult_21_C247_U610 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n1408, SL => mult_21_C247_n754, Z => 
                           mult_21_C247_n1057);
   mult_21_C247_U608 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n1408, SL => mult_21_C247_n753, Z => 
                           mult_21_C247_n1056);
   mult_21_C247_U606 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n1408, SL => mult_21_C247_n752, Z => 
                           mult_21_C247_n1055);
   mult_21_C247_U604 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n1408, SL => mult_21_C247_n751, Z => 
                           mult_21_C247_n1054);
   mult_21_C247_U602 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n1408, SL => mult_21_C247_n750, Z => 
                           mult_21_C247_n1053);
   mult_21_C247_U600 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n1408, SL => mult_21_C247_n749, Z => 
                           mult_21_C247_n1052);
   mult_21_C247_U598 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n1408, SL => mult_21_C247_n748, Z => 
                           mult_21_C247_n1051);
   mult_21_C247_U596 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n1408, SL => mult_21_C247_n747, Z => 
                           mult_21_C247_n1050);
   mult_21_C247_U594 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n1408, SL => mult_21_C247_n746, Z => 
                           mult_21_C247_n1049);
   mult_21_C247_U592 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n1408, SL => mult_21_C247_n745, Z => 
                           mult_21_C247_n1048);
   mult_21_C247_U590 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n1408, SL => mult_21_C247_n744, Z => 
                           mult_21_C247_n1047);
   mult_21_C247_U588 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n1408, SL => mult_21_C247_n743, Z => 
                           mult_21_C247_n1046);
   mult_21_C247_U586 : MUXB2DL port map( A0 => mult_21_C247_n50, A1 => 
                           mult_21_C247_n1408, SL => mult_21_C247_n742, Z => 
                           mult_21_C247_n1045);
   mult_21_C247_U583 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n1410, SL => mult_21_C247_n741, Z => 
                           mult_21_C247_n1044);
   mult_21_C247_U581 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n1410, SL => mult_21_C247_n740, Z => 
                           mult_21_C247_n1043);
   mult_21_C247_U579 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n1410, SL => mult_21_C247_n739, Z => 
                           mult_21_C247_n1042);
   mult_21_C247_U577 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n1410, SL => mult_21_C247_n738, Z => 
                           mult_21_C247_n1041);
   mult_21_C247_U575 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n1410, SL => mult_21_C247_n737, Z => 
                           mult_21_C247_n1040);
   mult_21_C247_U573 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n1410, SL => mult_21_C247_n736, Z => 
                           mult_21_C247_n1039);
   mult_21_C247_U571 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n1410, SL => mult_21_C247_n735, Z => 
                           mult_21_C247_n1038);
   mult_21_C247_U569 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n1410, SL => mult_21_C247_n734, Z => 
                           mult_21_C247_n1037);
   mult_21_C247_U567 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n1410, SL => mult_21_C247_n733, Z => 
                           mult_21_C247_n1036);
   mult_21_C247_U565 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n1410, SL => mult_21_C247_n732, Z => 
                           mult_21_C247_n1035);
   mult_21_C247_U563 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n1410, SL => mult_21_C247_n731, Z => 
                           mult_21_C247_n1034);
   mult_21_C247_U561 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n1410, SL => mult_21_C247_n730, Z => 
                           mult_21_C247_n1033);
   mult_21_C247_U559 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n1410, SL => mult_21_C247_n729, Z => 
                           mult_21_C247_n1032);
   mult_21_C247_U557 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n1410, SL => mult_21_C247_n728, Z => 
                           mult_21_C247_n1031);
   mult_21_C247_U555 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n1410, SL => mult_21_C247_n727, Z => 
                           mult_21_C247_n1030);
   mult_21_C247_U553 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n1410, SL => mult_21_C247_n726, Z => 
                           mult_21_C247_n1029);
   mult_21_C247_U551 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n1410, SL => mult_21_C247_n725, Z => 
                           mult_21_C247_n1028);
   mult_21_C247_U549 : MUXB2DL port map( A0 => mult_21_C247_n58, A1 => 
                           mult_21_C247_n1410, SL => mult_21_C247_n724, Z => 
                           mult_21_C247_n1027);
   mult_21_C247_U546 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n1412, SL => mult_21_C247_n723, Z => 
                           mult_21_C247_n1026);
   mult_21_C247_U544 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n1412, SL => mult_21_C247_n722, Z => 
                           mult_21_C247_n1025);
   mult_21_C247_U542 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n1412, SL => mult_21_C247_n721, Z => 
                           mult_21_C247_n1024);
   mult_21_C247_U540 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n1412, SL => mult_21_C247_n720, Z => 
                           mult_21_C247_n1023);
   mult_21_C247_U538 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n1412, SL => mult_21_C247_n719, Z => 
                           mult_21_C247_n1022);
   mult_21_C247_U536 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n1412, SL => mult_21_C247_n718, Z => 
                           mult_21_C247_n1021);
   mult_21_C247_U534 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n1412, SL => mult_21_C247_n717, Z => 
                           mult_21_C247_n1020);
   mult_21_C247_U532 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n1412, SL => mult_21_C247_n716, Z => 
                           mult_21_C247_n1019);
   mult_21_C247_U530 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n1412, SL => mult_21_C247_n715, Z => 
                           mult_21_C247_n1018);
   mult_21_C247_U528 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n1412, SL => mult_21_C247_n714, Z => 
                           mult_21_C247_n1017);
   mult_21_C247_U526 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n1412, SL => mult_21_C247_n713, Z => 
                           mult_21_C247_n1016);
   mult_21_C247_U524 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n1412, SL => mult_21_C247_n712, Z => 
                           mult_21_C247_n1015);
   mult_21_C247_U522 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n1412, SL => mult_21_C247_n711, Z => 
                           mult_21_C247_n1014);
   mult_21_C247_U520 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n1412, SL => mult_21_C247_n710, Z => 
                           mult_21_C247_n1013);
   mult_21_C247_U518 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n1412, SL => mult_21_C247_n709, Z => 
                           mult_21_C247_n1012);
   mult_21_C247_U516 : MUXB2DL port map( A0 => mult_21_C247_n66, A1 => 
                           mult_21_C247_n1412, SL => mult_21_C247_n708, Z => 
                           mult_21_C247_n1011);
   mult_21_C247_U513 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n1414, SL => mult_21_C247_n707, Z => 
                           mult_21_C247_n1010);
   mult_21_C247_U511 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n1414, SL => mult_21_C247_n706, Z => 
                           mult_21_C247_n1009);
   mult_21_C247_U509 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n1414, SL => mult_21_C247_n705, Z => 
                           mult_21_C247_n1008);
   mult_21_C247_U507 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n1414, SL => mult_21_C247_n704, Z => 
                           mult_21_C247_n1007);
   mult_21_C247_U505 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n1414, SL => mult_21_C247_n703, Z => 
                           mult_21_C247_n1006);
   mult_21_C247_U503 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n1414, SL => mult_21_C247_n702, Z => 
                           mult_21_C247_n1005);
   mult_21_C247_U501 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n1414, SL => mult_21_C247_n701, Z => 
                           mult_21_C247_n1004);
   mult_21_C247_U499 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n1414, SL => mult_21_C247_n700, Z => 
                           mult_21_C247_n1003);
   mult_21_C247_U497 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n1414, SL => mult_21_C247_n699, Z => 
                           mult_21_C247_n1002);
   mult_21_C247_U495 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n1414, SL => mult_21_C247_n698, Z => 
                           mult_21_C247_n1001);
   mult_21_C247_U493 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n1414, SL => mult_21_C247_n697, Z => 
                           mult_21_C247_n1000);
   mult_21_C247_U491 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n1414, SL => mult_21_C247_n696, Z => 
                           mult_21_C247_n999);
   mult_21_C247_U489 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n1414, SL => mult_21_C247_n695, Z => 
                           mult_21_C247_n998);
   mult_21_C247_U487 : MUXB2DL port map( A0 => mult_21_C247_n73, A1 => 
                           mult_21_C247_n1414, SL => mult_21_C247_n694, Z => 
                           mult_21_C247_n997);
   mult_21_C247_U484 : MUXB2DL port map( A0 => mult_21_C247_n80, A1 => 
                           mult_21_C247_n1416, SL => mult_21_C247_n693, Z => 
                           mult_21_C247_n996);
   mult_21_C247_U482 : MUXB2DL port map( A0 => mult_21_C247_n80, A1 => 
                           mult_21_C247_n1416, SL => mult_21_C247_n692, Z => 
                           mult_21_C247_n995);
   mult_21_C247_U480 : MUXB2DL port map( A0 => mult_21_C247_n80, A1 => 
                           mult_21_C247_n1416, SL => mult_21_C247_n691, Z => 
                           mult_21_C247_n994);
   mult_21_C247_U478 : MUXB2DL port map( A0 => mult_21_C247_n80, A1 => 
                           mult_21_C247_n1416, SL => mult_21_C247_n690, Z => 
                           mult_21_C247_n993);
   mult_21_C247_U476 : MUXB2DL port map( A0 => mult_21_C247_n80, A1 => 
                           mult_21_C247_n1416, SL => mult_21_C247_n689, Z => 
                           mult_21_C247_n992);
   mult_21_C247_U474 : MUXB2DL port map( A0 => mult_21_C247_n80, A1 => 
                           mult_21_C247_n1416, SL => mult_21_C247_n688, Z => 
                           mult_21_C247_n991);
   mult_21_C247_U472 : MUXB2DL port map( A0 => mult_21_C247_n80, A1 => 
                           mult_21_C247_n1416, SL => mult_21_C247_n687, Z => 
                           mult_21_C247_n990);
   mult_21_C247_U470 : MUXB2DL port map( A0 => mult_21_C247_n80, A1 => 
                           mult_21_C247_n1416, SL => mult_21_C247_n686, Z => 
                           mult_21_C247_n989);
   mult_21_C247_U468 : MUXB2DL port map( A0 => mult_21_C247_n80, A1 => 
                           mult_21_C247_n1416, SL => mult_21_C247_n685, Z => 
                           mult_21_C247_n988);
   mult_21_C247_U466 : MUXB2DL port map( A0 => mult_21_C247_n80, A1 => 
                           mult_21_C247_n1416, SL => mult_21_C247_n684, Z => 
                           mult_21_C247_n987);
   mult_21_C247_U464 : MUXB2DL port map( A0 => mult_21_C247_n80, A1 => 
                           mult_21_C247_n1416, SL => mult_21_C247_n683, Z => 
                           mult_21_C247_n986);
   mult_21_C247_U462 : MUXB2DL port map( A0 => mult_21_C247_n80, A1 => 
                           mult_21_C247_n1416, SL => mult_21_C247_n682, Z => 
                           mult_21_C247_n985);
   mult_21_C247_U459 : MUXB2DL port map( A0 => mult_21_C247_n84, A1 => 
                           mult_21_C247_n1418, SL => mult_21_C247_n681, Z => 
                           mult_21_C247_n984);
   mult_21_C247_U457 : MUXB2DL port map( A0 => mult_21_C247_n84, A1 => 
                           mult_21_C247_n1418, SL => mult_21_C247_n680, Z => 
                           mult_21_C247_n983);
   mult_21_C247_U455 : MUXB2DL port map( A0 => mult_21_C247_n84, A1 => 
                           mult_21_C247_n1418, SL => mult_21_C247_n679, Z => 
                           mult_21_C247_n982);
   mult_21_C247_U453 : MUXB2DL port map( A0 => mult_21_C247_n84, A1 => 
                           mult_21_C247_n1418, SL => mult_21_C247_n678, Z => 
                           mult_21_C247_n981);
   mult_21_C247_U451 : MUXB2DL port map( A0 => mult_21_C247_n84, A1 => 
                           mult_21_C247_n1418, SL => mult_21_C247_n677, Z => 
                           mult_21_C247_n980);
   mult_21_C247_U449 : MUXB2DL port map( A0 => mult_21_C247_n84, A1 => 
                           mult_21_C247_n1418, SL => mult_21_C247_n676, Z => 
                           mult_21_C247_n979);
   mult_21_C247_U447 : MUXB2DL port map( A0 => mult_21_C247_n84, A1 => 
                           mult_21_C247_n1418, SL => mult_21_C247_n675, Z => 
                           mult_21_C247_n978);
   mult_21_C247_U445 : MUXB2DL port map( A0 => mult_21_C247_n84, A1 => 
                           mult_21_C247_n1418, SL => mult_21_C247_n674, Z => 
                           mult_21_C247_n977);
   mult_21_C247_U443 : MUXB2DL port map( A0 => mult_21_C247_n84, A1 => 
                           mult_21_C247_n1418, SL => mult_21_C247_n673, Z => 
                           mult_21_C247_n976);
   mult_21_C247_U441 : MUXB2DL port map( A0 => mult_21_C247_n84, A1 => 
                           mult_21_C247_n1418, SL => mult_21_C247_n672, Z => 
                           mult_21_C247_n975);
   mult_21_C247_U438 : MUXB2DL port map( A0 => mult_21_C247_n89, A1 => 
                           mult_21_C247_n1420, SL => mult_21_C247_n671, Z => 
                           mult_21_C247_n974);
   mult_21_C247_U436 : MUXB2DL port map( A0 => mult_21_C247_n89, A1 => 
                           mult_21_C247_n1420, SL => mult_21_C247_n670, Z => 
                           mult_21_C247_n973);
   mult_21_C247_U434 : MUXB2DL port map( A0 => mult_21_C247_n89, A1 => 
                           mult_21_C247_n1420, SL => mult_21_C247_n669, Z => 
                           mult_21_C247_n972);
   mult_21_C247_U432 : MUXB2DL port map( A0 => mult_21_C247_n89, A1 => 
                           mult_21_C247_n1420, SL => mult_21_C247_n668, Z => 
                           mult_21_C247_n971);
   mult_21_C247_U430 : MUXB2DL port map( A0 => mult_21_C247_n89, A1 => 
                           mult_21_C247_n1420, SL => mult_21_C247_n667, Z => 
                           mult_21_C247_n970);
   mult_21_C247_U428 : MUXB2DL port map( A0 => mult_21_C247_n89, A1 => 
                           mult_21_C247_n1420, SL => mult_21_C247_n666, Z => 
                           mult_21_C247_n969);
   mult_21_C247_U426 : MUXB2DL port map( A0 => mult_21_C247_n89, A1 => 
                           mult_21_C247_n1420, SL => mult_21_C247_n665, Z => 
                           mult_21_C247_n968);
   mult_21_C247_U424 : MUXB2DL port map( A0 => mult_21_C247_n89, A1 => 
                           mult_21_C247_n1420, SL => mult_21_C247_n664, Z => 
                           mult_21_C247_n967);
   mult_21_C247_U421 : MUXB2DL port map( A0 => mult_21_C247_n94, A1 => 
                           mult_21_C247_n1422, SL => mult_21_C247_n663, Z => 
                           mult_21_C247_n966);
   mult_21_C247_U419 : MUXB2DL port map( A0 => mult_21_C247_n94, A1 => 
                           mult_21_C247_n1422, SL => mult_21_C247_n662, Z => 
                           mult_21_C247_n965);
   mult_21_C247_U417 : MUXB2DL port map( A0 => mult_21_C247_n94, A1 => 
                           mult_21_C247_n1422, SL => mult_21_C247_n661, Z => 
                           mult_21_C247_n964);
   mult_21_C247_U415 : MUXB2DL port map( A0 => mult_21_C247_n94, A1 => 
                           mult_21_C247_n1422, SL => mult_21_C247_n660, Z => 
                           mult_21_C247_n963);
   mult_21_C247_U413 : MUXB2DL port map( A0 => mult_21_C247_n94, A1 => 
                           mult_21_C247_n1422, SL => mult_21_C247_n659, Z => 
                           mult_21_C247_n962);
   mult_21_C247_U411 : MUXB2DL port map( A0 => mult_21_C247_n94, A1 => 
                           mult_21_C247_n1422, SL => mult_21_C247_n658, Z => 
                           mult_21_C247_n961);
   mult_21_C247_U408 : MUXB2DL port map( A0 => mult_21_C247_n99, A1 => 
                           mult_21_C247_n1425, SL => mult_21_C247_n657, Z => 
                           mult_21_C247_n960);
   mult_21_C247_U406 : MUXB2DL port map( A0 => mult_21_C247_n99, A1 => 
                           mult_21_C247_n1425, SL => mult_21_C247_n656, Z => 
                           mult_21_C247_n959);
   mult_21_C247_U404 : MUXB2DL port map( A0 => mult_21_C247_n99, A1 => 
                           mult_21_C247_n1425, SL => mult_21_C247_n655, Z => 
                           mult_21_C247_n958);
   mult_21_C247_U402 : MUXB2DL port map( A0 => mult_21_C247_n99, A1 => 
                           mult_21_C247_n1425, SL => mult_21_C247_n654, Z => 
                           mult_21_C247_n957);
   mult_21_C247_U399 : MUXB2DL port map( A0 => mult_21_C247_n104, A1 => 
                           mult_21_C247_n1426, SL => mult_21_C247_n653, Z => 
                           mult_21_C247_n956);
   mult_21_C247_U397 : MUXB2DL port map( A0 => mult_21_C247_n104, A1 => 
                           mult_21_C247_n1426, SL => mult_21_C247_n652, Z => 
                           mult_21_C247_n955);
   mult_21_C247_U395 : ADHALFDL port map( A => mult_21_C247_n1224, B => 
                           mult_21_C247_n953, CO => mult_21_C247_n650, S => 
                           mult_21_C247_n651);
   mult_21_C247_U394 : ADHALFDL port map( A => mult_21_C247_n650, B => 
                           mult_21_C247_n1223, CO => mult_21_C247_n648, S => 
                           mult_21_C247_n649);
   mult_21_C247_U393 : ADHALFDL port map( A => mult_21_C247_n1222, B => 
                           mult_21_C247_n952, CO => mult_21_C247_n646, S => 
                           mult_21_C247_n647);
   mult_21_C247_U392 : ADFULD1 port map( A => mult_21_C247_n1192, B => 
                           mult_21_C247_n1164, CI => mult_21_C247_n647, CO => 
                           mult_21_C247_n644, S => mult_21_C247_n645);
   mult_21_C247_U391 : ADHALFDL port map( A => mult_21_C247_n646, B => 
                           mult_21_C247_n1221, CO => mult_21_C247_n642, S => 
                           mult_21_C247_n643);
   mult_21_C247_U390 : ADFULD1 port map( A => mult_21_C247_n1163, B => 
                           mult_21_C247_n1191, CI => mult_21_C247_n643, CO => 
                           mult_21_C247_n640, S => mult_21_C247_n641);
   mult_21_C247_U389 : ADHALFDL port map( A => mult_21_C247_n1220, B => 
                           mult_21_C247_n951, CO => mult_21_C247_n638, S => 
                           mult_21_C247_n639);
   mult_21_C247_U388 : ADFULD1 port map( A => mult_21_C247_n1190, B => 
                           mult_21_C247_n1136, CI => mult_21_C247_n1162, CO => 
                           mult_21_C247_n636, S => mult_21_C247_n637);
   mult_21_C247_U387 : ADFULD1 port map( A => mult_21_C247_n642, B => 
                           mult_21_C247_n639, CI => mult_21_C247_n637, CO => 
                           mult_21_C247_n634, S => mult_21_C247_n635);
   mult_21_C247_U386 : ADHALFDL port map( A => mult_21_C247_n638, B => 
                           mult_21_C247_n1219, CO => mult_21_C247_n632, S => 
                           mult_21_C247_n633);
   mult_21_C247_U385 : ADFULD1 port map( A => mult_21_C247_n1135, B => 
                           mult_21_C247_n1189, CI => mult_21_C247_n1161, CO => 
                           mult_21_C247_n630, S => mult_21_C247_n631);
   mult_21_C247_U384 : ADFULD1 port map( A => mult_21_C247_n636, B => 
                           mult_21_C247_n633, CI => mult_21_C247_n631, CO => 
                           mult_21_C247_n628, S => mult_21_C247_n629);
   mult_21_C247_U383 : ADHALFDL port map( A => mult_21_C247_n1218, B => 
                           mult_21_C247_n950, CO => mult_21_C247_n626, S => 
                           mult_21_C247_n627);
   mult_21_C247_U382 : ADFULD1 port map( A => mult_21_C247_n1188, B => 
                           mult_21_C247_n1110, CI => mult_21_C247_n1134, CO => 
                           mult_21_C247_n624, S => mult_21_C247_n625);
   mult_21_C247_U381 : ADFULD1 port map( A => mult_21_C247_n627, B => 
                           mult_21_C247_n1160, CI => mult_21_C247_n632, CO => 
                           mult_21_C247_n622, S => mult_21_C247_n623);
   mult_21_C247_U380 : ADFULD1 port map( A => mult_21_C247_n625, B => 
                           mult_21_C247_n630, CI => mult_21_C247_n623, CO => 
                           mult_21_C247_n620, S => mult_21_C247_n621);
   mult_21_C247_U379 : ADHALFDL port map( A => mult_21_C247_n626, B => 
                           mult_21_C247_n1217, CO => mult_21_C247_n618, S => 
                           mult_21_C247_n619);
   mult_21_C247_U378 : ADFULD1 port map( A => mult_21_C247_n1109, B => 
                           mult_21_C247_n1133, CI => mult_21_C247_n1159, CO => 
                           mult_21_C247_n616, S => mult_21_C247_n617);
   mult_21_C247_U377 : ADFULD1 port map( A => mult_21_C247_n619, B => 
                           mult_21_C247_n1187, CI => mult_21_C247_n624, CO => 
                           mult_21_C247_n614, S => mult_21_C247_n615);
   mult_21_C247_U376 : ADFULD1 port map( A => mult_21_C247_n617, B => 
                           mult_21_C247_n622, CI => mult_21_C247_n615, CO => 
                           mult_21_C247_n612, S => mult_21_C247_n613);
   mult_21_C247_U375 : ADHALFDL port map( A => mult_21_C247_n1216, B => 
                           mult_21_C247_n949, CO => mult_21_C247_n610, S => 
                           mult_21_C247_n611);
   mult_21_C247_U374 : ADFULD1 port map( A => mult_21_C247_n1132, B => 
                           mult_21_C247_n1086, CI => mult_21_C247_n1186, CO => 
                           mult_21_C247_n608, S => mult_21_C247_n609);
   mult_21_C247_U373 : ADFULD1 port map( A => mult_21_C247_n1108, B => 
                           mult_21_C247_n1158, CI => mult_21_C247_n611, CO => 
                           mult_21_C247_n606, S => mult_21_C247_n607);
   mult_21_C247_U372 : ADFULD1 port map( A => mult_21_C247_n616, B => 
                           mult_21_C247_n618, CI => mult_21_C247_n609, CO => 
                           mult_21_C247_n604, S => mult_21_C247_n605);
   mult_21_C247_U371 : ADFULD1 port map( A => mult_21_C247_n614, B => 
                           mult_21_C247_n607, CI => mult_21_C247_n605, CO => 
                           mult_21_C247_n602, S => mult_21_C247_n603);
   mult_21_C247_U370 : ADHALFDL port map( A => mult_21_C247_n610, B => 
                           mult_21_C247_n1215, CO => mult_21_C247_n600, S => 
                           mult_21_C247_n601);
   mult_21_C247_U369 : ADFULD1 port map( A => mult_21_C247_n1085, B => 
                           mult_21_C247_n1131, CI => mult_21_C247_n1185, CO => 
                           mult_21_C247_n598, S => mult_21_C247_n599);
   mult_21_C247_U368 : ADFULD1 port map( A => mult_21_C247_n1107, B => 
                           mult_21_C247_n1157, CI => mult_21_C247_n601, CO => 
                           mult_21_C247_n596, S => mult_21_C247_n597);
   mult_21_C247_U367 : ADFULD1 port map( A => mult_21_C247_n606, B => 
                           mult_21_C247_n608, CI => mult_21_C247_n599, CO => 
                           mult_21_C247_n594, S => mult_21_C247_n595);
   mult_21_C247_U366 : ADFULD1 port map( A => mult_21_C247_n604, B => 
                           mult_21_C247_n597, CI => mult_21_C247_n595, CO => 
                           mult_21_C247_n592, S => mult_21_C247_n593);
   mult_21_C247_U365 : ADHALFDL port map( A => mult_21_C247_n1214, B => 
                           mult_21_C247_n948, CO => mult_21_C247_n590, S => 
                           mult_21_C247_n591);
   mult_21_C247_U364 : ADFULD1 port map( A => mult_21_C247_n1130, B => 
                           mult_21_C247_n1064, CI => mult_21_C247_n1184, CO => 
                           mult_21_C247_n588, S => mult_21_C247_n589);
   mult_21_C247_U363 : ADFULD1 port map( A => mult_21_C247_n1084, B => 
                           mult_21_C247_n1156, CI => mult_21_C247_n591, CO => 
                           mult_21_C247_n586, S => mult_21_C247_n587);
   mult_21_C247_U362 : ADFULD1 port map( A => mult_21_C247_n600, B => 
                           mult_21_C247_n1106, CI => mult_21_C247_n598, CO => 
                           mult_21_C247_n584, S => mult_21_C247_n585);
   mult_21_C247_U361 : ADFULD1 port map( A => mult_21_C247_n587, B => 
                           mult_21_C247_n589, CI => mult_21_C247_n596, CO => 
                           mult_21_C247_n582, S => mult_21_C247_n583);
   mult_21_C247_U360 : ADFULD1 port map( A => mult_21_C247_n585, B => 
                           mult_21_C247_n594, CI => mult_21_C247_n583, CO => 
                           mult_21_C247_n580, S => mult_21_C247_n581);
   mult_21_C247_U359 : ADHALFDL port map( A => mult_21_C247_n590, B => 
                           mult_21_C247_n1213, CO => mult_21_C247_n578, S => 
                           mult_21_C247_n579);
   mult_21_C247_U358 : ADFULD1 port map( A => mult_21_C247_n1183, B => 
                           mult_21_C247_n1105, CI => mult_21_C247_n1155, CO => 
                           mult_21_C247_n576, S => mult_21_C247_n577);
   mult_21_C247_U357 : ADFULD1 port map( A => mult_21_C247_n1063, B => 
                           mult_21_C247_n1129, CI => mult_21_C247_n1083, CO => 
                           mult_21_C247_n574, S => mult_21_C247_n575);
   mult_21_C247_U356 : ADFULD1 port map( A => mult_21_C247_n588, B => 
                           mult_21_C247_n579, CI => mult_21_C247_n586, CO => 
                           mult_21_C247_n572, S => mult_21_C247_n573);
   mult_21_C247_U355 : ADFULD1 port map( A => mult_21_C247_n577, B => 
                           mult_21_C247_n575, CI => mult_21_C247_n584, CO => 
                           mult_21_C247_n570, S => mult_21_C247_n571);
   mult_21_C247_U354 : ADFULD1 port map( A => mult_21_C247_n582, B => 
                           mult_21_C247_n573, CI => mult_21_C247_n571, CO => 
                           mult_21_C247_n568, S => mult_21_C247_n569);
   mult_21_C247_U353 : ADHALFDL port map( A => mult_21_C247_n1212, B => 
                           mult_21_C247_n947, CO => mult_21_C247_n566, S => 
                           mult_21_C247_n567);
   mult_21_C247_U352 : ADFULD1 port map( A => mult_21_C247_n1104, B => 
                           mult_21_C247_n1044, CI => mult_21_C247_n1182, CO => 
                           mult_21_C247_n564, S => mult_21_C247_n565);
   mult_21_C247_U351 : ADFULD1 port map( A => mult_21_C247_n1154, B => 
                           mult_21_C247_n1082, CI => mult_21_C247_n567, CO => 
                           mult_21_C247_n562, S => mult_21_C247_n563);
   mult_21_C247_U350 : ADFULD1 port map( A => mult_21_C247_n1062, B => 
                           mult_21_C247_n1128, CI => mult_21_C247_n578, CO => 
                           mult_21_C247_n560, S => mult_21_C247_n561);
   mult_21_C247_U349 : ADFULD1 port map( A => mult_21_C247_n574, B => 
                           mult_21_C247_n576, CI => mult_21_C247_n565, CO => 
                           mult_21_C247_n558, S => mult_21_C247_n559);
   mult_21_C247_U348 : ADFULD1 port map( A => mult_21_C247_n561, B => 
                           mult_21_C247_n563, CI => mult_21_C247_n572, CO => 
                           mult_21_C247_n556, S => mult_21_C247_n557);
   mult_21_C247_U347 : ADFULD1 port map( A => mult_21_C247_n570, B => 
                           mult_21_C247_n559, CI => mult_21_C247_n557, CO => 
                           mult_21_C247_n554, S => mult_21_C247_n555);
   mult_21_C247_U346 : ADHALFDL port map( A => mult_21_C247_n566, B => 
                           mult_21_C247_n1211, CO => mult_21_C247_n552, S => 
                           mult_21_C247_n553);
   mult_21_C247_U345 : ADFULD1 port map( A => mult_21_C247_n1043, B => 
                           mult_21_C247_n1103, CI => mult_21_C247_n1061, CO => 
                           mult_21_C247_n550, S => mult_21_C247_n551);
   mult_21_C247_U344 : ADFULD1 port map( A => mult_21_C247_n1181, B => 
                           mult_21_C247_n1081, CI => mult_21_C247_n1127, CO => 
                           mult_21_C247_n548, S => mult_21_C247_n549);
   mult_21_C247_U343 : ADFULD1 port map( A => mult_21_C247_n553, B => 
                           mult_21_C247_n1153, CI => mult_21_C247_n564, CO => 
                           mult_21_C247_n546, S => mult_21_C247_n547);
   mult_21_C247_U342 : ADFULD1 port map( A => mult_21_C247_n560, B => 
                           mult_21_C247_n562, CI => mult_21_C247_n549, CO => 
                           mult_21_C247_n544, S => mult_21_C247_n545);
   mult_21_C247_U341 : ADFULD1 port map( A => mult_21_C247_n547, B => 
                           mult_21_C247_n551, CI => mult_21_C247_n558, CO => 
                           mult_21_C247_n542, S => mult_21_C247_n543);
   mult_21_C247_U340 : ADFULD1 port map( A => mult_21_C247_n556, B => 
                           mult_21_C247_n545, CI => mult_21_C247_n543, CO => 
                           mult_21_C247_n540, S => mult_21_C247_n541);
   mult_21_C247_U339 : ADHALFDL port map( A => mult_21_C247_n1210, B => 
                           mult_21_C247_n946, CO => mult_21_C247_n538, S => 
                           mult_21_C247_n539);
   mult_21_C247_U338 : ADFULD1 port map( A => mult_21_C247_n1102, B => 
                           mult_21_C247_n1026, CI => mult_21_C247_n1180, CO => 
                           mult_21_C247_n536, S => mult_21_C247_n537);
   mult_21_C247_U337 : ADFULD1 port map( A => mult_21_C247_n1042, B => 
                           mult_21_C247_n1060, CI => mult_21_C247_n539, CO => 
                           mult_21_C247_n534, S => mult_21_C247_n535);
   mult_21_C247_U336 : ADFULD1 port map( A => mult_21_C247_n1080, B => 
                           mult_21_C247_n1152, CI => mult_21_C247_n1126, CO => 
                           mult_21_C247_n532, S => mult_21_C247_n533);
   mult_21_C247_U335 : ADFULD1 port map( A => mult_21_C247_n550, B => 
                           mult_21_C247_n552, CI => mult_21_C247_n548, CO => 
                           mult_21_C247_n530, S => mult_21_C247_n531);
   mult_21_C247_U334 : ADFULD1 port map( A => mult_21_C247_n533, B => 
                           mult_21_C247_n537, CI => mult_21_C247_n535, CO => 
                           mult_21_C247_n528, S => mult_21_C247_n529);
   mult_21_C247_U333 : ADFULD1 port map( A => mult_21_C247_n544, B => 
                           mult_21_C247_n546, CI => mult_21_C247_n531, CO => 
                           mult_21_C247_n526, S => mult_21_C247_n527);
   mult_21_C247_U332 : ADFULD1 port map( A => mult_21_C247_n542, B => 
                           mult_21_C247_n529, CI => mult_21_C247_n527, CO => 
                           mult_21_C247_n524, S => mult_21_C247_n525);
   mult_21_C247_U331 : ADHALFDL port map( A => mult_21_C247_n538, B => 
                           mult_21_C247_n1209, CO => mult_21_C247_n522, S => 
                           mult_21_C247_n523);
   mult_21_C247_U330 : ADFULD1 port map( A => mult_21_C247_n1179, B => 
                           mult_21_C247_n1079, CI => mult_21_C247_n1151, CO => 
                           mult_21_C247_n520, S => mult_21_C247_n521);
   mult_21_C247_U329 : ADFULD1 port map( A => mult_21_C247_n1025, B => 
                           mult_21_C247_n1041, CI => mult_21_C247_n1059, CO => 
                           mult_21_C247_n518, S => mult_21_C247_n519);
   mult_21_C247_U328 : ADFULD1 port map( A => mult_21_C247_n1101, B => 
                           mult_21_C247_n1125, CI => mult_21_C247_n523, CO => 
                           mult_21_C247_n516, S => mult_21_C247_n517);
   mult_21_C247_U327 : ADFULD1 port map( A => mult_21_C247_n534, B => 
                           mult_21_C247_n536, CI => mult_21_C247_n532, CO => 
                           mult_21_C247_n514, S => mult_21_C247_n515);
   mult_21_C247_U326 : ADFULD1 port map( A => mult_21_C247_n521, B => 
                           mult_21_C247_n519, CI => mult_21_C247_n517, CO => 
                           mult_21_C247_n512, S => mult_21_C247_n513);
   mult_21_C247_U325 : ADFULD1 port map( A => mult_21_C247_n528, B => 
                           mult_21_C247_n530, CI => mult_21_C247_n515, CO => 
                           mult_21_C247_n510, S => mult_21_C247_n511);
   mult_21_C247_U324 : ADFULD1 port map( A => mult_21_C247_n526, B => 
                           mult_21_C247_n513, CI => mult_21_C247_n511, CO => 
                           mult_21_C247_n508, S => mult_21_C247_n509);
   mult_21_C247_U323 : ADHALFDL port map( A => mult_21_C247_n1208, B => 
                           mult_21_C247_n945, CO => mult_21_C247_n506, S => 
                           mult_21_C247_n507);
   mult_21_C247_U322 : ADFULD1 port map( A => mult_21_C247_n1078, B => 
                           mult_21_C247_n1010, CI => mult_21_C247_n1024, CO => 
                           mult_21_C247_n504, S => mult_21_C247_n505);
   mult_21_C247_U321 : ADFULD1 port map( A => mult_21_C247_n1178, B => 
                           mult_21_C247_n1100, CI => mult_21_C247_n507, CO => 
                           mult_21_C247_n502, S => mult_21_C247_n503);
   mult_21_C247_U320 : ADFULD1 port map( A => mult_21_C247_n1040, B => 
                           mult_21_C247_n1150, CI => mult_21_C247_n1058, CO => 
                           mult_21_C247_n500, S => mult_21_C247_n501);
   mult_21_C247_U319 : ADFULD1 port map( A => mult_21_C247_n522, B => 
                           mult_21_C247_n1124, CI => mult_21_C247_n520, CO => 
                           mult_21_C247_n498, S => mult_21_C247_n499);
   mult_21_C247_U318 : ADFULD1 port map( A => mult_21_C247_n505, B => 
                           mult_21_C247_n518, CI => mult_21_C247_n501, CO => 
                           mult_21_C247_n496, S => mult_21_C247_n497);
   mult_21_C247_U317 : ADFULD1 port map( A => mult_21_C247_n516, B => 
                           mult_21_C247_n503, CI => mult_21_C247_n514, CO => 
                           mult_21_C247_n494, S => mult_21_C247_n495);
   mult_21_C247_U316 : ADFULD1 port map( A => mult_21_C247_n497, B => 
                           mult_21_C247_n499, CI => mult_21_C247_n512, CO => 
                           mult_21_C247_n492, S => mult_21_C247_n493);
   mult_21_C247_U315 : ADFULD1 port map( A => mult_21_C247_n510, B => 
                           mult_21_C247_n495, CI => mult_21_C247_n493, CO => 
                           mult_21_C247_n490, S => mult_21_C247_n491);
   mult_21_C247_U314 : ADHALFDL port map( A => mult_21_C247_n506, B => 
                           mult_21_C247_n1207, CO => mult_21_C247_n488, S => 
                           mult_21_C247_n489);
   mult_21_C247_U313 : ADFULD1 port map( A => mult_21_C247_n1009, B => 
                           mult_21_C247_n1077, CI => mult_21_C247_n1023, CO => 
                           mult_21_C247_n486, S => mult_21_C247_n487);
   mult_21_C247_U312 : ADFULD1 port map( A => mult_21_C247_n1177, B => 
                           mult_21_C247_n1099, CI => mult_21_C247_n1039, CO => 
                           mult_21_C247_n484, S => mult_21_C247_n485);
   mult_21_C247_U311 : ADFULD1 port map( A => mult_21_C247_n1057, B => 
                           mult_21_C247_n1149, CI => mult_21_C247_n1123, CO => 
                           mult_21_C247_n482, S => mult_21_C247_n483);
   mult_21_C247_U310 : ADFULD1 port map( A => mult_21_C247_n504, B => 
                           mult_21_C247_n489, CI => mult_21_C247_n502, CO => 
                           mult_21_C247_n480, S => mult_21_C247_n481);
   mult_21_C247_U309 : ADFULD1 port map( A => mult_21_C247_n483, B => 
                           mult_21_C247_n500, CI => mult_21_C247_n485, CO => 
                           mult_21_C247_n478, S => mult_21_C247_n479);
   mult_21_C247_U308 : ADFULD1 port map( A => mult_21_C247_n498, B => 
                           mult_21_C247_n487, CI => mult_21_C247_n496, CO => 
                           mult_21_C247_n476, S => mult_21_C247_n477);
   mult_21_C247_U307 : ADFULD1 port map( A => mult_21_C247_n479, B => 
                           mult_21_C247_n481, CI => mult_21_C247_n494, CO => 
                           mult_21_C247_n474, S => mult_21_C247_n475);
   mult_21_C247_U306 : ADFULD1 port map( A => mult_21_C247_n492, B => 
                           mult_21_C247_n477, CI => mult_21_C247_n475, CO => 
                           mult_21_C247_n472, S => mult_21_C247_n473);
   mult_21_C247_U305 : ADHALFDL port map( A => mult_21_C247_n1206, B => 
                           mult_21_C247_n944, CO => mult_21_C247_n470, S => 
                           mult_21_C247_n471);
   mult_21_C247_U304 : ADFULD1 port map( A => mult_21_C247_n1076, B => 
                           mult_21_C247_n996, CI => mult_21_C247_n1176, CO => 
                           mult_21_C247_n468, S => mult_21_C247_n469);
   mult_21_C247_U303 : ADFULD1 port map( A => mult_21_C247_n1008, B => 
                           mult_21_C247_n1038, CI => mult_21_C247_n471, CO => 
                           mult_21_C247_n466, S => mult_21_C247_n467);
   mult_21_C247_U302 : ADFULD1 port map( A => mult_21_C247_n1022, B => 
                           mult_21_C247_n1148, CI => mult_21_C247_n1056, CO => 
                           mult_21_C247_n464, S => mult_21_C247_n465);
   mult_21_C247_U301 : ADFULD1 port map( A => mult_21_C247_n1098, B => 
                           mult_21_C247_n1122, CI => mult_21_C247_n488, CO => 
                           mult_21_C247_n462, S => mult_21_C247_n463);
   mult_21_C247_U300 : ADFULD1 port map( A => mult_21_C247_n482, B => 
                           mult_21_C247_n486, CI => mult_21_C247_n484, CO => 
                           mult_21_C247_n460, S => mult_21_C247_n461);
   mult_21_C247_U299 : ADFULD1 port map( A => mult_21_C247_n465, B => 
                           mult_21_C247_n469, CI => mult_21_C247_n467, CO => 
                           mult_21_C247_n458, S => mult_21_C247_n459);
   mult_21_C247_U298 : ADFULD1 port map( A => mult_21_C247_n480, B => 
                           mult_21_C247_n463, CI => mult_21_C247_n478, CO => 
                           mult_21_C247_n456, S => mult_21_C247_n457);
   mult_21_C247_U297 : ADFULD1 port map( A => mult_21_C247_n459, B => 
                           mult_21_C247_n461, CI => mult_21_C247_n476, CO => 
                           mult_21_C247_n454, S => mult_21_C247_n455);
   mult_21_C247_U296 : ADFULD1 port map( A => mult_21_C247_n474, B => 
                           mult_21_C247_n457, CI => mult_21_C247_n455, CO => 
                           mult_21_C247_n452, S => mult_21_C247_n453);
   mult_21_C247_U295 : ADHALFDL port map( A => mult_21_C247_n470, B => 
                           mult_21_C247_n1205, CO => mult_21_C247_n450, S => 
                           mult_21_C247_n451);
   mult_21_C247_U294 : ADFULD1 port map( A => mult_21_C247_n1175, B => 
                           mult_21_C247_n1055, CI => mult_21_C247_n1147, CO => 
                           mult_21_C247_n448, S => mult_21_C247_n449);
   mult_21_C247_U293 : ADFULD1 port map( A => mult_21_C247_n1121, B => 
                           mult_21_C247_n1021, CI => mult_21_C247_n1097, CO => 
                           mult_21_C247_n446, S => mult_21_C247_n447);
   mult_21_C247_U292 : ADFULD1 port map( A => mult_21_C247_n995, B => 
                           mult_21_C247_n1075, CI => mult_21_C247_n1007, CO => 
                           mult_21_C247_n444, S => mult_21_C247_n445);
   mult_21_C247_U291 : ADFULD1 port map( A => mult_21_C247_n451, B => 
                           mult_21_C247_n1037, CI => mult_21_C247_n468, CO => 
                           mult_21_C247_n442, S => mult_21_C247_n443);
   mult_21_C247_U290 : ADFULD1 port map( A => mult_21_C247_n464, B => 
                           mult_21_C247_n466, CI => mult_21_C247_n462, CO => 
                           mult_21_C247_n440, S => mult_21_C247_n441);
   mult_21_C247_U289 : ADFULD1 port map( A => mult_21_C247_n449, B => 
                           mult_21_C247_n445, CI => mult_21_C247_n447, CO => 
                           mult_21_C247_n438, S => mult_21_C247_n439);
   mult_21_C247_U288 : ADFULD1 port map( A => mult_21_C247_n443, B => 
                           mult_21_C247_n460, CI => mult_21_C247_n458, CO => 
                           mult_21_C247_n436, S => mult_21_C247_n437);
   mult_21_C247_U287 : ADFULD1 port map( A => mult_21_C247_n439, B => 
                           mult_21_C247_n441, CI => mult_21_C247_n456, CO => 
                           mult_21_C247_n434, S => mult_21_C247_n435);
   mult_21_C247_U286 : ADFULD1 port map( A => mult_21_C247_n454, B => 
                           mult_21_C247_n437, CI => mult_21_C247_n435, CO => 
                           mult_21_C247_n432, S => mult_21_C247_n433);
   mult_21_C247_U285 : ADHALFDL port map( A => mult_21_C247_n1204, B => 
                           mult_21_C247_n943, CO => mult_21_C247_n430, S => 
                           mult_21_C247_n431);
   mult_21_C247_U284 : ADFULD1 port map( A => mult_21_C247_n1054, B => 
                           mult_21_C247_n984, CI => mult_21_C247_n994, CO => 
                           mult_21_C247_n428, S => mult_21_C247_n429);
   mult_21_C247_U283 : ADFULD1 port map( A => mult_21_C247_n1174, B => 
                           mult_21_C247_n1036, CI => mult_21_C247_n431, CO => 
                           mult_21_C247_n426, S => mult_21_C247_n427);
   mult_21_C247_U282 : ADFULD1 port map( A => mult_21_C247_n1006, B => 
                           mult_21_C247_n1146, CI => mult_21_C247_n1020, CO => 
                           mult_21_C247_n424, S => mult_21_C247_n425);
   mult_21_C247_U281 : ADFULD1 port map( A => mult_21_C247_n1074, B => 
                           mult_21_C247_n1120, CI => mult_21_C247_n1096, CO => 
                           mult_21_C247_n422, S => mult_21_C247_n423);
   mult_21_C247_U280 : ADFULD1 port map( A => mult_21_C247_n448, B => 
                           mult_21_C247_n450, CI => mult_21_C247_n446, CO => 
                           mult_21_C247_n420, S => mult_21_C247_n421);
   mult_21_C247_U279 : ADFULD1 port map( A => mult_21_C247_n429, B => 
                           mult_21_C247_n444, CI => mult_21_C247_n423, CO => 
                           mult_21_C247_n418, S => mult_21_C247_n419);
   mult_21_C247_U278 : ADFULD1 port map( A => mult_21_C247_n427, B => 
                           mult_21_C247_n425, CI => mult_21_C247_n442, CO => 
                           mult_21_C247_n416, S => mult_21_C247_n417);
   mult_21_C247_U277 : ADFULD1 port map( A => mult_21_C247_n421, B => 
                           mult_21_C247_n440, CI => mult_21_C247_n438, CO => 
                           mult_21_C247_n414, S => mult_21_C247_n415);
   mult_21_C247_U276 : ADFULD1 port map( A => mult_21_C247_n417, B => 
                           mult_21_C247_n419, CI => mult_21_C247_n436, CO => 
                           mult_21_C247_n412, S => mult_21_C247_n413);
   mult_21_C247_U275 : ADFULD1 port map( A => mult_21_C247_n434, B => 
                           mult_21_C247_n415, CI => mult_21_C247_n413, CO => 
                           mult_21_C247_n410, S => mult_21_C247_n411);
   mult_21_C247_U274 : ADHALFDL port map( A => mult_21_C247_n430, B => 
                           mult_21_C247_n1203, CO => mult_21_C247_n408, S => 
                           mult_21_C247_n409);
   mult_21_C247_U273 : ADFULD1 port map( A => mult_21_C247_n983, B => 
                           mult_21_C247_n1053, CI => mult_21_C247_n993, CO => 
                           mult_21_C247_n406, S => mult_21_C247_n407);
   mult_21_C247_U272 : ADFULD1 port map( A => mult_21_C247_n1173, B => 
                           mult_21_C247_n1035, CI => mult_21_C247_n1145, CO => 
                           mult_21_C247_n404, S => mult_21_C247_n405);
   mult_21_C247_U271 : ADFULD1 port map( A => mult_21_C247_n1005, B => 
                           mult_21_C247_n1119, CI => mult_21_C247_n1019, CO => 
                           mult_21_C247_n402, S => mult_21_C247_n403);
   mult_21_C247_U270 : ADFULD1 port map( A => mult_21_C247_n1073, B => 
                           mult_21_C247_n1095, CI => mult_21_C247_n409, CO => 
                           mult_21_C247_n400, S => mult_21_C247_n401);
   mult_21_C247_U269 : ADFULD1 port map( A => mult_21_C247_n426, B => 
                           mult_21_C247_n428, CI => mult_21_C247_n422, CO => 
                           mult_21_C247_n398, S => mult_21_C247_n399);
   mult_21_C247_U268 : ADFULD1 port map( A => mult_21_C247_n403, B => 
                           mult_21_C247_n424, CI => mult_21_C247_n405, CO => 
                           mult_21_C247_n396, S => mult_21_C247_n397);
   mult_21_C247_U267 : ADFULD1 port map( A => mult_21_C247_n401, B => 
                           mult_21_C247_n407, CI => mult_21_C247_n420, CO => 
                           mult_21_C247_n394, S => mult_21_C247_n395);
   mult_21_C247_U266 : ADFULD1 port map( A => mult_21_C247_n399, B => 
                           mult_21_C247_n418, CI => mult_21_C247_n416, CO => 
                           mult_21_C247_n392, S => mult_21_C247_n393);
   mult_21_C247_U265 : ADFULD1 port map( A => mult_21_C247_n395, B => 
                           mult_21_C247_n397, CI => mult_21_C247_n414, CO => 
                           mult_21_C247_n390, S => mult_21_C247_n391);
   mult_21_C247_U264 : ADFULD1 port map( A => mult_21_C247_n412, B => 
                           mult_21_C247_n393, CI => mult_21_C247_n391, CO => 
                           mult_21_C247_n388, S => mult_21_C247_n389);
   mult_21_C247_U263 : ADHALFDL port map( A => mult_21_C247_n1202, B => 
                           mult_21_C247_n942, CO => mult_21_C247_n386, S => 
                           mult_21_C247_n387);
   mult_21_C247_U262 : ADFULD1 port map( A => mult_21_C247_n1052, B => 
                           mult_21_C247_n974, CI => mult_21_C247_n1172, CO => 
                           mult_21_C247_n384, S => mult_21_C247_n385);
   mult_21_C247_U261 : ADFULD1 port map( A => mult_21_C247_n982, B => 
                           mult_21_C247_n1018, CI => mult_21_C247_n387, CO => 
                           mult_21_C247_n382, S => mult_21_C247_n383);
   mult_21_C247_U260 : ADFULD1 port map( A => mult_21_C247_n992, B => 
                           mult_21_C247_n1144, CI => mult_21_C247_n1118, CO => 
                           mult_21_C247_n380, S => mult_21_C247_n381);
   mult_21_C247_U259 : ADFULD1 port map( A => mult_21_C247_n1004, B => 
                           mult_21_C247_n1094, CI => mult_21_C247_n1034, CO => 
                           mult_21_C247_n378, S => mult_21_C247_n379);
   mult_21_C247_U258 : ADFULD1 port map( A => mult_21_C247_n408, B => 
                           mult_21_C247_n1072, CI => mult_21_C247_n406, CO => 
                           mult_21_C247_n376, S => mult_21_C247_n377);
   mult_21_C247_U257 : ADFULD1 port map( A => mult_21_C247_n402, B => 
                           mult_21_C247_n404, CI => mult_21_C247_n385, CO => 
                           mult_21_C247_n374, S => mult_21_C247_n375);
   mult_21_C247_U256 : ADFULD1 port map( A => mult_21_C247_n383, B => 
                           mult_21_C247_n379, CI => mult_21_C247_n381, CO => 
                           mult_21_C247_n372, S => mult_21_C247_n373);
   mult_21_C247_U255 : ADFULD1 port map( A => mult_21_C247_n398, B => 
                           mult_21_C247_n400, CI => mult_21_C247_n377, CO => 
                           mult_21_C247_n370, S => mult_21_C247_n371);
   mult_21_C247_U254 : ADFULD1 port map( A => mult_21_C247_n375, B => 
                           mult_21_C247_n396, CI => mult_21_C247_n373, CO => 
                           mult_21_C247_n368, S => mult_21_C247_n369);
   mult_21_C247_U253 : ADFULD1 port map( A => mult_21_C247_n371, B => 
                           mult_21_C247_n394, CI => mult_21_C247_n392, CO => 
                           mult_21_C247_n366, S => mult_21_C247_n367);
   mult_21_C247_U252 : ADFULD1 port map( A => mult_21_C247_n390, B => 
                           mult_21_C247_n369, CI => mult_21_C247_n367, CO => 
                           mult_21_C247_n364, S => mult_21_C247_n365);
   mult_21_C247_U251 : ADHALFDL port map( A => mult_21_C247_n386, B => 
                           mult_21_C247_n1201, CO => mult_21_C247_n362, S => 
                           mult_21_C247_n363);
   mult_21_C247_U250 : ADFULD1 port map( A => mult_21_C247_n1171, B => 
                           mult_21_C247_n1051, CI => mult_21_C247_n1143, CO => 
                           mult_21_C247_n360, S => mult_21_C247_n361);
   mult_21_C247_U249 : ADFULD1 port map( A => mult_21_C247_n973, B => 
                           mult_21_C247_n1003, CI => mult_21_C247_n981, CO => 
                           mult_21_C247_n358, S => mult_21_C247_n359);
   mult_21_C247_U248 : ADFULD1 port map( A => mult_21_C247_n991, B => 
                           mult_21_C247_n1117, CI => mult_21_C247_n1017, CO => 
                           mult_21_C247_n356, S => mult_21_C247_n357);
   mult_21_C247_U247 : ADFULD1 port map( A => mult_21_C247_n1033, B => 
                           mult_21_C247_n1093, CI => mult_21_C247_n1071, CO => 
                           mult_21_C247_n354, S => mult_21_C247_n355);
   mult_21_C247_U246 : ADFULD1 port map( A => mult_21_C247_n384, B => 
                           mult_21_C247_n363, CI => mult_21_C247_n382, CO => 
                           mult_21_C247_n352, S => mult_21_C247_n353);
   mult_21_C247_U245 : ADFULD1 port map( A => mult_21_C247_n378, B => 
                           mult_21_C247_n380, CI => mult_21_C247_n355, CO => 
                           mult_21_C247_n350, S => mult_21_C247_n351);
   mult_21_C247_U244 : ADFULD1 port map( A => mult_21_C247_n361, B => 
                           mult_21_C247_n357, CI => mult_21_C247_n359, CO => 
                           mult_21_C247_n348, S => mult_21_C247_n349);
   mult_21_C247_U243 : ADFULD1 port map( A => mult_21_C247_n374, B => 
                           mult_21_C247_n376, CI => mult_21_C247_n353, CO => 
                           mult_21_C247_n346, S => mult_21_C247_n347);
   mult_21_C247_U242 : ADFULD1 port map( A => mult_21_C247_n351, B => 
                           mult_21_C247_n372, CI => mult_21_C247_n349, CO => 
                           mult_21_C247_n344, S => mult_21_C247_n345);
   mult_21_C247_U241 : ADFULD1 port map( A => mult_21_C247_n347, B => 
                           mult_21_C247_n370, CI => mult_21_C247_n368, CO => 
                           mult_21_C247_n342, S => mult_21_C247_n343);
   mult_21_C247_U240 : ADFULD1 port map( A => mult_21_C247_n366, B => 
                           mult_21_C247_n345, CI => mult_21_C247_n343, CO => 
                           mult_21_C247_n340, S => mult_21_C247_n341);
   mult_21_C247_U239 : ADHALFDL port map( A => mult_21_C247_n1200, B => 
                           mult_21_C247_n941, CO => mult_21_C247_n338, S => 
                           mult_21_C247_n339);
   mult_21_C247_U238 : ADFULD1 port map( A => mult_21_C247_n1050, B => 
                           mult_21_C247_n966, CI => mult_21_C247_n972, CO => 
                           mult_21_C247_n336, S => mult_21_C247_n337);
   mult_21_C247_U237 : ADFULD1 port map( A => mult_21_C247_n980, B => 
                           mult_21_C247_n1032, CI => mult_21_C247_n339, CO => 
                           mult_21_C247_n334, S => mult_21_C247_n335);
   mult_21_C247_U236 : ADFULD1 port map( A => mult_21_C247_n990, B => 
                           mult_21_C247_n1170, CI => mult_21_C247_n1002, CO => 
                           mult_21_C247_n332, S => mult_21_C247_n333);
   mult_21_C247_U235 : ADFULD1 port map( A => mult_21_C247_n1016, B => 
                           mult_21_C247_n1142, CI => mult_21_C247_n1070, CO => 
                           mult_21_C247_n330, S => mult_21_C247_n331);
   mult_21_C247_U234 : ADFULD1 port map( A => mult_21_C247_n1092, B => 
                           mult_21_C247_n1116, CI => mult_21_C247_n362, CO => 
                           mult_21_C247_n328, S => mult_21_C247_n329);
   mult_21_C247_U233 : ADFULD1 port map( A => mult_21_C247_n354, B => 
                           mult_21_C247_n360, CI => mult_21_C247_n356, CO => 
                           mult_21_C247_n326, S => mult_21_C247_n327);
   mult_21_C247_U232 : ADFULD1 port map( A => mult_21_C247_n337, B => 
                           mult_21_C247_n358, CI => mult_21_C247_n331, CO => 
                           mult_21_C247_n324, S => mult_21_C247_n325);
   mult_21_C247_U231 : ADFULD1 port map( A => mult_21_C247_n333, B => 
                           mult_21_C247_n335, CI => mult_21_C247_n329, CO => 
                           mult_21_C247_n322, S => mult_21_C247_n323);
   mult_21_C247_U230 : ADFULD1 port map( A => mult_21_C247_n350, B => 
                           mult_21_C247_n352, CI => mult_21_C247_n348, CO => 
                           mult_21_C247_n320, S => mult_21_C247_n321);
   mult_21_C247_U229 : ADFULD1 port map( A => mult_21_C247_n325, B => 
                           mult_21_C247_n327, CI => mult_21_C247_n323, CO => 
                           mult_21_C247_n318, S => mult_21_C247_n319);
   mult_21_C247_U228 : ADFULD1 port map( A => mult_21_C247_n344, B => 
                           mult_21_C247_n346, CI => mult_21_C247_n321, CO => 
                           mult_21_C247_n316, S => mult_21_C247_n317);
   mult_21_C247_U227 : ADFULD1 port map( A => mult_21_C247_n342, B => 
                           mult_21_C247_n319, CI => mult_21_C247_n317, CO => 
                           mult_21_C247_n314, S => mult_21_C247_n315);
   mult_21_C247_U226 : ADHALFDL port map( A => mult_21_C247_n338, B => 
                           mult_21_C247_n1199, CO => mult_21_C247_n312, S => 
                           mult_21_C247_n313);
   mult_21_C247_U225 : ADFULD1 port map( A => mult_21_C247_n965, B => 
                           mult_21_C247_n1031, CI => mult_21_C247_n971, CO => 
                           mult_21_C247_n310, S => mult_21_C247_n311);
   mult_21_C247_U224 : ADFULD1 port map( A => mult_21_C247_n979, B => 
                           mult_21_C247_n1049, CI => mult_21_C247_n1169, CO => 
                           mult_21_C247_n308, S => mult_21_C247_n309);
   mult_21_C247_U223 : ADFULD1 port map( A => mult_21_C247_n1141, B => 
                           mult_21_C247_n1001, CI => mult_21_C247_n989, CO => 
                           mult_21_C247_n306, S => mult_21_C247_n307);
   mult_21_C247_U222 : ADFULD1 port map( A => mult_21_C247_n1015, B => 
                           mult_21_C247_n1115, CI => mult_21_C247_n1069, CO => 
                           mult_21_C247_n304, S => mult_21_C247_n305);
   mult_21_C247_U221 : ADFULD1 port map( A => mult_21_C247_n313, B => 
                           mult_21_C247_n1091, CI => mult_21_C247_n336, CO => 
                           mult_21_C247_n302, S => mult_21_C247_n303);
   mult_21_C247_U220 : ADFULD1 port map( A => mult_21_C247_n332, B => 
                           mult_21_C247_n330, CI => mult_21_C247_n334, CO => 
                           mult_21_C247_n300, S => mult_21_C247_n301);
   mult_21_C247_U219 : ADFULD1 port map( A => mult_21_C247_n305, B => 
                           mult_21_C247_n328, CI => mult_21_C247_n311, CO => 
                           mult_21_C247_n298, S => mult_21_C247_n299);
   mult_21_C247_U218 : ADFULD1 port map( A => mult_21_C247_n307, B => 
                           mult_21_C247_n309, CI => mult_21_C247_n326, CO => 
                           mult_21_C247_n296, S => mult_21_C247_n297);
   mult_21_C247_U217 : ADFULD1 port map( A => mult_21_C247_n324, B => 
                           mult_21_C247_n303, CI => mult_21_C247_n301, CO => 
                           mult_21_C247_n294, S => mult_21_C247_n295);
   mult_21_C247_U216 : ADFULD1 port map( A => mult_21_C247_n299, B => 
                           mult_21_C247_n322, CI => mult_21_C247_n320, CO => 
                           mult_21_C247_n292, S => mult_21_C247_n293);
   mult_21_C247_U215 : ADFULD1 port map( A => mult_21_C247_n318, B => 
                           mult_21_C247_n297, CI => mult_21_C247_n295, CO => 
                           mult_21_C247_n290, S => mult_21_C247_n291);
   mult_21_C247_U214 : ADFULD1 port map( A => mult_21_C247_n316, B => 
                           mult_21_C247_n293, CI => mult_21_C247_n291, CO => 
                           mult_21_C247_n288, S => mult_21_C247_n289);
   mult_21_C247_U213 : ADHALFDL port map( A => mult_21_C247_n1198, B => 
                           mult_21_C247_n940, CO => mult_21_C247_n286, S => 
                           mult_21_C247_n287);
   mult_21_C247_U212 : ADFULD1 port map( A => mult_21_C247_n1030, B => 
                           mult_21_C247_n960, CI => mult_21_C247_n1168, CO => 
                           mult_21_C247_n284, S => mult_21_C247_n285);
   mult_21_C247_U211 : ADFULD1 port map( A => mult_21_C247_n1140, B => 
                           mult_21_C247_n1000, CI => mult_21_C247_n287, CO => 
                           mult_21_C247_n282, S => mult_21_C247_n283);
   mult_21_C247_U210 : ADFULD1 port map( A => mult_21_C247_n964, B => 
                           mult_21_C247_n1114, CI => mult_21_C247_n970, CO => 
                           mult_21_C247_n280, S => mult_21_C247_n281);
   mult_21_C247_U209 : ADFULD1 port map( A => mult_21_C247_n978, B => 
                           mult_21_C247_n1090, CI => mult_21_C247_n988, CO => 
                           mult_21_C247_n278, S => mult_21_C247_n279);
   mult_21_C247_U208 : ADFULD1 port map( A => mult_21_C247_n1014, B => 
                           mult_21_C247_n1068, CI => mult_21_C247_n1048, CO => 
                           mult_21_C247_n276, S => mult_21_C247_n277);
   mult_21_C247_U207 : ADFULD1 port map( A => mult_21_C247_n304, B => 
                           mult_21_C247_n312, CI => mult_21_C247_n306, CO => 
                           mult_21_C247_n274, S => mult_21_C247_n275);
   mult_21_C247_U206 : ADFULD1 port map( A => mult_21_C247_n310, B => 
                           mult_21_C247_n308, CI => mult_21_C247_n285, CO => 
                           mult_21_C247_n272, S => mult_21_C247_n273);
   mult_21_C247_U205 : ADFULD1 port map( A => mult_21_C247_n283, B => 
                           mult_21_C247_n277, CI => mult_21_C247_n279, CO => 
                           mult_21_C247_n270, S => mult_21_C247_n271);
   mult_21_C247_U204 : ADFULD1 port map( A => mult_21_C247_n302, B => 
                           mult_21_C247_n281, CI => mult_21_C247_n300, CO => 
                           mult_21_C247_n268, S => mult_21_C247_n269);
   mult_21_C247_U203 : ADFULD1 port map( A => mult_21_C247_n275, B => 
                           mult_21_C247_n298, CI => mult_21_C247_n273, CO => 
                           mult_21_C247_n266, S => mult_21_C247_n267);
   mult_21_C247_U202 : ADFULD1 port map( A => mult_21_C247_n296, B => 
                           mult_21_C247_n271, CI => mult_21_C247_n269, CO => 
                           mult_21_C247_n264, S => mult_21_C247_n265);
   mult_21_C247_U201 : ADFULD1 port map( A => mult_21_C247_n267, B => 
                           mult_21_C247_n294, CI => mult_21_C247_n292, CO => 
                           mult_21_C247_n262, S => mult_21_C247_n263);
   mult_21_C247_U200 : ADFULD1 port map( A => mult_21_C247_n290, B => 
                           mult_21_C247_n265, CI => mult_21_C247_n263, CO => 
                           mult_21_C247_n260, S => mult_21_C247_n261);
   mult_21_C247_U199 : ADHALFDL port map( A => mult_21_C247_n286, B => 
                           mult_21_C247_n1197, CO => mult_21_C247_n258, S => 
                           mult_21_C247_n259);
   mult_21_C247_U198 : ADFULD1 port map( A => mult_21_C247_n1167, B => 
                           mult_21_C247_n1029, CI => mult_21_C247_n1139, CO => 
                           mult_21_C247_n256, S => mult_21_C247_n257);
   mult_21_C247_U197 : ADFULD1 port map( A => mult_21_C247_n1113, B => 
                           mult_21_C247_n987, CI => mult_21_C247_n1089, CO => 
                           mult_21_C247_n254, S => mult_21_C247_n255);
   mult_21_C247_U196 : ADFULD1 port map( A => mult_21_C247_n959, B => 
                           mult_21_C247_n969, CI => mult_21_C247_n963, CO => 
                           mult_21_C247_n252, S => mult_21_C247_n253);
   mult_21_C247_U195 : ADFULD1 port map( A => mult_21_C247_n977, B => 
                           mult_21_C247_n1067, CI => mult_21_C247_n999, CO => 
                           mult_21_C247_n250, S => mult_21_C247_n251);
   mult_21_C247_U194 : ADFULD1 port map( A => mult_21_C247_n1047, B => 
                           mult_21_C247_n1013, CI => mult_21_C247_n259, CO => 
                           mult_21_C247_n248, S => mult_21_C247_n249);
   mult_21_C247_U193 : ADFULD1 port map( A => mult_21_C247_n278, B => 
                           mult_21_C247_n284, CI => mult_21_C247_n282, CO => 
                           mult_21_C247_n246, S => mult_21_C247_n247);
   mult_21_C247_U192 : ADFULD1 port map( A => mult_21_C247_n280, B => 
                           mult_21_C247_n276, CI => mult_21_C247_n251, CO => 
                           mult_21_C247_n244, S => mult_21_C247_n245);
   mult_21_C247_U191 : ADFULD1 port map( A => mult_21_C247_n253, B => 
                           mult_21_C247_n255, CI => mult_21_C247_n257, CO => 
                           mult_21_C247_n242, S => mult_21_C247_n243);
   mult_21_C247_U190 : ADFULD1 port map( A => mult_21_C247_n274, B => 
                           mult_21_C247_n249, CI => mult_21_C247_n272, CO => 
                           mult_21_C247_n240, S => mult_21_C247_n241);
   mult_21_C247_U189 : ADFULD1 port map( A => mult_21_C247_n270, B => 
                           mult_21_C247_n247, CI => mult_21_C247_n245, CO => 
                           mult_21_C247_n238, S => mult_21_C247_n239);
   mult_21_C247_U188 : ADFULD1 port map( A => mult_21_C247_n268, B => 
                           mult_21_C247_n243, CI => mult_21_C247_n241, CO => 
                           mult_21_C247_n236, S => mult_21_C247_n237);
   mult_21_C247_U187 : ADFULD1 port map( A => mult_21_C247_n239, B => 
                           mult_21_C247_n266, CI => mult_21_C247_n264, CO => 
                           mult_21_C247_n234, S => mult_21_C247_n235);
   mult_21_C247_U186 : ADFULD1 port map( A => mult_21_C247_n262, B => 
                           mult_21_C247_n237, CI => mult_21_C247_n235, CO => 
                           mult_21_C247_n232, S => mult_21_C247_n233);
   mult_21_C247_U185 : ADHALFDL port map( A => mult_21_C247_n1196, B => 
                           mult_21_C247_n939, CO => mult_21_C247_n230, S => 
                           mult_21_C247_n231);
   mult_21_C247_U184 : ADFULD1 port map( A => mult_21_C247_n1028, B => 
                           mult_21_C247_n956, CI => mult_21_C247_n958, CO => 
                           mult_21_C247_n228, S => mult_21_C247_n229);
   mult_21_C247_U183 : ADFULD1 port map( A => mult_21_C247_n1166, B => 
                           mult_21_C247_n1012, CI => mult_21_C247_n231, CO => 
                           mult_21_C247_n226, S => mult_21_C247_n227);
   mult_21_C247_U182 : ADFULD1 port map( A => mult_21_C247_n962, B => 
                           mult_21_C247_n1138, CI => mult_21_C247_n968, CO => 
                           mult_21_C247_n224, S => mult_21_C247_n225);
   mult_21_C247_U181 : ADFULD1 port map( A => mult_21_C247_n986, B => 
                           mult_21_C247_n976, CI => mult_21_C247_n998, CO => 
                           mult_21_C247_n222, S => mult_21_C247_n223);
   mult_21_C247_U180 : ADFULD1 port map( A => mult_21_C247_n1046, B => 
                           mult_21_C247_n1112, CI => mult_21_C247_n1066, CO => 
                           mult_21_C247_n220, S => mult_21_C247_n221);
   mult_21_C247_U179 : ADFULD1 port map( A => mult_21_C247_n258, B => 
                           mult_21_C247_n1088, CI => mult_21_C247_n250, CO => 
                           mult_21_C247_n218, S => mult_21_C247_n219);
   mult_21_C247_U178 : ADFULD1 port map( A => mult_21_C247_n256, B => 
                           mult_21_C247_n252, CI => mult_21_C247_n254, CO => 
                           mult_21_C247_n216, S => mult_21_C247_n217);
   mult_21_C247_U177 : ADFULD1 port map( A => mult_21_C247_n221, B => 
                           mult_21_C247_n229, CI => mult_21_C247_n227, CO => 
                           mult_21_C247_n214, S => mult_21_C247_n215);
   mult_21_C247_U176 : ADFULD1 port map( A => mult_21_C247_n225, B => 
                           mult_21_C247_n223, CI => mult_21_C247_n248, CO => 
                           mult_21_C247_n212, S => mult_21_C247_n213);
   mult_21_C247_U175 : ADFULD1 port map( A => mult_21_C247_n244, B => 
                           mult_21_C247_n246, CI => mult_21_C247_n219, CO => 
                           mult_21_C247_n210, S => mult_21_C247_n211);
   mult_21_C247_U174 : ADFULD1 port map( A => mult_21_C247_n217, B => 
                           mult_21_C247_n242, CI => mult_21_C247_n215, CO => 
                           mult_21_C247_n208, S => mult_21_C247_n209);
   mult_21_C247_U173 : ADFULD1 port map( A => mult_21_C247_n240, B => 
                           mult_21_C247_n213, CI => mult_21_C247_n238, CO => 
                           mult_21_C247_n206, S => mult_21_C247_n207);
   mult_21_C247_U172 : ADFULD1 port map( A => mult_21_C247_n209, B => 
                           mult_21_C247_n211, CI => mult_21_C247_n236, CO => 
                           mult_21_C247_n204, S => mult_21_C247_n205);
   mult_21_C247_U171 : ADFULD1 port map( A => mult_21_C247_n234, B => 
                           mult_21_C247_n207, CI => mult_21_C247_n205, CO => 
                           mult_21_C247_n202, S => mult_21_C247_n203);
   mult_21_C247_U155 : ADHALFDL port map( A => mult_21_C247_n1226, B => N3010, 
                           CO => mult_21_C247_n186, S => N3329);
   mult_21_C247_U154 : ADHALFDL port map( A => mult_21_C247_n186, B => 
                           mult_21_C247_n1225, CO => mult_21_C247_n185, S => 
                           N3330);
   mult_21_C247_U153 : ADFULD1 port map( A => mult_21_C247_n651, B => 
                           mult_21_C247_n1194, CI => mult_21_C247_n185, CO => 
                           mult_21_C247_n184, S => N3331);
   mult_21_C247_U152 : ADFULD1 port map( A => mult_21_C247_n649, B => 
                           mult_21_C247_n1193, CI => mult_21_C247_n184, CO => 
                           mult_21_C247_n183, S => N3332);
   mult_21_C247_U151 : ADFULD1 port map( A => mult_21_C247_n645, B => 
                           mult_21_C247_n648, CI => mult_21_C247_n183, CO => 
                           mult_21_C247_n182, S => N3333);
   mult_21_C247_U150 : ADFULD1 port map( A => mult_21_C247_n641, B => 
                           mult_21_C247_n644, CI => mult_21_C247_n182, CO => 
                           mult_21_C247_n181, S => N3334);
   mult_21_C247_U149 : ADFULD1 port map( A => mult_21_C247_n635, B => 
                           mult_21_C247_n640, CI => mult_21_C247_n181, CO => 
                           mult_21_C247_n180, S => N3335);
   mult_21_C247_U148 : ADFULD1 port map( A => mult_21_C247_n629, B => 
                           mult_21_C247_n634, CI => mult_21_C247_n180, CO => 
                           mult_21_C247_n179, S => N3336);
   mult_21_C247_U147 : ADFULD1 port map( A => mult_21_C247_n621, B => 
                           mult_21_C247_n628, CI => mult_21_C247_n179, CO => 
                           mult_21_C247_n178, S => N3337);
   mult_21_C247_U146 : ADFULD1 port map( A => mult_21_C247_n613, B => 
                           mult_21_C247_n620, CI => mult_21_C247_n178, CO => 
                           mult_21_C247_n177, S => N3338);
   mult_21_C247_U145 : ADFULD1 port map( A => mult_21_C247_n603, B => 
                           mult_21_C247_n612, CI => mult_21_C247_n177, CO => 
                           mult_21_C247_n176, S => N3339);
   mult_21_C247_U144 : ADFULD1 port map( A => mult_21_C247_n593, B => 
                           mult_21_C247_n602, CI => mult_21_C247_n176, CO => 
                           mult_21_C247_n175, S => N3340);
   mult_21_C247_U143 : ADFULD1 port map( A => mult_21_C247_n581, B => 
                           mult_21_C247_n592, CI => mult_21_C247_n175, CO => 
                           mult_21_C247_n174, S => N3341);
   mult_21_C247_U142 : ADFULD1 port map( A => mult_21_C247_n569, B => 
                           mult_21_C247_n580, CI => mult_21_C247_n174, CO => 
                           mult_21_C247_n173, S => N3342);
   mult_21_C247_U141 : ADFULD1 port map( A => mult_21_C247_n555, B => 
                           mult_21_C247_n568, CI => mult_21_C247_n173, CO => 
                           mult_21_C247_n172, S => N3343);
   mult_21_C247_U140 : ADFULD1 port map( A => mult_21_C247_n541, B => 
                           mult_21_C247_n554, CI => mult_21_C247_n172, CO => 
                           mult_21_C247_n171, S => N3344);
   mult_21_C247_U139 : ADFULD1 port map( A => mult_21_C247_n525, B => 
                           mult_21_C247_n540, CI => mult_21_C247_n171, CO => 
                           mult_21_C247_n170, S => N3345);
   mult_21_C247_U138 : ADFULD1 port map( A => mult_21_C247_n509, B => 
                           mult_21_C247_n524, CI => mult_21_C247_n170, CO => 
                           mult_21_C247_n169, S => N3346);
   mult_21_C247_U137 : ADFULD1 port map( A => mult_21_C247_n491, B => 
                           mult_21_C247_n508, CI => mult_21_C247_n169, CO => 
                           mult_21_C247_n168, S => N3347);
   mult_21_C247_U136 : ADFULD1 port map( A => mult_21_C247_n473, B => 
                           mult_21_C247_n490, CI => mult_21_C247_n168, CO => 
                           mult_21_C247_n167, S => N3348);
   mult_21_C247_U135 : ADFULD1 port map( A => mult_21_C247_n453, B => 
                           mult_21_C247_n472, CI => mult_21_C247_n167, CO => 
                           mult_21_C247_n166, S => N3349);
   mult_21_C247_U134 : ADFULD1 port map( A => mult_21_C247_n433, B => 
                           mult_21_C247_n452, CI => mult_21_C247_n166, CO => 
                           mult_21_C247_n165, S => N3350);
   mult_21_C247_U133 : ADFULD1 port map( A => mult_21_C247_n411, B => 
                           mult_21_C247_n432, CI => mult_21_C247_n165, CO => 
                           mult_21_C247_n164, S => N3351);
   mult_21_C247_U132 : ADFULD1 port map( A => mult_21_C247_n389, B => 
                           mult_21_C247_n410, CI => mult_21_C247_n164, CO => 
                           mult_21_C247_n163, S => N3352);
   mult_21_C247_U131 : ADFULD1 port map( A => mult_21_C247_n365, B => 
                           mult_21_C247_n388, CI => mult_21_C247_n163, CO => 
                           mult_21_C247_n162, S => N3353);
   mult_21_C247_U130 : ADFULD1 port map( A => mult_21_C247_n341, B => 
                           mult_21_C247_n364, CI => mult_21_C247_n162, CO => 
                           mult_21_C247_n161, S => N3354);
   mult_21_C247_U129 : ADFULD1 port map( A => mult_21_C247_n315, B => 
                           mult_21_C247_n340, CI => mult_21_C247_n161, CO => 
                           mult_21_C247_n160, S => N3355);
   mult_21_C247_U128 : ADFULD1 port map( A => mult_21_C247_n289, B => 
                           mult_21_C247_n314, CI => mult_21_C247_n160, CO => 
                           mult_21_C247_n159, S => N3356);
   mult_21_C247_U127 : ADFULD1 port map( A => mult_21_C247_n261, B => 
                           mult_21_C247_n288, CI => mult_21_C247_n159, CO => 
                           mult_21_C247_n158, S => N3357);
   mult_21_C247_U126 : ADFULD1 port map( A => mult_21_C247_n233, B => 
                           mult_21_C247_n260, CI => mult_21_C247_n158, CO => 
                           mult_21_C247_n157, S => N3358);
   mult_21_C247_U125 : ADFULD1 port map( A => mult_21_C247_n203, B => 
                           mult_21_C247_n232, CI => mult_21_C247_n157, CO => 
                           mult_21_C247_n156, S => N3359);
   mult_21_C249_U1399 : AOI21D1 port map( A1 => N3068, A2 => N3069, B => 
                           mult_21_C249_n1424, Z => mult_21_C249_n940);
   mult_21_C249_U1398 : OAI21D1 port map( A1 => N3071, A2 => N3070, B => 
                           mult_21_C249_n1425, Z => mult_21_C249_n104);
   mult_21_C249_U1397 : AOI21D1 port map( A1 => N3070, A2 => N3071, B => 
                           mult_21_C249_n1425, Z => mult_21_C249_n939);
   mult_21_C249_U1396 : AOI21D1 port map( A1 => N3042, A2 => N3043, B => 
                           mult_21_C249_n1398, Z => mult_21_C249_n953);
   mult_21_C249_U1395 : AOI21D1 port map( A1 => N3044, A2 => N3045, B => 
                           mult_21_C249_n1400, Z => mult_21_C249_n952);
   mult_21_C249_U1394 : AOI21D1 port map( A1 => N3046, A2 => N3047, B => 
                           mult_21_C249_n1402, Z => mult_21_C249_n951);
   mult_21_C249_U1393 : AOI21D1 port map( A1 => N3048, A2 => N3049, B => 
                           mult_21_C249_n1404, Z => mult_21_C249_n950);
   mult_21_C249_U1392 : AOI21D1 port map( A1 => N3050, A2 => N3051, B => 
                           mult_21_C249_n1406, Z => mult_21_C249_n949);
   mult_21_C249_U1391 : AOI21D1 port map( A1 => N3052, A2 => N3053, B => 
                           mult_21_C249_n1408, Z => mult_21_C249_n948);
   mult_21_C249_U1390 : AOI21D1 port map( A1 => N3054, A2 => N3055, B => 
                           mult_21_C249_n1410, Z => mult_21_C249_n947);
   mult_21_C249_U1389 : EXOR2D1 port map( A1 => N3071, A2 => N3070, Z => 
                           mult_21_C249_n1454);
   mult_21_C249_U1388 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C249_n1454, Z => mult_21_C249_n652);
   mult_21_C249_U1387 : NAN2D1 port map( A1 => N3201, A2 => mult_21_C249_n1454,
                           Z => mult_21_C249_n653);
   mult_21_C249_U1386 : EXOR2D1 port map( A1 => N3069, A2 => N3068, Z => 
                           mult_21_C249_n1453);
   mult_21_C249_U1385 : MUXB2DL port map( A0 => N3203, A1 => N3204, SL => 
                           mult_21_C249_n1453, Z => mult_21_C249_n654);
   mult_21_C249_U1384 : MUXB2DL port map( A0 => mult_21_C249_n1391, A1 => 
                           mult_21_C249_n1389, SL => mult_21_C249_n1453, Z => 
                           mult_21_C249_n655);
   mult_21_C249_U1383 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C249_n1453, Z => mult_21_C249_n656);
   mult_21_C249_U1382 : NAN2D1 port map( A1 => N3201, A2 => mult_21_C249_n1453,
                           Z => mult_21_C249_n657);
   mult_21_C249_U1381 : EXOR2D1 port map( A1 => N3067, A2 => N3066, Z => 
                           mult_21_C249_n1452);
   mult_21_C249_U1380 : MUXB2DL port map( A0 => N3205, A1 => mult_21_C249_n1385
                           , SL => mult_21_C249_n1452, Z => mult_21_C249_n658);
   mult_21_C249_U1379 : MUXB2DL port map( A0 => mult_21_C249_n1387, A1 => N3205
                           , SL => mult_21_C249_n1452, Z => mult_21_C249_n659);
   mult_21_C249_U1378 : MUXB2DL port map( A0 => N3203, A1 => N3204, SL => 
                           mult_21_C249_n1452, Z => mult_21_C249_n660);
   mult_21_C249_U1377 : MUXB2DL port map( A0 => mult_21_C249_n1391, A1 => N3203
                           , SL => mult_21_C249_n1452, Z => mult_21_C249_n661);
   mult_21_C249_U1376 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C249_n1452, Z => mult_21_C249_n662);
   mult_21_C249_U1375 : NAN2D1 port map( A1 => N3201, A2 => mult_21_C249_n1452,
                           Z => mult_21_C249_n663);
   mult_21_C249_U1374 : EXOR2D1 port map( A1 => N3065, A2 => N3064, Z => 
                           mult_21_C249_n1451);
   mult_21_C249_U1373 : MUXB2DL port map( A0 => N3207, A1 => N3208, SL => 
                           mult_21_C249_n1451, Z => mult_21_C249_n664);
   mult_21_C249_U1372 : MUXB2DL port map( A0 => N3206, A1 => N3207, SL => 
                           mult_21_C249_n1451, Z => mult_21_C249_n665);
   mult_21_C249_U1371 : MUXB2DL port map( A0 => N3205, A1 => N3206, SL => 
                           mult_21_C249_n1451, Z => mult_21_C249_n666);
   mult_21_C249_U1370 : MUXB2DL port map( A0 => mult_21_C249_n1387, A1 => N3205
                           , SL => mult_21_C249_n1451, Z => mult_21_C249_n667);
   mult_21_C249_U1369 : MUXB2DL port map( A0 => N3203, A1 => N3204, SL => 
                           mult_21_C249_n1451, Z => mult_21_C249_n668);
   mult_21_C249_U1368 : MUXB2DL port map( A0 => mult_21_C249_n1391, A1 => N3203
                           , SL => mult_21_C249_n1451, Z => mult_21_C249_n669);
   mult_21_C249_U1367 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C249_n1451, Z => mult_21_C249_n670);
   mult_21_C249_U1366 : NAN2D1 port map( A1 => N3201, A2 => mult_21_C249_n1451,
                           Z => mult_21_C249_n671);
   mult_21_C249_U1365 : MUXB2DL port map( A0 => N3209, A1 => N3210, SL => 
                           mult_21_C249_n1450, Z => mult_21_C249_n672);
   mult_21_C249_U1364 : MUXB2DL port map( A0 => N3208, A1 => N3209, SL => 
                           mult_21_C249_n1450, Z => mult_21_C249_n673);
   mult_21_C249_U1363 : MUXB2DL port map( A0 => N3207, A1 => N3208, SL => 
                           mult_21_C249_n1450, Z => mult_21_C249_n674);
   mult_21_C249_U1362 : MUXB2DL port map( A0 => N3206, A1 => N3207, SL => 
                           mult_21_C249_n1450, Z => mult_21_C249_n675);
   mult_21_C249_U1361 : MUXB2DL port map( A0 => N3205, A1 => mult_21_C249_n1385
                           , SL => mult_21_C249_n1450, Z => mult_21_C249_n676);
   mult_21_C249_U1360 : MUXB2DL port map( A0 => mult_21_C249_n1387, A1 => N3205
                           , SL => mult_21_C249_n1450, Z => mult_21_C249_n677);
   mult_21_C249_U1359 : MUXB2DL port map( A0 => N3203, A1 => N3204, SL => 
                           mult_21_C249_n1450, Z => mult_21_C249_n678);
   mult_21_C249_U1358 : MUXB2DL port map( A0 => mult_21_C249_n1391, A1 => N3203
                           , SL => mult_21_C249_n1450, Z => mult_21_C249_n679);
   mult_21_C249_U1357 : AOI21D1 port map( A1 => N3056, A2 => N3057, B => 
                           mult_21_C249_n1412, Z => mult_21_C249_n946);
   mult_21_C249_U1356 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C249_n1450, Z => mult_21_C249_n680);
   mult_21_C249_U1355 : NAN2D1 port map( A1 => mult_21_C249_n1393, A2 => 
                           mult_21_C249_n1450, Z => mult_21_C249_n681);
   mult_21_C249_U1354 : MUXB2DL port map( A0 => N3211, A1 => N3212, SL => 
                           mult_21_C249_n1449, Z => mult_21_C249_n682);
   mult_21_C249_U1353 : MUXB2DL port map( A0 => N3210, A1 => N3211, SL => 
                           mult_21_C249_n1449, Z => mult_21_C249_n683);
   mult_21_C249_U1352 : MUXB2DL port map( A0 => N3209, A1 => N3210, SL => 
                           mult_21_C249_n1449, Z => mult_21_C249_n684);
   mult_21_C249_U1351 : MUXB2DL port map( A0 => N3208, A1 => N3209, SL => 
                           mult_21_C249_n1449, Z => mult_21_C249_n685);
   mult_21_C249_U1350 : MUXB2DL port map( A0 => N3207, A1 => N3208, SL => 
                           mult_21_C249_n1449, Z => mult_21_C249_n686);
   mult_21_C249_U1349 : MUXB2DL port map( A0 => N3206, A1 => N3207, SL => 
                           mult_21_C249_n1449, Z => mult_21_C249_n687);
   mult_21_C249_U1348 : MUXB2DL port map( A0 => N3205, A1 => mult_21_C249_n1385
                           , SL => mult_21_C249_n1449, Z => mult_21_C249_n688);
   mult_21_C249_U1347 : MUXB2DL port map( A0 => mult_21_C249_n1387, A1 => N3205
                           , SL => mult_21_C249_n1449, Z => mult_21_C249_n689);
   mult_21_C249_U1346 : MUXB2DL port map( A0 => N3203, A1 => N3204, SL => 
                           mult_21_C249_n1449, Z => mult_21_C249_n690);
   mult_21_C249_U1345 : MUXB2DL port map( A0 => mult_21_C249_n1391, A1 => N3203
                           , SL => mult_21_C249_n1449, Z => mult_21_C249_n691);
   mult_21_C249_U1344 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C249_n1449, Z => mult_21_C249_n692);
   mult_21_C249_U1343 : NAN2D1 port map( A1 => mult_21_C249_n1393, A2 => 
                           mult_21_C249_n1449, Z => mult_21_C249_n693);
   mult_21_C249_U1342 : MUXB2DL port map( A0 => N3213, A1 => N3214, SL => 
                           mult_21_C249_n1448, Z => mult_21_C249_n694);
   mult_21_C249_U1341 : MUXB2DL port map( A0 => N3212, A1 => N3213, SL => 
                           mult_21_C249_n1448, Z => mult_21_C249_n695);
   mult_21_C249_U1340 : MUXB2DL port map( A0 => N3211, A1 => N3212, SL => 
                           mult_21_C249_n1448, Z => mult_21_C249_n696);
   mult_21_C249_U1339 : MUXB2DL port map( A0 => N3210, A1 => N3211, SL => 
                           mult_21_C249_n1448, Z => mult_21_C249_n697);
   mult_21_C249_U1338 : MUXB2DL port map( A0 => N3209, A1 => N3210, SL => 
                           mult_21_C249_n1448, Z => mult_21_C249_n698);
   mult_21_C249_U1337 : MUXB2DL port map( A0 => N3208, A1 => N3209, SL => 
                           mult_21_C249_n1448, Z => mult_21_C249_n699);
   mult_21_C249_U1336 : MUXB2DL port map( A0 => N3207, A1 => N3208, SL => 
                           mult_21_C249_n1448, Z => mult_21_C249_n700);
   mult_21_C249_U1335 : MUXB2DL port map( A0 => N3206, A1 => N3207, SL => 
                           mult_21_C249_n1448, Z => mult_21_C249_n701);
   mult_21_C249_U1334 : MUXB2DL port map( A0 => N3205, A1 => mult_21_C249_n1385
                           , SL => mult_21_C249_n1448, Z => mult_21_C249_n702);
   mult_21_C249_U1333 : MUXB2DL port map( A0 => mult_21_C249_n1387, A1 => N3205
                           , SL => mult_21_C249_n1448, Z => mult_21_C249_n703);
   mult_21_C249_U1332 : MUXB2DL port map( A0 => N3203, A1 => N3204, SL => 
                           mult_21_C249_n1448, Z => mult_21_C249_n704);
   mult_21_C249_U1331 : MUXB2DL port map( A0 => mult_21_C249_n1391, A1 => 
                           mult_21_C249_n1389, SL => mult_21_C249_n1448, Z => 
                           mult_21_C249_n705);
   mult_21_C249_U1330 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C249_n1448, Z => mult_21_C249_n706);
   mult_21_C249_U1329 : NAN2D1 port map( A1 => mult_21_C249_n1393, A2 => 
                           mult_21_C249_n1448, Z => mult_21_C249_n707);
   mult_21_C249_U1328 : MUXB2DL port map( A0 => N3215, A1 => N3216, SL => 
                           mult_21_C249_n1447, Z => mult_21_C249_n708);
   mult_21_C249_U1327 : MUXB2DL port map( A0 => N3214, A1 => N3215, SL => 
                           mult_21_C249_n1447, Z => mult_21_C249_n709);
   mult_21_C249_U1326 : MUXB2DL port map( A0 => N3213, A1 => N3214, SL => 
                           mult_21_C249_n1447, Z => mult_21_C249_n710);
   mult_21_C249_U1325 : MUXB2DL port map( A0 => N3212, A1 => N3213, SL => 
                           mult_21_C249_n1447, Z => mult_21_C249_n711);
   mult_21_C249_U1324 : MUXB2DL port map( A0 => N3211, A1 => N3212, SL => 
                           mult_21_C249_n1447, Z => mult_21_C249_n712);
   mult_21_C249_U1323 : MUXB2DL port map( A0 => N3210, A1 => N3211, SL => 
                           mult_21_C249_n1447, Z => mult_21_C249_n713);
   mult_21_C249_U1322 : MUXB2DL port map( A0 => N3209, A1 => N3210, SL => 
                           mult_21_C249_n1447, Z => mult_21_C249_n714);
   mult_21_C249_U1321 : MUXB2DL port map( A0 => N3208, A1 => N3209, SL => 
                           mult_21_C249_n1447, Z => mult_21_C249_n715);
   mult_21_C249_U1320 : MUXB2DL port map( A0 => N3207, A1 => N3208, SL => 
                           mult_21_C249_n1447, Z => mult_21_C249_n716);
   mult_21_C249_U1319 : MUXB2DL port map( A0 => N3206, A1 => N3207, SL => 
                           mult_21_C249_n1447, Z => mult_21_C249_n717);
   mult_21_C249_U1318 : MUXB2DL port map( A0 => N3205, A1 => mult_21_C249_n1385
                           , SL => mult_21_C249_n1447, Z => mult_21_C249_n718);
   mult_21_C249_U1317 : MUXB2DL port map( A0 => mult_21_C249_n1387, A1 => N3205
                           , SL => mult_21_C249_n1447, Z => mult_21_C249_n719);
   mult_21_C249_U1316 : MUXB2DL port map( A0 => N3203, A1 => N3204, SL => 
                           mult_21_C249_n1447, Z => mult_21_C249_n720);
   mult_21_C249_U1315 : MUXB2DL port map( A0 => mult_21_C249_n1391, A1 => 
                           mult_21_C249_n1389, SL => mult_21_C249_n1447, Z => 
                           mult_21_C249_n721);
   mult_21_C249_U1314 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C249_n1447, Z => mult_21_C249_n722);
   mult_21_C249_U1313 : NAN2D1 port map( A1 => mult_21_C249_n1393, A2 => 
                           mult_21_C249_n1447, Z => mult_21_C249_n723);
   mult_21_C249_U1312 : MUXB2DL port map( A0 => N3217, A1 => N3218, SL => 
                           mult_21_C249_n1446, Z => mult_21_C249_n724);
   mult_21_C249_U1311 : MUXB2DL port map( A0 => N3216, A1 => N3217, SL => 
                           mult_21_C249_n1446, Z => mult_21_C249_n725);
   mult_21_C249_U1310 : MUXB2DL port map( A0 => N3215, A1 => N3216, SL => 
                           mult_21_C249_n1446, Z => mult_21_C249_n726);
   mult_21_C249_U1309 : MUXB2DL port map( A0 => N3214, A1 => N3215, SL => 
                           mult_21_C249_n1446, Z => mult_21_C249_n727);
   mult_21_C249_U1308 : MUXB2DL port map( A0 => N3213, A1 => N3214, SL => 
                           mult_21_C249_n1446, Z => mult_21_C249_n728);
   mult_21_C249_U1307 : MUXB2DL port map( A0 => N3212, A1 => N3213, SL => 
                           mult_21_C249_n1446, Z => mult_21_C249_n729);
   mult_21_C249_U1306 : MUXB2DL port map( A0 => N3211, A1 => N3212, SL => 
                           mult_21_C249_n1446, Z => mult_21_C249_n730);
   mult_21_C249_U1305 : MUXB2DL port map( A0 => N3210, A1 => N3211, SL => 
                           mult_21_C249_n1446, Z => mult_21_C249_n731);
   mult_21_C249_U1304 : MUXB2DL port map( A0 => N3209, A1 => N3210, SL => 
                           mult_21_C249_n1446, Z => mult_21_C249_n732);
   mult_21_C249_U1303 : MUXB2DL port map( A0 => N3208, A1 => N3209, SL => 
                           mult_21_C249_n1446, Z => mult_21_C249_n733);
   mult_21_C249_U1302 : MUXB2DL port map( A0 => N3207, A1 => N3208, SL => 
                           mult_21_C249_n1446, Z => mult_21_C249_n734);
   mult_21_C249_U1301 : MUXB2DL port map( A0 => N3206, A1 => N3207, SL => 
                           mult_21_C249_n1446, Z => mult_21_C249_n735);
   mult_21_C249_U1300 : MUXB2DL port map( A0 => N3205, A1 => mult_21_C249_n1385
                           , SL => mult_21_C249_n1446, Z => mult_21_C249_n736);
   mult_21_C249_U1299 : MUXB2DL port map( A0 => mult_21_C249_n1387, A1 => N3205
                           , SL => mult_21_C249_n1446, Z => mult_21_C249_n737);
   mult_21_C249_U1298 : MUXB2DL port map( A0 => N3203, A1 => N3204, SL => 
                           mult_21_C249_n1446, Z => mult_21_C249_n738);
   mult_21_C249_U1297 : MUXB2DL port map( A0 => mult_21_C249_n1391, A1 => 
                           mult_21_C249_n1389, SL => mult_21_C249_n1446, Z => 
                           mult_21_C249_n739);
   mult_21_C249_U1296 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C249_n1446, Z => mult_21_C249_n740);
   mult_21_C249_U1295 : NAN2D1 port map( A1 => mult_21_C249_n1393, A2 => 
                           mult_21_C249_n1446, Z => mult_21_C249_n741);
   mult_21_C249_U1294 : MUXB2DL port map( A0 => N3219, A1 => N3220, SL => 
                           mult_21_C249_n1445, Z => mult_21_C249_n742);
   mult_21_C249_U1293 : MUXB2DL port map( A0 => N3218, A1 => N3219, SL => 
                           mult_21_C249_n1445, Z => mult_21_C249_n743);
   mult_21_C249_U1292 : MUXB2DL port map( A0 => N3217, A1 => N3218, SL => 
                           mult_21_C249_n1445, Z => mult_21_C249_n744);
   mult_21_C249_U1291 : MUXB2DL port map( A0 => N3216, A1 => N3217, SL => 
                           mult_21_C249_n1445, Z => mult_21_C249_n745);
   mult_21_C249_U1290 : MUXB2DL port map( A0 => N3215, A1 => N3216, SL => 
                           mult_21_C249_n1445, Z => mult_21_C249_n746);
   mult_21_C249_U1289 : MUXB2DL port map( A0 => N3214, A1 => N3215, SL => 
                           mult_21_C249_n1445, Z => mult_21_C249_n747);
   mult_21_C249_U1288 : MUXB2DL port map( A0 => N3213, A1 => N3214, SL => 
                           mult_21_C249_n1445, Z => mult_21_C249_n748);
   mult_21_C249_U1287 : MUXB2DL port map( A0 => N3212, A1 => N3213, SL => 
                           mult_21_C249_n1445, Z => mult_21_C249_n749);
   mult_21_C249_U1286 : AOI21D1 port map( A1 => N3058, A2 => N3059, B => 
                           mult_21_C249_n1414, Z => mult_21_C249_n945);
   mult_21_C249_U1285 : MUXB2DL port map( A0 => N3211, A1 => N3212, SL => 
                           mult_21_C249_n1445, Z => mult_21_C249_n750);
   mult_21_C249_U1284 : MUXB2DL port map( A0 => N3210, A1 => N3211, SL => 
                           mult_21_C249_n1445, Z => mult_21_C249_n751);
   mult_21_C249_U1283 : MUXB2DL port map( A0 => N3209, A1 => N3210, SL => 
                           mult_21_C249_n1445, Z => mult_21_C249_n752);
   mult_21_C249_U1282 : MUXB2DL port map( A0 => N3208, A1 => N3209, SL => 
                           mult_21_C249_n1445, Z => mult_21_C249_n753);
   mult_21_C249_U1281 : MUXB2DL port map( A0 => N3207, A1 => N3208, SL => 
                           mult_21_C249_n1445, Z => mult_21_C249_n754);
   mult_21_C249_U1280 : MUXB2DL port map( A0 => N3206, A1 => N3207, SL => 
                           mult_21_C249_n1445, Z => mult_21_C249_n755);
   mult_21_C249_U1279 : MUXB2DL port map( A0 => N3205, A1 => mult_21_C249_n1385
                           , SL => mult_21_C249_n1445, Z => mult_21_C249_n756);
   mult_21_C249_U1278 : MUXB2DL port map( A0 => mult_21_C249_n1387, A1 => N3205
                           , SL => mult_21_C249_n1445, Z => mult_21_C249_n757);
   mult_21_C249_U1277 : MUXB2DL port map( A0 => N3203, A1 => N3204, SL => 
                           mult_21_C249_n1445, Z => mult_21_C249_n758);
   mult_21_C249_U1276 : MUXB2DL port map( A0 => N3202, A1 => mult_21_C249_n1389
                           , SL => mult_21_C249_n1445, Z => mult_21_C249_n759);
   mult_21_C249_U1275 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C249_n1445, Z => mult_21_C249_n760);
   mult_21_C249_U1274 : NAN2D1 port map( A1 => mult_21_C249_n1393, A2 => 
                           mult_21_C249_n1445, Z => mult_21_C249_n761);
   mult_21_C249_U1273 : MUXB2DL port map( A0 => N3221, A1 => N3222, SL => 
                           mult_21_C249_n1444, Z => mult_21_C249_n762);
   mult_21_C249_U1272 : MUXB2DL port map( A0 => N3220, A1 => N3221, SL => 
                           mult_21_C249_n1444, Z => mult_21_C249_n763);
   mult_21_C249_U1271 : MUXB2DL port map( A0 => N3219, A1 => N3220, SL => 
                           mult_21_C249_n1444, Z => mult_21_C249_n764);
   mult_21_C249_U1270 : MUXB2DL port map( A0 => N3218, A1 => N3219, SL => 
                           mult_21_C249_n1444, Z => mult_21_C249_n765);
   mult_21_C249_U1269 : MUXB2DL port map( A0 => N3217, A1 => N3218, SL => 
                           mult_21_C249_n1444, Z => mult_21_C249_n766);
   mult_21_C249_U1268 : MUXB2DL port map( A0 => N3216, A1 => N3217, SL => 
                           mult_21_C249_n1444, Z => mult_21_C249_n767);
   mult_21_C249_U1267 : MUXB2DL port map( A0 => N3215, A1 => N3216, SL => 
                           mult_21_C249_n1444, Z => mult_21_C249_n768);
   mult_21_C249_U1266 : MUXB2DL port map( A0 => N3214, A1 => N3215, SL => 
                           mult_21_C249_n1444, Z => mult_21_C249_n769);
   mult_21_C249_U1265 : MUXB2DL port map( A0 => N3213, A1 => N3214, SL => 
                           mult_21_C249_n1444, Z => mult_21_C249_n770);
   mult_21_C249_U1264 : MUXB2DL port map( A0 => N3212, A1 => N3213, SL => 
                           mult_21_C249_n1444, Z => mult_21_C249_n771);
   mult_21_C249_U1263 : MUXB2DL port map( A0 => N3211, A1 => N3212, SL => 
                           mult_21_C249_n1444, Z => mult_21_C249_n772);
   mult_21_C249_U1262 : MUXB2DL port map( A0 => N3210, A1 => N3211, SL => 
                           mult_21_C249_n1444, Z => mult_21_C249_n773);
   mult_21_C249_U1261 : MUXB2DL port map( A0 => N3209, A1 => N3210, SL => 
                           mult_21_C249_n1444, Z => mult_21_C249_n774);
   mult_21_C249_U1260 : MUXB2DL port map( A0 => N3208, A1 => N3209, SL => 
                           mult_21_C249_n1444, Z => mult_21_C249_n775);
   mult_21_C249_U1259 : MUXB2DL port map( A0 => N3207, A1 => N3208, SL => 
                           mult_21_C249_n1444, Z => mult_21_C249_n776);
   mult_21_C249_U1258 : MUXB2DL port map( A0 => N3206, A1 => N3207, SL => 
                           mult_21_C249_n1444, Z => mult_21_C249_n777);
   mult_21_C249_U1257 : MUXB2DL port map( A0 => N3205, A1 => mult_21_C249_n1385
                           , SL => mult_21_C249_n1444, Z => mult_21_C249_n778);
   mult_21_C249_U1256 : MUXB2DL port map( A0 => N3204, A1 => N3205, SL => 
                           mult_21_C249_n1444, Z => mult_21_C249_n779);
   mult_21_C249_U1255 : MUXB2DL port map( A0 => mult_21_C249_n1389, A1 => N3204
                           , SL => mult_21_C249_n1444, Z => mult_21_C249_n780);
   mult_21_C249_U1254 : MUXB2DL port map( A0 => mult_21_C249_n1391, A1 => 
                           mult_21_C249_n1389, SL => mult_21_C249_n1444, Z => 
                           mult_21_C249_n781);
   mult_21_C249_U1253 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C249_n1444, Z => mult_21_C249_n782);
   mult_21_C249_U1252 : NAN2D1 port map( A1 => mult_21_C249_n1393, A2 => 
                           mult_21_C249_n1444, Z => mult_21_C249_n783);
   mult_21_C249_U1251 : MUXB2DL port map( A0 => N3223, A1 => N3224, SL => 
                           mult_21_C249_n1377, Z => mult_21_C249_n784);
   mult_21_C249_U1250 : MUXB2DL port map( A0 => N3222, A1 => N3223, SL => 
                           mult_21_C249_n1377, Z => mult_21_C249_n785);
   mult_21_C249_U1249 : MUXB2DL port map( A0 => N3221, A1 => N3222, SL => 
                           mult_21_C249_n1377, Z => mult_21_C249_n786);
   mult_21_C249_U1248 : MUXB2DL port map( A0 => N3220, A1 => N3221, SL => 
                           mult_21_C249_n1377, Z => mult_21_C249_n787);
   mult_21_C249_U1247 : MUXB2DL port map( A0 => N3219, A1 => N3220, SL => 
                           mult_21_C249_n1377, Z => mult_21_C249_n788);
   mult_21_C249_U1246 : MUXB2DL port map( A0 => N3218, A1 => N3219, SL => 
                           mult_21_C249_n1377, Z => mult_21_C249_n789);
   mult_21_C249_U1245 : MUXB2DL port map( A0 => N3217, A1 => N3218, SL => 
                           mult_21_C249_n1377, Z => mult_21_C249_n790);
   mult_21_C249_U1244 : MUXB2DL port map( A0 => N3216, A1 => N3217, SL => 
                           mult_21_C249_n1377, Z => mult_21_C249_n791);
   mult_21_C249_U1243 : MUXB2DL port map( A0 => N3215, A1 => N3216, SL => 
                           mult_21_C249_n1377, Z => mult_21_C249_n792);
   mult_21_C249_U1242 : MUXB2DL port map( A0 => N3214, A1 => N3215, SL => 
                           mult_21_C249_n1377, Z => mult_21_C249_n793);
   mult_21_C249_U1241 : MUXB2DL port map( A0 => N3213, A1 => N3214, SL => 
                           mult_21_C249_n1377, Z => mult_21_C249_n794);
   mult_21_C249_U1240 : MUXB2DL port map( A0 => N3212, A1 => N3213, SL => 
                           mult_21_C249_n1377, Z => mult_21_C249_n795);
   mult_21_C249_U1239 : MUXB2DL port map( A0 => N3211, A1 => N3212, SL => 
                           mult_21_C249_n1377, Z => mult_21_C249_n796);
   mult_21_C249_U1238 : MUXB2DL port map( A0 => N3210, A1 => N3211, SL => 
                           mult_21_C249_n1377, Z => mult_21_C249_n797);
   mult_21_C249_U1237 : MUXB2DL port map( A0 => N3209, A1 => N3210, SL => 
                           mult_21_C249_n1377, Z => mult_21_C249_n798);
   mult_21_C249_U1236 : MUXB2DL port map( A0 => N3208, A1 => N3209, SL => 
                           mult_21_C249_n1377, Z => mult_21_C249_n799);
   mult_21_C249_U1235 : MUXB2DL port map( A0 => N3207, A1 => N3208, SL => 
                           mult_21_C249_n1377, Z => mult_21_C249_n800);
   mult_21_C249_U1234 : MUXB2DL port map( A0 => N3206, A1 => N3207, SL => 
                           mult_21_C249_n1377, Z => mult_21_C249_n801);
   mult_21_C249_U1233 : MUXB2DL port map( A0 => N3205, A1 => mult_21_C249_n1385
                           , SL => mult_21_C249_n1377, Z => mult_21_C249_n802);
   mult_21_C249_U1232 : MUXB2DL port map( A0 => mult_21_C249_n1387, A1 => N3205
                           , SL => mult_21_C249_n1377, Z => mult_21_C249_n803);
   mult_21_C249_U1231 : MUXB2DL port map( A0 => N3203, A1 => N3204, SL => 
                           mult_21_C249_n1377, Z => mult_21_C249_n804);
   mult_21_C249_U1230 : MUXB2DL port map( A0 => N3202, A1 => mult_21_C249_n1389
                           , SL => mult_21_C249_n1377, Z => mult_21_C249_n805);
   mult_21_C249_U1229 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C249_n1377, Z => mult_21_C249_n806);
   mult_21_C249_U1228 : NAN2D1 port map( A1 => mult_21_C249_n1393, A2 => 
                           mult_21_C249_n1377, Z => mult_21_C249_n807);
   mult_21_C249_U1227 : MUXB2DL port map( A0 => N3225, A1 => N3226, SL => 
                           mult_21_C249_n1376, Z => mult_21_C249_n808);
   mult_21_C249_U1226 : MUXB2DL port map( A0 => N3224, A1 => N3225, SL => 
                           mult_21_C249_n1376, Z => mult_21_C249_n809);
   mult_21_C249_U1225 : AOI21D1 port map( A1 => N3060, A2 => N3061, B => 
                           mult_21_C249_n1416, Z => mult_21_C249_n944);
   mult_21_C249_U1224 : MUXB2DL port map( A0 => N3223, A1 => N3224, SL => 
                           mult_21_C249_n1376, Z => mult_21_C249_n810);
   mult_21_C249_U1223 : MUXB2DL port map( A0 => N3222, A1 => N3223, SL => 
                           mult_21_C249_n1376, Z => mult_21_C249_n811);
   mult_21_C249_U1222 : MUXB2DL port map( A0 => N3221, A1 => N3222, SL => 
                           mult_21_C249_n1376, Z => mult_21_C249_n812);
   mult_21_C249_U1221 : MUXB2DL port map( A0 => N3220, A1 => N3221, SL => 
                           mult_21_C249_n1376, Z => mult_21_C249_n813);
   mult_21_C249_U1220 : MUXB2DL port map( A0 => N3219, A1 => N3220, SL => 
                           mult_21_C249_n1376, Z => mult_21_C249_n814);
   mult_21_C249_U1219 : MUXB2DL port map( A0 => N3218, A1 => N3219, SL => 
                           mult_21_C249_n1376, Z => mult_21_C249_n815);
   mult_21_C249_U1218 : MUXB2DL port map( A0 => N3217, A1 => N3218, SL => 
                           mult_21_C249_n1376, Z => mult_21_C249_n816);
   mult_21_C249_U1217 : MUXB2DL port map( A0 => N3216, A1 => N3217, SL => 
                           mult_21_C249_n1376, Z => mult_21_C249_n817);
   mult_21_C249_U1216 : MUXB2DL port map( A0 => N3215, A1 => N3216, SL => 
                           mult_21_C249_n1376, Z => mult_21_C249_n818);
   mult_21_C249_U1215 : MUXB2DL port map( A0 => N3214, A1 => N3215, SL => 
                           mult_21_C249_n1376, Z => mult_21_C249_n819);
   mult_21_C249_U1214 : MUXB2DL port map( A0 => N3213, A1 => N3214, SL => 
                           mult_21_C249_n1376, Z => mult_21_C249_n820);
   mult_21_C249_U1213 : MUXB2DL port map( A0 => N3212, A1 => N3213, SL => 
                           mult_21_C249_n1376, Z => mult_21_C249_n821);
   mult_21_C249_U1212 : MUXB2DL port map( A0 => N3211, A1 => N3212, SL => 
                           mult_21_C249_n1376, Z => mult_21_C249_n822);
   mult_21_C249_U1211 : MUXB2DL port map( A0 => N3210, A1 => N3211, SL => 
                           mult_21_C249_n1376, Z => mult_21_C249_n823);
   mult_21_C249_U1210 : MUXB2DL port map( A0 => N3209, A1 => N3210, SL => 
                           mult_21_C249_n1376, Z => mult_21_C249_n824);
   mult_21_C249_U1209 : MUXB2DL port map( A0 => N3208, A1 => N3209, SL => 
                           mult_21_C249_n1376, Z => mult_21_C249_n825);
   mult_21_C249_U1208 : MUXB2DL port map( A0 => N3207, A1 => N3208, SL => 
                           mult_21_C249_n1376, Z => mult_21_C249_n826);
   mult_21_C249_U1207 : MUXB2DL port map( A0 => N3206, A1 => N3207, SL => 
                           mult_21_C249_n1376, Z => mult_21_C249_n827);
   mult_21_C249_U1206 : MUXB2DL port map( A0 => N3205, A1 => mult_21_C249_n1385
                           , SL => mult_21_C249_n1376, Z => mult_21_C249_n828);
   mult_21_C249_U1205 : MUXB2DL port map( A0 => mult_21_C249_n1387, A1 => N3205
                           , SL => mult_21_C249_n1376, Z => mult_21_C249_n829);
   mult_21_C249_U1204 : MUXB2DL port map( A0 => mult_21_C249_n1389, A1 => N3204
                           , SL => mult_21_C249_n1376, Z => mult_21_C249_n830);
   mult_21_C249_U1203 : MUXB2DL port map( A0 => mult_21_C249_n1391, A1 => 
                           mult_21_C249_n1389, SL => mult_21_C249_n1376, Z => 
                           mult_21_C249_n831);
   mult_21_C249_U1202 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C249_n1376, Z => mult_21_C249_n832);
   mult_21_C249_U1201 : NAN2D1 port map( A1 => mult_21_C249_n1393, A2 => 
                           mult_21_C249_n1376, Z => mult_21_C249_n833);
   mult_21_C249_U1200 : MUXB2DL port map( A0 => N3227, A1 => N3228, SL => 
                           mult_21_C249_n1375, Z => mult_21_C249_n834);
   mult_21_C249_U1199 : MUXB2DL port map( A0 => N3226, A1 => N3227, SL => 
                           mult_21_C249_n1375, Z => mult_21_C249_n835);
   mult_21_C249_U1198 : MUXB2DL port map( A0 => N3225, A1 => N3226, SL => 
                           mult_21_C249_n1375, Z => mult_21_C249_n836);
   mult_21_C249_U1197 : MUXB2DL port map( A0 => N3224, A1 => N3225, SL => 
                           mult_21_C249_n1375, Z => mult_21_C249_n837);
   mult_21_C249_U1196 : MUXB2DL port map( A0 => N3223, A1 => N3224, SL => 
                           mult_21_C249_n1375, Z => mult_21_C249_n838);
   mult_21_C249_U1195 : MUXB2DL port map( A0 => N3222, A1 => N3223, SL => 
                           mult_21_C249_n1375, Z => mult_21_C249_n839);
   mult_21_C249_U1194 : MUXB2DL port map( A0 => N3221, A1 => N3222, SL => 
                           mult_21_C249_n1375, Z => mult_21_C249_n840);
   mult_21_C249_U1193 : MUXB2DL port map( A0 => N3220, A1 => N3221, SL => 
                           mult_21_C249_n1375, Z => mult_21_C249_n841);
   mult_21_C249_U1192 : MUXB2DL port map( A0 => N3219, A1 => N3220, SL => 
                           mult_21_C249_n1375, Z => mult_21_C249_n842);
   mult_21_C249_U1191 : MUXB2DL port map( A0 => N3218, A1 => N3219, SL => 
                           mult_21_C249_n1375, Z => mult_21_C249_n843);
   mult_21_C249_U1190 : MUXB2DL port map( A0 => N3217, A1 => N3218, SL => 
                           mult_21_C249_n1375, Z => mult_21_C249_n844);
   mult_21_C249_U1189 : MUXB2DL port map( A0 => N3216, A1 => N3217, SL => 
                           mult_21_C249_n1375, Z => mult_21_C249_n845);
   mult_21_C249_U1188 : MUXB2DL port map( A0 => N3215, A1 => N3216, SL => 
                           mult_21_C249_n1375, Z => mult_21_C249_n846);
   mult_21_C249_U1187 : MUXB2DL port map( A0 => N3214, A1 => N3215, SL => 
                           mult_21_C249_n1375, Z => mult_21_C249_n847);
   mult_21_C249_U1186 : MUXB2DL port map( A0 => N3213, A1 => N3214, SL => 
                           mult_21_C249_n1375, Z => mult_21_C249_n848);
   mult_21_C249_U1185 : MUXB2DL port map( A0 => N3212, A1 => N3213, SL => 
                           mult_21_C249_n1375, Z => mult_21_C249_n849);
   mult_21_C249_U1184 : MUXB2DL port map( A0 => N3211, A1 => N3212, SL => 
                           mult_21_C249_n1375, Z => mult_21_C249_n850);
   mult_21_C249_U1183 : MUXB2DL port map( A0 => N3210, A1 => N3211, SL => 
                           mult_21_C249_n1375, Z => mult_21_C249_n851);
   mult_21_C249_U1182 : MUXB2DL port map( A0 => N3209, A1 => N3210, SL => 
                           mult_21_C249_n1375, Z => mult_21_C249_n852);
   mult_21_C249_U1181 : MUXB2DL port map( A0 => N3208, A1 => N3209, SL => 
                           mult_21_C249_n1375, Z => mult_21_C249_n853);
   mult_21_C249_U1180 : MUXB2DL port map( A0 => N3207, A1 => N3208, SL => 
                           mult_21_C249_n1375, Z => mult_21_C249_n854);
   mult_21_C249_U1179 : MUXB2DL port map( A0 => N3206, A1 => N3207, SL => 
                           mult_21_C249_n1375, Z => mult_21_C249_n855);
   mult_21_C249_U1178 : MUXB2DL port map( A0 => N3205, A1 => mult_21_C249_n1385
                           , SL => mult_21_C249_n1375, Z => mult_21_C249_n856);
   mult_21_C249_U1177 : MUXB2DL port map( A0 => mult_21_C249_n1387, A1 => N3205
                           , SL => mult_21_C249_n1375, Z => mult_21_C249_n857);
   mult_21_C249_U1176 : MUXB2DL port map( A0 => N3203, A1 => N3204, SL => 
                           mult_21_C249_n1375, Z => mult_21_C249_n858);
   mult_21_C249_U1175 : MUXB2DL port map( A0 => mult_21_C249_n1391, A1 => 
                           mult_21_C249_n1389, SL => mult_21_C249_n1375, Z => 
                           mult_21_C249_n859);
   mult_21_C249_U1174 : AOI21D1 port map( A1 => N3062, A2 => N3063, B => 
                           mult_21_C249_n1418, Z => mult_21_C249_n943);
   mult_21_C249_U1173 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C249_n1375, Z => mult_21_C249_n860);
   mult_21_C249_U1172 : NAN2D1 port map( A1 => mult_21_C249_n1393, A2 => 
                           mult_21_C249_n1375, Z => mult_21_C249_n861);
   mult_21_C249_U1171 : MUXB2DL port map( A0 => N3228, A1 => N3229, SL => 
                           mult_21_C249_n1384, Z => mult_21_C249_n863);
   mult_21_C249_U1170 : MUXB2DL port map( A0 => N3227, A1 => N3228, SL => 
                           mult_21_C249_n1384, Z => mult_21_C249_n864);
   mult_21_C249_U1169 : MUXB2DL port map( A0 => N3226, A1 => N3227, SL => 
                           mult_21_C249_n1384, Z => mult_21_C249_n865);
   mult_21_C249_U1168 : MUXB2DL port map( A0 => N3225, A1 => N3226, SL => 
                           mult_21_C249_n1384, Z => mult_21_C249_n866);
   mult_21_C249_U1167 : MUXB2DL port map( A0 => N3224, A1 => N3225, SL => 
                           mult_21_C249_n1384, Z => mult_21_C249_n867);
   mult_21_C249_U1166 : MUXB2DL port map( A0 => N3223, A1 => N3224, SL => 
                           mult_21_C249_n1384, Z => mult_21_C249_n868);
   mult_21_C249_U1165 : MUXB2DL port map( A0 => N3222, A1 => N3223, SL => 
                           mult_21_C249_n1384, Z => mult_21_C249_n869);
   mult_21_C249_U1164 : MUXB2DL port map( A0 => N3221, A1 => N3222, SL => 
                           mult_21_C249_n1384, Z => mult_21_C249_n870);
   mult_21_C249_U1163 : MUXB2DL port map( A0 => N3220, A1 => N3221, SL => 
                           mult_21_C249_n1384, Z => mult_21_C249_n871);
   mult_21_C249_U1162 : MUXB2DL port map( A0 => N3219, A1 => N3220, SL => 
                           mult_21_C249_n1384, Z => mult_21_C249_n872);
   mult_21_C249_U1161 : MUXB2DL port map( A0 => N3218, A1 => N3219, SL => 
                           mult_21_C249_n1384, Z => mult_21_C249_n873);
   mult_21_C249_U1160 : MUXB2DL port map( A0 => N3217, A1 => N3218, SL => 
                           mult_21_C249_n1384, Z => mult_21_C249_n874);
   mult_21_C249_U1159 : MUXB2DL port map( A0 => N3216, A1 => N3217, SL => 
                           mult_21_C249_n1384, Z => mult_21_C249_n875);
   mult_21_C249_U1158 : MUXB2DL port map( A0 => N3215, A1 => N3216, SL => 
                           mult_21_C249_n1384, Z => mult_21_C249_n876);
   mult_21_C249_U1157 : MUXB2DL port map( A0 => N3214, A1 => N3215, SL => 
                           mult_21_C249_n1384, Z => mult_21_C249_n877);
   mult_21_C249_U1156 : MUXB2DL port map( A0 => N3213, A1 => N3214, SL => 
                           mult_21_C249_n1384, Z => mult_21_C249_n878);
   mult_21_C249_U1155 : MUXB2DL port map( A0 => N3212, A1 => N3213, SL => 
                           mult_21_C249_n1384, Z => mult_21_C249_n879);
   mult_21_C249_U1154 : MUXB2DL port map( A0 => N3211, A1 => N3212, SL => 
                           mult_21_C249_n1384, Z => mult_21_C249_n880);
   mult_21_C249_U1153 : MUXB2DL port map( A0 => N3210, A1 => N3211, SL => 
                           mult_21_C249_n1384, Z => mult_21_C249_n881);
   mult_21_C249_U1152 : MUXB2DL port map( A0 => N3209, A1 => N3210, SL => 
                           mult_21_C249_n1384, Z => mult_21_C249_n882);
   mult_21_C249_U1151 : MUXB2DL port map( A0 => N3208, A1 => N3209, SL => 
                           mult_21_C249_n1384, Z => mult_21_C249_n883);
   mult_21_C249_U1150 : MUXB2DL port map( A0 => N3207, A1 => N3208, SL => 
                           mult_21_C249_n1384, Z => mult_21_C249_n884);
   mult_21_C249_U1149 : MUXB2DL port map( A0 => N3206, A1 => N3207, SL => 
                           mult_21_C249_n1384, Z => mult_21_C249_n885);
   mult_21_C249_U1148 : MUXB2DL port map( A0 => N3205, A1 => mult_21_C249_n1385
                           , SL => mult_21_C249_n1384, Z => mult_21_C249_n886);
   mult_21_C249_U1147 : MUXB2DL port map( A0 => mult_21_C249_n1387, A1 => N3205
                           , SL => mult_21_C249_n1384, Z => mult_21_C249_n887);
   mult_21_C249_U1146 : MUXB2DL port map( A0 => N3203, A1 => N3204, SL => 
                           mult_21_C249_n1384, Z => mult_21_C249_n888);
   mult_21_C249_U1145 : MUXB2DL port map( A0 => mult_21_C249_n1391, A1 => 
                           mult_21_C249_n1389, SL => mult_21_C249_n1384, Z => 
                           mult_21_C249_n889);
   mult_21_C249_U1144 : OAI21D1 port map( A1 => N3065, A2 => N3064, B => 
                           mult_21_C249_n1420, Z => mult_21_C249_n89);
   mult_21_C249_U1143 : MUXB2DL port map( A0 => N3201, A1 => N3202, SL => 
                           mult_21_C249_n1384, Z => mult_21_C249_n890);
   mult_21_C249_U1142 : NAN2D1 port map( A1 => mult_21_C249_n1393, A2 => 
                           mult_21_C249_n1384, Z => mult_21_C249_n891);
   mult_21_C249_U1141 : MUXB2DL port map( A0 => N3231, A1 => N3232, SL => N3041
                           , Z => mult_21_C249_n892);
   mult_21_C249_U1140 : MUXB2DL port map( A0 => N3230, A1 => N3231, SL => N3041
                           , Z => mult_21_C249_n893);
   mult_21_C249_U1139 : MUXB2DL port map( A0 => N3229, A1 => N3230, SL => N3041
                           , Z => mult_21_C249_n894);
   mult_21_C249_U1138 : MUXB2DL port map( A0 => N3228, A1 => N3229, SL => N3041
                           , Z => mult_21_C249_n895);
   mult_21_C249_U1137 : MUXB2DL port map( A0 => N3227, A1 => N3228, SL => N3041
                           , Z => mult_21_C249_n896);
   mult_21_C249_U1136 : MUXB2DL port map( A0 => N3226, A1 => N3227, SL => N3041
                           , Z => mult_21_C249_n897);
   mult_21_C249_U1135 : MUXB2DL port map( A0 => N3225, A1 => N3226, SL => N3041
                           , Z => mult_21_C249_n898);
   mult_21_C249_U1134 : MUXB2DL port map( A0 => N3224, A1 => N3225, SL => N3041
                           , Z => mult_21_C249_n899);
   mult_21_C249_U1133 : MUXB2DL port map( A0 => N3223, A1 => N3224, SL => N3041
                           , Z => mult_21_C249_n900);
   mult_21_C249_U1132 : MUXB2DL port map( A0 => N3222, A1 => N3223, SL => N3041
                           , Z => mult_21_C249_n901);
   mult_21_C249_U1131 : MUXB2DL port map( A0 => N3221, A1 => N3222, SL => N3041
                           , Z => mult_21_C249_n902);
   mult_21_C249_U1130 : MUXB2DL port map( A0 => N3220, A1 => N3221, SL => N3041
                           , Z => mult_21_C249_n903);
   mult_21_C249_U1129 : MUXB2DL port map( A0 => N3219, A1 => N3220, SL => N3041
                           , Z => mult_21_C249_n904);
   mult_21_C249_U1128 : MUXB2DL port map( A0 => N3218, A1 => N3219, SL => N3041
                           , Z => mult_21_C249_n905);
   mult_21_C249_U1127 : MUXB2DL port map( A0 => N3217, A1 => N3218, SL => N3041
                           , Z => mult_21_C249_n906);
   mult_21_C249_U1126 : MUXB2DL port map( A0 => N3216, A1 => N3217, SL => N3041
                           , Z => mult_21_C249_n907);
   mult_21_C249_U1125 : MUXB2DL port map( A0 => N3215, A1 => N3216, SL => N3041
                           , Z => mult_21_C249_n908);
   mult_21_C249_U1124 : MUXB2DL port map( A0 => N3214, A1 => N3215, SL => N3041
                           , Z => mult_21_C249_n909);
   mult_21_C249_U1123 : AOI21D1 port map( A1 => N3064, A2 => N3065, B => 
                           mult_21_C249_n1420, Z => mult_21_C249_n942);
   mult_21_C249_U1122 : MUXB2DL port map( A0 => N3213, A1 => N3214, SL => N3041
                           , Z => mult_21_C249_n910);
   mult_21_C249_U1121 : MUXB2DL port map( A0 => N3212, A1 => N3213, SL => N3041
                           , Z => mult_21_C249_n911);
   mult_21_C249_U1120 : MUXB2DL port map( A0 => N3211, A1 => N3212, SL => N3041
                           , Z => mult_21_C249_n912);
   mult_21_C249_U1119 : MUXB2DL port map( A0 => N3210, A1 => N3211, SL => N3041
                           , Z => mult_21_C249_n913);
   mult_21_C249_U1118 : MUXB2DL port map( A0 => N3209, A1 => N3210, SL => N3041
                           , Z => mult_21_C249_n914);
   mult_21_C249_U1117 : MUXB2DL port map( A0 => N3208, A1 => N3209, SL => N3041
                           , Z => mult_21_C249_n915);
   mult_21_C249_U1116 : MUXB2DL port map( A0 => N3207, A1 => N3208, SL => N3041
                           , Z => mult_21_C249_n916);
   mult_21_C249_U1115 : MUXB2DL port map( A0 => mult_21_C249_n1385, A1 => N3207
                           , SL => N3041, Z => mult_21_C249_n917);
   mult_21_C249_U1114 : MUXB2DL port map( A0 => N3205, A1 => mult_21_C249_n1385
                           , SL => N3041, Z => mult_21_C249_n918);
   mult_21_C249_U1113 : MUXB2DL port map( A0 => mult_21_C249_n1387, A1 => N3205
                           , SL => N3041, Z => mult_21_C249_n919);
   mult_21_C249_U1112 : MUXB2DL port map( A0 => N3203, A1 => mult_21_C249_n1387
                           , SL => N3041, Z => mult_21_C249_n920);
   mult_21_C249_U1111 : MUXB2DL port map( A0 => mult_21_C249_n1391, A1 => 
                           mult_21_C249_n1389, SL => N3041, Z => 
                           mult_21_C249_n921);
   mult_21_C249_U1110 : MUXB2DL port map( A0 => N3201, A1 => mult_21_C249_n1391
                           , SL => N3041, Z => mult_21_C249_n922);
   mult_21_C249_U1109 : NAN2D1 port map( A1 => mult_21_C249_n1393, A2 => N3041,
                           Z => mult_21_C249_n923);
   mult_21_C249_U1108 : OAI21D1 port map( A1 => N3067, A2 => N3066, B => 
                           mult_21_C249_n1421, Z => mult_21_C249_n94);
   mult_21_C249_U1107 : AOI21D1 port map( A1 => N3066, A2 => N3067, B => 
                           mult_21_C249_n1421, Z => mult_21_C249_n941);
   mult_21_C249_U1106 : OAI21D1 port map( A1 => N3069, A2 => N3068, B => 
                           mult_21_C249_n1424, Z => mult_21_C249_n99);
   mult_21_C249_U1105 : EXOR2D1 port map( A1 => mult_21_C249_n230, A2 => 
                           mult_21_C249_n228, Z => mult_21_C249_n1443);
   mult_21_C249_U1104 : EXOR3D1 port map( A1 => mult_21_C249_n226, A2 => 
                           mult_21_C249_n224, A3 => mult_21_C249_n1443, Z => 
                           mult_21_C249_n1438);
   mult_21_C249_U1103 : EXOR2D1 port map( A1 => mult_21_C249_n222, A2 => 
                           mult_21_C249_n220, Z => mult_21_C249_n1442);
   mult_21_C249_U1102 : EXOR3D1 port map( A1 => mult_21_C249_n216, A2 => 
                           mult_21_C249_n1195, A3 => mult_21_C249_n1442, Z => 
                           mult_21_C249_n1439);
   mult_21_C249_U1101 : EXOR3D1 port map( A1 => mult_21_C249_n1165, A2 => 
                           mult_21_C249_n1137, A3 => mult_21_C249_n1045, Z => 
                           mult_21_C249_n1441);
   mult_21_C249_U1100 : EXOR3D1 port map( A1 => mult_21_C249_n1027, A2 => 
                           mult_21_C249_n1011, A3 => mult_21_C249_n1441, Z => 
                           mult_21_C249_n1440);
   mult_21_C249_U1099 : EXOR3D1 port map( A1 => mult_21_C249_n1438, A2 => 
                           mult_21_C249_n1439, A3 => mult_21_C249_n1440, Z => 
                           mult_21_C249_n1430);
   mult_21_C249_U1098 : EXOR2D1 port map( A1 => mult_21_C249_n985, A2 => 
                           mult_21_C249_n967, Z => mult_21_C249_n1437);
   mult_21_C249_U1097 : EXOR3D1 port map( A1 => mult_21_C249_n961, A2 => 
                           mult_21_C249_n218, A3 => mult_21_C249_n1437, Z => 
                           mult_21_C249_n1434);
   mult_21_C249_U1096 : EXNOR2D1 port map( A1 => mult_21_C249_n210, A2 => 
                           mult_21_C249_n1111, Z => mult_21_C249_n1436);
   mult_21_C249_U1095 : EXOR3D1 port map( A1 => mult_21_C249_n1087, A2 => 
                           mult_21_C249_n1065, A3 => mult_21_C249_n1436, Z => 
                           mult_21_C249_n1435);
   mult_21_C249_U1094 : EXOR3D1 port map( A1 => mult_21_C249_n1434, A2 => 
                           mult_21_C249_n204, A3 => mult_21_C249_n1435, Z => 
                           mult_21_C249_n1431);
   mult_21_C249_U1093 : EXNOR2D1 port map( A1 => mult_21_C249_n997, A2 => 
                           mult_21_C249_n975, Z => mult_21_C249_n1433);
   mult_21_C249_U1092 : EXOR3D1 port map( A1 => mult_21_C249_n957, A2 => 
                           mult_21_C249_n955, A3 => mult_21_C249_n1433, Z => 
                           mult_21_C249_n1432);
   mult_21_C249_U1091 : EXOR3D1 port map( A1 => mult_21_C249_n1430, A2 => 
                           mult_21_C249_n1431, A3 => mult_21_C249_n1432, Z => 
                           mult_21_C249_n1426);
   mult_21_C249_U1090 : EXOR2D1 port map( A1 => mult_21_C249_n202, A2 => 
                           mult_21_C249_n156, Z => mult_21_C249_n1427);
   mult_21_C249_U1089 : EXOR2D1 port map( A1 => mult_21_C249_n214, A2 => 
                           mult_21_C249_n212, Z => mult_21_C249_n1429);
   mult_21_C249_U1088 : EXOR3D1 port map( A1 => mult_21_C249_n208, A2 => 
                           mult_21_C249_n206, A3 => mult_21_C249_n1429, Z => 
                           mult_21_C249_n1428);
   mult_21_C249_U1087 : EXOR3D1 port map( A1 => mult_21_C249_n1426, A2 => 
                           mult_21_C249_n1427, A3 => mult_21_C249_n1428, Z => 
                           N3392);
   mult_21_C249_U1086 : INVD1 port map( A => N3072, Z => mult_21_C249_n1425);
   mult_21_C249_U1085 : MUXB2DL port map( A0 => N3230, A1 => N3229, SL => 
                           mult_21_C249_n1383, Z => mult_21_C249_n862);
   mult_21_C249_U1084 : INVD1 port map( A => N3070, Z => mult_21_C249_n1424);
   mult_21_C249_U1083 : INVD1 port map( A => N3068, Z => mult_21_C249_n1421);
   mult_21_C249_U1082 : INVD1 port map( A => N3066, Z => mult_21_C249_n1420);
   mult_21_C249_U1081 : OAI21D1 port map( A1 => N3063, A2 => N3062, B => 
                           mult_21_C249_n1418, Z => mult_21_C249_n84);
   mult_21_C249_U1080 : INVD1 port map( A => N3064, Z => mult_21_C249_n1418);
   mult_21_C249_U1079 : EXOR2D1 port map( A1 => N3063, A2 => N3062, Z => 
                           mult_21_C249_n1450);
   mult_21_C249_U1078 : OAI21D1 port map( A1 => N3061, A2 => N3060, B => 
                           mult_21_C249_n1416, Z => mult_21_C249_n80);
   mult_21_C249_U1077 : INVD1 port map( A => N3062, Z => mult_21_C249_n1416);
   mult_21_C249_U1076 : EXOR2D1 port map( A1 => N3061, A2 => N3060, Z => 
                           mult_21_C249_n1449);
   mult_21_C249_U1075 : OAI21D1 port map( A1 => N3059, A2 => N3058, B => 
                           mult_21_C249_n1414, Z => mult_21_C249_n73);
   mult_21_C249_U1074 : INVD1 port map( A => N3060, Z => mult_21_C249_n1414);
   mult_21_C249_U1073 : EXOR2D1 port map( A1 => N3059, A2 => N3058, Z => 
                           mult_21_C249_n1448);
   mult_21_C249_U1072 : OAI21D1 port map( A1 => N3057, A2 => N3056, B => 
                           mult_21_C249_n1412, Z => mult_21_C249_n66);
   mult_21_C249_U1071 : INVD1 port map( A => N3058, Z => mult_21_C249_n1412);
   mult_21_C249_U1070 : EXOR2D1 port map( A1 => N3057, A2 => N3056, Z => 
                           mult_21_C249_n1447);
   mult_21_C249_U1069 : OAI21D1 port map( A1 => N3055, A2 => N3054, B => 
                           mult_21_C249_n1410, Z => mult_21_C249_n58);
   mult_21_C249_U1068 : INVD1 port map( A => N3056, Z => mult_21_C249_n1410);
   mult_21_C249_U1067 : EXOR2D1 port map( A1 => N3055, A2 => N3054, Z => 
                           mult_21_C249_n1446);
   mult_21_C249_U1066 : OAI21D1 port map( A1 => N3053, A2 => N3052, B => 
                           mult_21_C249_n1408, Z => mult_21_C249_n50);
   mult_21_C249_U1065 : INVD1 port map( A => N3054, Z => mult_21_C249_n1408);
   mult_21_C249_U1064 : EXOR2D1 port map( A1 => N3053, A2 => N3052, Z => 
                           mult_21_C249_n1445);
   mult_21_C249_U1063 : OAI21D1 port map( A1 => N3050, A2 => N3051, B => 
                           mult_21_C249_n1406, Z => mult_21_C249_n42);
   mult_21_C249_U1062 : INVD1 port map( A => N3052, Z => mult_21_C249_n1406);
   mult_21_C249_U1061 : EXOR2D1 port map( A1 => N3051, A2 => N3050, Z => 
                           mult_21_C249_n1444);
   mult_21_C249_U1060 : INVD1 port map( A => N3050, Z => mult_21_C249_n1404);
   mult_21_C249_U1059 : INVD1 port map( A => N3048, Z => mult_21_C249_n1402);
   mult_21_C249_U1058 : INVD1 port map( A => N3206, Z => mult_21_C249_n1386);
   mult_21_C249_U1057 : INVD1 port map( A => N3046, Z => mult_21_C249_n1400);
   mult_21_C249_U1056 : INVD1 port map( A => N3044, Z => mult_21_C249_n1398);
   mult_21_C249_U1055 : INVD1 port map( A => N3204, Z => mult_21_C249_n1388);
   mult_21_C249_U1054 : INVD1 port map( A => N3201, Z => mult_21_C249_n1394);
   mult_21_C249_U1053 : INVD1 port map( A => N3202, Z => mult_21_C249_n1392);
   mult_21_C249_U1052 : INVD1 port map( A => N3203, Z => mult_21_C249_n1390);
   mult_21_C249_U1051 : EXNOR2D1 port map( A1 => N3043, A2 => N3042, Z => 
                           mult_21_C249_n1383);
   mult_21_C249_U1050 : INVD1 port map( A => N3042, Z => mult_21_C249_n1395);
   mult_21_C249_U1049 : INVD1 port map( A => mult_21_C249_n939, Z => 
                           mult_21_C249_n1423);
   mult_21_C249_U1048 : INVD1 port map( A => mult_21_C249_n940, Z => 
                           mult_21_C249_n1422);
   mult_21_C249_U1047 : INVD1 port map( A => mult_21_C249_n941, Z => 
                           mult_21_C249_n1419);
   mult_21_C249_U1046 : INVD1 port map( A => mult_21_C249_n942, Z => 
                           mult_21_C249_n1417);
   mult_21_C249_U1045 : INVD1 port map( A => mult_21_C249_n943, Z => 
                           mult_21_C249_n1415);
   mult_21_C249_U1044 : INVD1 port map( A => mult_21_C249_n944, Z => 
                           mult_21_C249_n1413);
   mult_21_C249_U1043 : INVD1 port map( A => mult_21_C249_n945, Z => 
                           mult_21_C249_n1411);
   mult_21_C249_U1042 : INVD1 port map( A => mult_21_C249_n946, Z => 
                           mult_21_C249_n1409);
   mult_21_C249_U1041 : INVD1 port map( A => mult_21_C249_n947, Z => 
                           mult_21_C249_n1407);
   mult_21_C249_U1040 : INVD1 port map( A => mult_21_C249_n948, Z => 
                           mult_21_C249_n1405);
   mult_21_C249_U1039 : INVD1 port map( A => mult_21_C249_n949, Z => 
                           mult_21_C249_n1403);
   mult_21_C249_U1038 : INVD1 port map( A => mult_21_C249_n950, Z => 
                           mult_21_C249_n1401);
   mult_21_C249_U1037 : INVD1 port map( A => mult_21_C249_n951, Z => 
                           mult_21_C249_n1399);
   mult_21_C249_U1036 : INVD1 port map( A => mult_21_C249_n952, Z => 
                           mult_21_C249_n1397);
   mult_21_C249_U1035 : INVD1 port map( A => mult_21_C249_n1386, Z => 
                           mult_21_C249_n1385);
   mult_21_C249_U1034 : INVD1 port map( A => mult_21_C249_n953, Z => 
                           mult_21_C249_n1396);
   mult_21_C249_U1033 : INVD1 port map( A => mult_21_C249_n1388, Z => 
                           mult_21_C249_n1387);
   mult_21_C249_U1032 : INVD1 port map( A => mult_21_C249_n1394, Z => 
                           mult_21_C249_n1393);
   mult_21_C249_U1031 : INVD1 port map( A => mult_21_C249_n1392, Z => 
                           mult_21_C249_n1391);
   mult_21_C249_U1030 : INVD1 port map( A => mult_21_C249_n1390, Z => 
                           mult_21_C249_n1389);
   mult_21_C249_U1029 : INVD1 port map( A => mult_21_C249_n1383, Z => 
                           mult_21_C249_n1384);
   mult_21_C249_U1028 : OAI21D1 port map( A1 => N3049, A2 => N3048, B => 
                           mult_21_C249_n1404, Z => mult_21_C249_n1382);
   mult_21_C249_U1027 : OAI21D1 port map( A1 => N3047, A2 => N3046, B => 
                           mult_21_C249_n1402, Z => mult_21_C249_n1381);
   mult_21_C249_U1026 : OAI21D1 port map( A1 => N3045, A2 => N3044, B => 
                           mult_21_C249_n1400, Z => mult_21_C249_n1380);
   mult_21_C249_U1025 : OAI21D1 port map( A1 => N3043, A2 => N3042, B => 
                           mult_21_C249_n1398, Z => mult_21_C249_n1379);
   mult_21_C249_U1024 : NAN2D1 port map( A1 => N3041, A2 => mult_21_C249_n1395,
                           Z => mult_21_C249_n1378);
   mult_21_C249_U1023 : EXOR2D1 port map( A1 => N3049, A2 => N3048, Z => 
                           mult_21_C249_n1377);
   mult_21_C249_U1022 : EXOR2D1 port map( A1 => N3047, A2 => N3046, Z => 
                           mult_21_C249_n1376);
   mult_21_C249_U1021 : EXOR2D1 port map( A1 => N3045, A2 => N3044, Z => 
                           mult_21_C249_n1375);
   mult_21_C249_U954 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n923, Z => 
                           mult_21_C249_n1226);
   mult_21_C249_U952 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n922, Z => 
                           mult_21_C249_n1225);
   mult_21_C249_U950 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n921, Z => 
                           mult_21_C249_n1224);
   mult_21_C249_U948 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n920, Z => 
                           mult_21_C249_n1223);
   mult_21_C249_U946 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n919, Z => 
                           mult_21_C249_n1222);
   mult_21_C249_U944 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n918, Z => 
                           mult_21_C249_n1221);
   mult_21_C249_U942 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n917, Z => 
                           mult_21_C249_n1220);
   mult_21_C249_U940 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n916, Z => 
                           mult_21_C249_n1219);
   mult_21_C249_U938 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n915, Z => 
                           mult_21_C249_n1218);
   mult_21_C249_U936 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n914, Z => 
                           mult_21_C249_n1217);
   mult_21_C249_U934 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n913, Z => 
                           mult_21_C249_n1216);
   mult_21_C249_U932 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n912, Z => 
                           mult_21_C249_n1215);
   mult_21_C249_U930 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n911, Z => 
                           mult_21_C249_n1214);
   mult_21_C249_U928 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n910, Z => 
                           mult_21_C249_n1213);
   mult_21_C249_U926 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n909, Z => 
                           mult_21_C249_n1212);
   mult_21_C249_U924 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n908, Z => 
                           mult_21_C249_n1211);
   mult_21_C249_U922 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n907, Z => 
                           mult_21_C249_n1210);
   mult_21_C249_U920 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n906, Z => 
                           mult_21_C249_n1209);
   mult_21_C249_U918 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n905, Z => 
                           mult_21_C249_n1208);
   mult_21_C249_U916 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n904, Z => 
                           mult_21_C249_n1207);
   mult_21_C249_U914 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n903, Z => 
                           mult_21_C249_n1206);
   mult_21_C249_U912 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n902, Z => 
                           mult_21_C249_n1205);
   mult_21_C249_U910 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n901, Z => 
                           mult_21_C249_n1204);
   mult_21_C249_U908 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n900, Z => 
                           mult_21_C249_n1203);
   mult_21_C249_U906 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n899, Z => 
                           mult_21_C249_n1202);
   mult_21_C249_U904 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n898, Z => 
                           mult_21_C249_n1201);
   mult_21_C249_U902 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n897, Z => 
                           mult_21_C249_n1200);
   mult_21_C249_U900 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n896, Z => 
                           mult_21_C249_n1199);
   mult_21_C249_U898 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n895, Z => 
                           mult_21_C249_n1198);
   mult_21_C249_U896 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n894, Z => 
                           mult_21_C249_n1197);
   mult_21_C249_U894 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n893, Z => 
                           mult_21_C249_n1196);
   mult_21_C249_U892 : MUXB2DL port map( A0 => mult_21_C249_n1378, A1 => 
                           mult_21_C249_n1395, SL => mult_21_C249_n892, Z => 
                           mult_21_C249_n1195);
   mult_21_C249_U889 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n891, Z => 
                           mult_21_C249_n1194);
   mult_21_C249_U887 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n890, Z => 
                           mult_21_C249_n1193);
   mult_21_C249_U885 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n889, Z => 
                           mult_21_C249_n1192);
   mult_21_C249_U883 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n888, Z => 
                           mult_21_C249_n1191);
   mult_21_C249_U881 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n887, Z => 
                           mult_21_C249_n1190);
   mult_21_C249_U879 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n886, Z => 
                           mult_21_C249_n1189);
   mult_21_C249_U877 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n885, Z => 
                           mult_21_C249_n1188);
   mult_21_C249_U875 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n884, Z => 
                           mult_21_C249_n1187);
   mult_21_C249_U873 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n883, Z => 
                           mult_21_C249_n1186);
   mult_21_C249_U871 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n882, Z => 
                           mult_21_C249_n1185);
   mult_21_C249_U869 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n881, Z => 
                           mult_21_C249_n1184);
   mult_21_C249_U867 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n880, Z => 
                           mult_21_C249_n1183);
   mult_21_C249_U865 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n879, Z => 
                           mult_21_C249_n1182);
   mult_21_C249_U863 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n878, Z => 
                           mult_21_C249_n1181);
   mult_21_C249_U861 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n877, Z => 
                           mult_21_C249_n1180);
   mult_21_C249_U859 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n876, Z => 
                           mult_21_C249_n1179);
   mult_21_C249_U857 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n875, Z => 
                           mult_21_C249_n1178);
   mult_21_C249_U855 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n874, Z => 
                           mult_21_C249_n1177);
   mult_21_C249_U853 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n873, Z => 
                           mult_21_C249_n1176);
   mult_21_C249_U851 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n872, Z => 
                           mult_21_C249_n1175);
   mult_21_C249_U849 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n871, Z => 
                           mult_21_C249_n1174);
   mult_21_C249_U847 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n870, Z => 
                           mult_21_C249_n1173);
   mult_21_C249_U845 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n869, Z => 
                           mult_21_C249_n1172);
   mult_21_C249_U843 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n868, Z => 
                           mult_21_C249_n1171);
   mult_21_C249_U841 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n867, Z => 
                           mult_21_C249_n1170);
   mult_21_C249_U839 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n866, Z => 
                           mult_21_C249_n1169);
   mult_21_C249_U837 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n865, Z => 
                           mult_21_C249_n1168);
   mult_21_C249_U835 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n864, Z => 
                           mult_21_C249_n1167);
   mult_21_C249_U833 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n863, Z => 
                           mult_21_C249_n1166);
   mult_21_C249_U831 : MUXB2DL port map( A0 => mult_21_C249_n1379, A1 => 
                           mult_21_C249_n1396, SL => mult_21_C249_n862, Z => 
                           mult_21_C249_n1165);
   mult_21_C249_U828 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n861, Z => 
                           mult_21_C249_n1164);
   mult_21_C249_U826 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n860, Z => 
                           mult_21_C249_n1163);
   mult_21_C249_U824 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n859, Z => 
                           mult_21_C249_n1162);
   mult_21_C249_U822 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n858, Z => 
                           mult_21_C249_n1161);
   mult_21_C249_U820 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n857, Z => 
                           mult_21_C249_n1160);
   mult_21_C249_U818 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n856, Z => 
                           mult_21_C249_n1159);
   mult_21_C249_U816 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n855, Z => 
                           mult_21_C249_n1158);
   mult_21_C249_U814 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n854, Z => 
                           mult_21_C249_n1157);
   mult_21_C249_U812 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n853, Z => 
                           mult_21_C249_n1156);
   mult_21_C249_U810 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n852, Z => 
                           mult_21_C249_n1155);
   mult_21_C249_U808 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n851, Z => 
                           mult_21_C249_n1154);
   mult_21_C249_U806 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n850, Z => 
                           mult_21_C249_n1153);
   mult_21_C249_U804 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n849, Z => 
                           mult_21_C249_n1152);
   mult_21_C249_U802 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n848, Z => 
                           mult_21_C249_n1151);
   mult_21_C249_U800 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n847, Z => 
                           mult_21_C249_n1150);
   mult_21_C249_U798 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n846, Z => 
                           mult_21_C249_n1149);
   mult_21_C249_U796 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n845, Z => 
                           mult_21_C249_n1148);
   mult_21_C249_U794 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n844, Z => 
                           mult_21_C249_n1147);
   mult_21_C249_U792 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n843, Z => 
                           mult_21_C249_n1146);
   mult_21_C249_U790 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n842, Z => 
                           mult_21_C249_n1145);
   mult_21_C249_U788 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n841, Z => 
                           mult_21_C249_n1144);
   mult_21_C249_U786 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n840, Z => 
                           mult_21_C249_n1143);
   mult_21_C249_U784 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n839, Z => 
                           mult_21_C249_n1142);
   mult_21_C249_U782 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n838, Z => 
                           mult_21_C249_n1141);
   mult_21_C249_U780 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n837, Z => 
                           mult_21_C249_n1140);
   mult_21_C249_U778 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n836, Z => 
                           mult_21_C249_n1139);
   mult_21_C249_U776 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n835, Z => 
                           mult_21_C249_n1138);
   mult_21_C249_U774 : MUXB2DL port map( A0 => mult_21_C249_n1380, A1 => 
                           mult_21_C249_n1397, SL => mult_21_C249_n834, Z => 
                           mult_21_C249_n1137);
   mult_21_C249_U771 : MUXB2DL port map( A0 => mult_21_C249_n1381, A1 => 
                           mult_21_C249_n1399, SL => mult_21_C249_n833, Z => 
                           mult_21_C249_n1136);
   mult_21_C249_U769 : MUXB2DL port map( A0 => mult_21_C249_n1381, A1 => 
                           mult_21_C249_n1399, SL => mult_21_C249_n832, Z => 
                           mult_21_C249_n1135);
   mult_21_C249_U767 : MUXB2DL port map( A0 => mult_21_C249_n1381, A1 => 
                           mult_21_C249_n1399, SL => mult_21_C249_n831, Z => 
                           mult_21_C249_n1134);
   mult_21_C249_U765 : MUXB2DL port map( A0 => mult_21_C249_n1381, A1 => 
                           mult_21_C249_n1399, SL => mult_21_C249_n830, Z => 
                           mult_21_C249_n1133);
   mult_21_C249_U763 : MUXB2DL port map( A0 => mult_21_C249_n1381, A1 => 
                           mult_21_C249_n1399, SL => mult_21_C249_n829, Z => 
                           mult_21_C249_n1132);
   mult_21_C249_U761 : MUXB2DL port map( A0 => mult_21_C249_n1381, A1 => 
                           mult_21_C249_n1399, SL => mult_21_C249_n828, Z => 
                           mult_21_C249_n1131);
   mult_21_C249_U759 : MUXB2DL port map( A0 => mult_21_C249_n1381, A1 => 
                           mult_21_C249_n1399, SL => mult_21_C249_n827, Z => 
                           mult_21_C249_n1130);
   mult_21_C249_U757 : MUXB2DL port map( A0 => mult_21_C249_n1381, A1 => 
                           mult_21_C249_n1399, SL => mult_21_C249_n826, Z => 
                           mult_21_C249_n1129);
   mult_21_C249_U755 : MUXB2DL port map( A0 => mult_21_C249_n1381, A1 => 
                           mult_21_C249_n1399, SL => mult_21_C249_n825, Z => 
                           mult_21_C249_n1128);
   mult_21_C249_U753 : MUXB2DL port map( A0 => mult_21_C249_n1381, A1 => 
                           mult_21_C249_n1399, SL => mult_21_C249_n824, Z => 
                           mult_21_C249_n1127);
   mult_21_C249_U751 : MUXB2DL port map( A0 => mult_21_C249_n1381, A1 => 
                           mult_21_C249_n1399, SL => mult_21_C249_n823, Z => 
                           mult_21_C249_n1126);
   mult_21_C249_U749 : MUXB2DL port map( A0 => mult_21_C249_n1381, A1 => 
                           mult_21_C249_n1399, SL => mult_21_C249_n822, Z => 
                           mult_21_C249_n1125);
   mult_21_C249_U747 : MUXB2DL port map( A0 => mult_21_C249_n1381, A1 => 
                           mult_21_C249_n1399, SL => mult_21_C249_n821, Z => 
                           mult_21_C249_n1124);
   mult_21_C249_U745 : MUXB2DL port map( A0 => mult_21_C249_n1381, A1 => 
                           mult_21_C249_n1399, SL => mult_21_C249_n820, Z => 
                           mult_21_C249_n1123);
   mult_21_C249_U743 : MUXB2DL port map( A0 => mult_21_C249_n1381, A1 => 
                           mult_21_C249_n1399, SL => mult_21_C249_n819, Z => 
                           mult_21_C249_n1122);
   mult_21_C249_U741 : MUXB2DL port map( A0 => mult_21_C249_n1381, A1 => 
                           mult_21_C249_n1399, SL => mult_21_C249_n818, Z => 
                           mult_21_C249_n1121);
   mult_21_C249_U739 : MUXB2DL port map( A0 => mult_21_C249_n1381, A1 => 
                           mult_21_C249_n1399, SL => mult_21_C249_n817, Z => 
                           mult_21_C249_n1120);
   mult_21_C249_U737 : MUXB2DL port map( A0 => mult_21_C249_n1381, A1 => 
                           mult_21_C249_n1399, SL => mult_21_C249_n816, Z => 
                           mult_21_C249_n1119);
   mult_21_C249_U735 : MUXB2DL port map( A0 => mult_21_C249_n1381, A1 => 
                           mult_21_C249_n1399, SL => mult_21_C249_n815, Z => 
                           mult_21_C249_n1118);
   mult_21_C249_U733 : MUXB2DL port map( A0 => mult_21_C249_n1381, A1 => 
                           mult_21_C249_n1399, SL => mult_21_C249_n814, Z => 
                           mult_21_C249_n1117);
   mult_21_C249_U731 : MUXB2DL port map( A0 => mult_21_C249_n1381, A1 => 
                           mult_21_C249_n1399, SL => mult_21_C249_n813, Z => 
                           mult_21_C249_n1116);
   mult_21_C249_U729 : MUXB2DL port map( A0 => mult_21_C249_n1381, A1 => 
                           mult_21_C249_n1399, SL => mult_21_C249_n812, Z => 
                           mult_21_C249_n1115);
   mult_21_C249_U727 : MUXB2DL port map( A0 => mult_21_C249_n1381, A1 => 
                           mult_21_C249_n1399, SL => mult_21_C249_n811, Z => 
                           mult_21_C249_n1114);
   mult_21_C249_U725 : MUXB2DL port map( A0 => mult_21_C249_n1381, A1 => 
                           mult_21_C249_n1399, SL => mult_21_C249_n810, Z => 
                           mult_21_C249_n1113);
   mult_21_C249_U723 : MUXB2DL port map( A0 => mult_21_C249_n1381, A1 => 
                           mult_21_C249_n1399, SL => mult_21_C249_n809, Z => 
                           mult_21_C249_n1112);
   mult_21_C249_U721 : MUXB2DL port map( A0 => mult_21_C249_n1381, A1 => 
                           mult_21_C249_n1399, SL => mult_21_C249_n808, Z => 
                           mult_21_C249_n1111);
   mult_21_C249_U718 : MUXB2DL port map( A0 => mult_21_C249_n1382, A1 => 
                           mult_21_C249_n1401, SL => mult_21_C249_n807, Z => 
                           mult_21_C249_n1110);
   mult_21_C249_U716 : MUXB2DL port map( A0 => mult_21_C249_n1382, A1 => 
                           mult_21_C249_n1401, SL => mult_21_C249_n806, Z => 
                           mult_21_C249_n1109);
   mult_21_C249_U714 : MUXB2DL port map( A0 => mult_21_C249_n1382, A1 => 
                           mult_21_C249_n1401, SL => mult_21_C249_n805, Z => 
                           mult_21_C249_n1108);
   mult_21_C249_U712 : MUXB2DL port map( A0 => mult_21_C249_n1382, A1 => 
                           mult_21_C249_n1401, SL => mult_21_C249_n804, Z => 
                           mult_21_C249_n1107);
   mult_21_C249_U710 : MUXB2DL port map( A0 => mult_21_C249_n1382, A1 => 
                           mult_21_C249_n1401, SL => mult_21_C249_n803, Z => 
                           mult_21_C249_n1106);
   mult_21_C249_U708 : MUXB2DL port map( A0 => mult_21_C249_n1382, A1 => 
                           mult_21_C249_n1401, SL => mult_21_C249_n802, Z => 
                           mult_21_C249_n1105);
   mult_21_C249_U706 : MUXB2DL port map( A0 => mult_21_C249_n1382, A1 => 
                           mult_21_C249_n1401, SL => mult_21_C249_n801, Z => 
                           mult_21_C249_n1104);
   mult_21_C249_U704 : MUXB2DL port map( A0 => mult_21_C249_n1382, A1 => 
                           mult_21_C249_n1401, SL => mult_21_C249_n800, Z => 
                           mult_21_C249_n1103);
   mult_21_C249_U702 : MUXB2DL port map( A0 => mult_21_C249_n1382, A1 => 
                           mult_21_C249_n1401, SL => mult_21_C249_n799, Z => 
                           mult_21_C249_n1102);
   mult_21_C249_U700 : MUXB2DL port map( A0 => mult_21_C249_n1382, A1 => 
                           mult_21_C249_n1401, SL => mult_21_C249_n798, Z => 
                           mult_21_C249_n1101);
   mult_21_C249_U698 : MUXB2DL port map( A0 => mult_21_C249_n1382, A1 => 
                           mult_21_C249_n1401, SL => mult_21_C249_n797, Z => 
                           mult_21_C249_n1100);
   mult_21_C249_U696 : MUXB2DL port map( A0 => mult_21_C249_n1382, A1 => 
                           mult_21_C249_n1401, SL => mult_21_C249_n796, Z => 
                           mult_21_C249_n1099);
   mult_21_C249_U694 : MUXB2DL port map( A0 => mult_21_C249_n1382, A1 => 
                           mult_21_C249_n1401, SL => mult_21_C249_n795, Z => 
                           mult_21_C249_n1098);
   mult_21_C249_U692 : MUXB2DL port map( A0 => mult_21_C249_n1382, A1 => 
                           mult_21_C249_n1401, SL => mult_21_C249_n794, Z => 
                           mult_21_C249_n1097);
   mult_21_C249_U690 : MUXB2DL port map( A0 => mult_21_C249_n1382, A1 => 
                           mult_21_C249_n1401, SL => mult_21_C249_n793, Z => 
                           mult_21_C249_n1096);
   mult_21_C249_U688 : MUXB2DL port map( A0 => mult_21_C249_n1382, A1 => 
                           mult_21_C249_n1401, SL => mult_21_C249_n792, Z => 
                           mult_21_C249_n1095);
   mult_21_C249_U686 : MUXB2DL port map( A0 => mult_21_C249_n1382, A1 => 
                           mult_21_C249_n1401, SL => mult_21_C249_n791, Z => 
                           mult_21_C249_n1094);
   mult_21_C249_U684 : MUXB2DL port map( A0 => mult_21_C249_n1382, A1 => 
                           mult_21_C249_n1401, SL => mult_21_C249_n790, Z => 
                           mult_21_C249_n1093);
   mult_21_C249_U682 : MUXB2DL port map( A0 => mult_21_C249_n1382, A1 => 
                           mult_21_C249_n1401, SL => mult_21_C249_n789, Z => 
                           mult_21_C249_n1092);
   mult_21_C249_U680 : MUXB2DL port map( A0 => mult_21_C249_n1382, A1 => 
                           mult_21_C249_n1401, SL => mult_21_C249_n788, Z => 
                           mult_21_C249_n1091);
   mult_21_C249_U678 : MUXB2DL port map( A0 => mult_21_C249_n1382, A1 => 
                           mult_21_C249_n1401, SL => mult_21_C249_n787, Z => 
                           mult_21_C249_n1090);
   mult_21_C249_U676 : MUXB2DL port map( A0 => mult_21_C249_n1382, A1 => 
                           mult_21_C249_n1401, SL => mult_21_C249_n786, Z => 
                           mult_21_C249_n1089);
   mult_21_C249_U674 : MUXB2DL port map( A0 => mult_21_C249_n1382, A1 => 
                           mult_21_C249_n1401, SL => mult_21_C249_n785, Z => 
                           mult_21_C249_n1088);
   mult_21_C249_U672 : MUXB2DL port map( A0 => mult_21_C249_n1382, A1 => 
                           mult_21_C249_n1401, SL => mult_21_C249_n784, Z => 
                           mult_21_C249_n1087);
   mult_21_C249_U669 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n1403, SL => mult_21_C249_n783, Z => 
                           mult_21_C249_n1086);
   mult_21_C249_U667 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n1403, SL => mult_21_C249_n782, Z => 
                           mult_21_C249_n1085);
   mult_21_C249_U665 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n1403, SL => mult_21_C249_n781, Z => 
                           mult_21_C249_n1084);
   mult_21_C249_U663 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n1403, SL => mult_21_C249_n780, Z => 
                           mult_21_C249_n1083);
   mult_21_C249_U661 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n1403, SL => mult_21_C249_n779, Z => 
                           mult_21_C249_n1082);
   mult_21_C249_U659 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n1403, SL => mult_21_C249_n778, Z => 
                           mult_21_C249_n1081);
   mult_21_C249_U657 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n1403, SL => mult_21_C249_n777, Z => 
                           mult_21_C249_n1080);
   mult_21_C249_U655 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n1403, SL => mult_21_C249_n776, Z => 
                           mult_21_C249_n1079);
   mult_21_C249_U653 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n1403, SL => mult_21_C249_n775, Z => 
                           mult_21_C249_n1078);
   mult_21_C249_U651 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n1403, SL => mult_21_C249_n774, Z => 
                           mult_21_C249_n1077);
   mult_21_C249_U649 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n1403, SL => mult_21_C249_n773, Z => 
                           mult_21_C249_n1076);
   mult_21_C249_U647 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n1403, SL => mult_21_C249_n772, Z => 
                           mult_21_C249_n1075);
   mult_21_C249_U645 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n1403, SL => mult_21_C249_n771, Z => 
                           mult_21_C249_n1074);
   mult_21_C249_U643 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n1403, SL => mult_21_C249_n770, Z => 
                           mult_21_C249_n1073);
   mult_21_C249_U641 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n1403, SL => mult_21_C249_n769, Z => 
                           mult_21_C249_n1072);
   mult_21_C249_U639 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n1403, SL => mult_21_C249_n768, Z => 
                           mult_21_C249_n1071);
   mult_21_C249_U637 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n1403, SL => mult_21_C249_n767, Z => 
                           mult_21_C249_n1070);
   mult_21_C249_U635 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n1403, SL => mult_21_C249_n766, Z => 
                           mult_21_C249_n1069);
   mult_21_C249_U633 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n1403, SL => mult_21_C249_n765, Z => 
                           mult_21_C249_n1068);
   mult_21_C249_U631 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n1403, SL => mult_21_C249_n764, Z => 
                           mult_21_C249_n1067);
   mult_21_C249_U629 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n1403, SL => mult_21_C249_n763, Z => 
                           mult_21_C249_n1066);
   mult_21_C249_U627 : MUXB2DL port map( A0 => mult_21_C249_n42, A1 => 
                           mult_21_C249_n1403, SL => mult_21_C249_n762, Z => 
                           mult_21_C249_n1065);
   mult_21_C249_U624 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n1405, SL => mult_21_C249_n761, Z => 
                           mult_21_C249_n1064);
   mult_21_C249_U622 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n1405, SL => mult_21_C249_n760, Z => 
                           mult_21_C249_n1063);
   mult_21_C249_U620 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n1405, SL => mult_21_C249_n759, Z => 
                           mult_21_C249_n1062);
   mult_21_C249_U618 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n1405, SL => mult_21_C249_n758, Z => 
                           mult_21_C249_n1061);
   mult_21_C249_U616 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n1405, SL => mult_21_C249_n757, Z => 
                           mult_21_C249_n1060);
   mult_21_C249_U614 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n1405, SL => mult_21_C249_n756, Z => 
                           mult_21_C249_n1059);
   mult_21_C249_U612 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n1405, SL => mult_21_C249_n755, Z => 
                           mult_21_C249_n1058);
   mult_21_C249_U610 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n1405, SL => mult_21_C249_n754, Z => 
                           mult_21_C249_n1057);
   mult_21_C249_U608 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n1405, SL => mult_21_C249_n753, Z => 
                           mult_21_C249_n1056);
   mult_21_C249_U606 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n1405, SL => mult_21_C249_n752, Z => 
                           mult_21_C249_n1055);
   mult_21_C249_U604 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n1405, SL => mult_21_C249_n751, Z => 
                           mult_21_C249_n1054);
   mult_21_C249_U602 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n1405, SL => mult_21_C249_n750, Z => 
                           mult_21_C249_n1053);
   mult_21_C249_U600 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n1405, SL => mult_21_C249_n749, Z => 
                           mult_21_C249_n1052);
   mult_21_C249_U598 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n1405, SL => mult_21_C249_n748, Z => 
                           mult_21_C249_n1051);
   mult_21_C249_U596 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n1405, SL => mult_21_C249_n747, Z => 
                           mult_21_C249_n1050);
   mult_21_C249_U594 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n1405, SL => mult_21_C249_n746, Z => 
                           mult_21_C249_n1049);
   mult_21_C249_U592 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n1405, SL => mult_21_C249_n745, Z => 
                           mult_21_C249_n1048);
   mult_21_C249_U590 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n1405, SL => mult_21_C249_n744, Z => 
                           mult_21_C249_n1047);
   mult_21_C249_U588 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n1405, SL => mult_21_C249_n743, Z => 
                           mult_21_C249_n1046);
   mult_21_C249_U586 : MUXB2DL port map( A0 => mult_21_C249_n50, A1 => 
                           mult_21_C249_n1405, SL => mult_21_C249_n742, Z => 
                           mult_21_C249_n1045);
   mult_21_C249_U583 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n1407, SL => mult_21_C249_n741, Z => 
                           mult_21_C249_n1044);
   mult_21_C249_U581 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n1407, SL => mult_21_C249_n740, Z => 
                           mult_21_C249_n1043);
   mult_21_C249_U579 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n1407, SL => mult_21_C249_n739, Z => 
                           mult_21_C249_n1042);
   mult_21_C249_U577 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n1407, SL => mult_21_C249_n738, Z => 
                           mult_21_C249_n1041);
   mult_21_C249_U575 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n1407, SL => mult_21_C249_n737, Z => 
                           mult_21_C249_n1040);
   mult_21_C249_U573 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n1407, SL => mult_21_C249_n736, Z => 
                           mult_21_C249_n1039);
   mult_21_C249_U571 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n1407, SL => mult_21_C249_n735, Z => 
                           mult_21_C249_n1038);
   mult_21_C249_U569 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n1407, SL => mult_21_C249_n734, Z => 
                           mult_21_C249_n1037);
   mult_21_C249_U567 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n1407, SL => mult_21_C249_n733, Z => 
                           mult_21_C249_n1036);
   mult_21_C249_U565 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n1407, SL => mult_21_C249_n732, Z => 
                           mult_21_C249_n1035);
   mult_21_C249_U563 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n1407, SL => mult_21_C249_n731, Z => 
                           mult_21_C249_n1034);
   mult_21_C249_U561 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n1407, SL => mult_21_C249_n730, Z => 
                           mult_21_C249_n1033);
   mult_21_C249_U559 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n1407, SL => mult_21_C249_n729, Z => 
                           mult_21_C249_n1032);
   mult_21_C249_U557 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n1407, SL => mult_21_C249_n728, Z => 
                           mult_21_C249_n1031);
   mult_21_C249_U555 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n1407, SL => mult_21_C249_n727, Z => 
                           mult_21_C249_n1030);
   mult_21_C249_U553 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n1407, SL => mult_21_C249_n726, Z => 
                           mult_21_C249_n1029);
   mult_21_C249_U551 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n1407, SL => mult_21_C249_n725, Z => 
                           mult_21_C249_n1028);
   mult_21_C249_U549 : MUXB2DL port map( A0 => mult_21_C249_n58, A1 => 
                           mult_21_C249_n1407, SL => mult_21_C249_n724, Z => 
                           mult_21_C249_n1027);
   mult_21_C249_U546 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n1409, SL => mult_21_C249_n723, Z => 
                           mult_21_C249_n1026);
   mult_21_C249_U544 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n1409, SL => mult_21_C249_n722, Z => 
                           mult_21_C249_n1025);
   mult_21_C249_U542 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n1409, SL => mult_21_C249_n721, Z => 
                           mult_21_C249_n1024);
   mult_21_C249_U540 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n1409, SL => mult_21_C249_n720, Z => 
                           mult_21_C249_n1023);
   mult_21_C249_U538 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n1409, SL => mult_21_C249_n719, Z => 
                           mult_21_C249_n1022);
   mult_21_C249_U536 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n1409, SL => mult_21_C249_n718, Z => 
                           mult_21_C249_n1021);
   mult_21_C249_U534 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n1409, SL => mult_21_C249_n717, Z => 
                           mult_21_C249_n1020);
   mult_21_C249_U532 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n1409, SL => mult_21_C249_n716, Z => 
                           mult_21_C249_n1019);
   mult_21_C249_U530 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n1409, SL => mult_21_C249_n715, Z => 
                           mult_21_C249_n1018);
   mult_21_C249_U528 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n1409, SL => mult_21_C249_n714, Z => 
                           mult_21_C249_n1017);
   mult_21_C249_U526 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n1409, SL => mult_21_C249_n713, Z => 
                           mult_21_C249_n1016);
   mult_21_C249_U524 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n1409, SL => mult_21_C249_n712, Z => 
                           mult_21_C249_n1015);
   mult_21_C249_U522 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n1409, SL => mult_21_C249_n711, Z => 
                           mult_21_C249_n1014);
   mult_21_C249_U520 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n1409, SL => mult_21_C249_n710, Z => 
                           mult_21_C249_n1013);
   mult_21_C249_U518 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n1409, SL => mult_21_C249_n709, Z => 
                           mult_21_C249_n1012);
   mult_21_C249_U516 : MUXB2DL port map( A0 => mult_21_C249_n66, A1 => 
                           mult_21_C249_n1409, SL => mult_21_C249_n708, Z => 
                           mult_21_C249_n1011);
   mult_21_C249_U513 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n1411, SL => mult_21_C249_n707, Z => 
                           mult_21_C249_n1010);
   mult_21_C249_U511 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n1411, SL => mult_21_C249_n706, Z => 
                           mult_21_C249_n1009);
   mult_21_C249_U509 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n1411, SL => mult_21_C249_n705, Z => 
                           mult_21_C249_n1008);
   mult_21_C249_U507 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n1411, SL => mult_21_C249_n704, Z => 
                           mult_21_C249_n1007);
   mult_21_C249_U505 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n1411, SL => mult_21_C249_n703, Z => 
                           mult_21_C249_n1006);
   mult_21_C249_U503 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n1411, SL => mult_21_C249_n702, Z => 
                           mult_21_C249_n1005);
   mult_21_C249_U501 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n1411, SL => mult_21_C249_n701, Z => 
                           mult_21_C249_n1004);
   mult_21_C249_U499 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n1411, SL => mult_21_C249_n700, Z => 
                           mult_21_C249_n1003);
   mult_21_C249_U497 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n1411, SL => mult_21_C249_n699, Z => 
                           mult_21_C249_n1002);
   mult_21_C249_U495 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n1411, SL => mult_21_C249_n698, Z => 
                           mult_21_C249_n1001);
   mult_21_C249_U493 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n1411, SL => mult_21_C249_n697, Z => 
                           mult_21_C249_n1000);
   mult_21_C249_U491 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n1411, SL => mult_21_C249_n696, Z => 
                           mult_21_C249_n999);
   mult_21_C249_U489 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n1411, SL => mult_21_C249_n695, Z => 
                           mult_21_C249_n998);
   mult_21_C249_U487 : MUXB2DL port map( A0 => mult_21_C249_n73, A1 => 
                           mult_21_C249_n1411, SL => mult_21_C249_n694, Z => 
                           mult_21_C249_n997);
   mult_21_C249_U484 : MUXB2DL port map( A0 => mult_21_C249_n80, A1 => 
                           mult_21_C249_n1413, SL => mult_21_C249_n693, Z => 
                           mult_21_C249_n996);
   mult_21_C249_U482 : MUXB2DL port map( A0 => mult_21_C249_n80, A1 => 
                           mult_21_C249_n1413, SL => mult_21_C249_n692, Z => 
                           mult_21_C249_n995);
   mult_21_C249_U480 : MUXB2DL port map( A0 => mult_21_C249_n80, A1 => 
                           mult_21_C249_n1413, SL => mult_21_C249_n691, Z => 
                           mult_21_C249_n994);
   mult_21_C249_U478 : MUXB2DL port map( A0 => mult_21_C249_n80, A1 => 
                           mult_21_C249_n1413, SL => mult_21_C249_n690, Z => 
                           mult_21_C249_n993);
   mult_21_C249_U476 : MUXB2DL port map( A0 => mult_21_C249_n80, A1 => 
                           mult_21_C249_n1413, SL => mult_21_C249_n689, Z => 
                           mult_21_C249_n992);
   mult_21_C249_U474 : MUXB2DL port map( A0 => mult_21_C249_n80, A1 => 
                           mult_21_C249_n1413, SL => mult_21_C249_n688, Z => 
                           mult_21_C249_n991);
   mult_21_C249_U472 : MUXB2DL port map( A0 => mult_21_C249_n80, A1 => 
                           mult_21_C249_n1413, SL => mult_21_C249_n687, Z => 
                           mult_21_C249_n990);
   mult_21_C249_U470 : MUXB2DL port map( A0 => mult_21_C249_n80, A1 => 
                           mult_21_C249_n1413, SL => mult_21_C249_n686, Z => 
                           mult_21_C249_n989);
   mult_21_C249_U468 : MUXB2DL port map( A0 => mult_21_C249_n80, A1 => 
                           mult_21_C249_n1413, SL => mult_21_C249_n685, Z => 
                           mult_21_C249_n988);
   mult_21_C249_U466 : MUXB2DL port map( A0 => mult_21_C249_n80, A1 => 
                           mult_21_C249_n1413, SL => mult_21_C249_n684, Z => 
                           mult_21_C249_n987);
   mult_21_C249_U464 : MUXB2DL port map( A0 => mult_21_C249_n80, A1 => 
                           mult_21_C249_n1413, SL => mult_21_C249_n683, Z => 
                           mult_21_C249_n986);
   mult_21_C249_U462 : MUXB2DL port map( A0 => mult_21_C249_n80, A1 => 
                           mult_21_C249_n1413, SL => mult_21_C249_n682, Z => 
                           mult_21_C249_n985);
   mult_21_C249_U459 : MUXB2DL port map( A0 => mult_21_C249_n84, A1 => 
                           mult_21_C249_n1415, SL => mult_21_C249_n681, Z => 
                           mult_21_C249_n984);
   mult_21_C249_U457 : MUXB2DL port map( A0 => mult_21_C249_n84, A1 => 
                           mult_21_C249_n1415, SL => mult_21_C249_n680, Z => 
                           mult_21_C249_n983);
   mult_21_C249_U455 : MUXB2DL port map( A0 => mult_21_C249_n84, A1 => 
                           mult_21_C249_n1415, SL => mult_21_C249_n679, Z => 
                           mult_21_C249_n982);
   mult_21_C249_U453 : MUXB2DL port map( A0 => mult_21_C249_n84, A1 => 
                           mult_21_C249_n1415, SL => mult_21_C249_n678, Z => 
                           mult_21_C249_n981);
   mult_21_C249_U451 : MUXB2DL port map( A0 => mult_21_C249_n84, A1 => 
                           mult_21_C249_n1415, SL => mult_21_C249_n677, Z => 
                           mult_21_C249_n980);
   mult_21_C249_U449 : MUXB2DL port map( A0 => mult_21_C249_n84, A1 => 
                           mult_21_C249_n1415, SL => mult_21_C249_n676, Z => 
                           mult_21_C249_n979);
   mult_21_C249_U447 : MUXB2DL port map( A0 => mult_21_C249_n84, A1 => 
                           mult_21_C249_n1415, SL => mult_21_C249_n675, Z => 
                           mult_21_C249_n978);
   mult_21_C249_U445 : MUXB2DL port map( A0 => mult_21_C249_n84, A1 => 
                           mult_21_C249_n1415, SL => mult_21_C249_n674, Z => 
                           mult_21_C249_n977);
   mult_21_C249_U443 : MUXB2DL port map( A0 => mult_21_C249_n84, A1 => 
                           mult_21_C249_n1415, SL => mult_21_C249_n673, Z => 
                           mult_21_C249_n976);
   mult_21_C249_U441 : MUXB2DL port map( A0 => mult_21_C249_n84, A1 => 
                           mult_21_C249_n1415, SL => mult_21_C249_n672, Z => 
                           mult_21_C249_n975);
   mult_21_C249_U438 : MUXB2DL port map( A0 => mult_21_C249_n89, A1 => 
                           mult_21_C249_n1417, SL => mult_21_C249_n671, Z => 
                           mult_21_C249_n974);
   mult_21_C249_U436 : MUXB2DL port map( A0 => mult_21_C249_n89, A1 => 
                           mult_21_C249_n1417, SL => mult_21_C249_n670, Z => 
                           mult_21_C249_n973);
   mult_21_C249_U434 : MUXB2DL port map( A0 => mult_21_C249_n89, A1 => 
                           mult_21_C249_n1417, SL => mult_21_C249_n669, Z => 
                           mult_21_C249_n972);
   mult_21_C249_U432 : MUXB2DL port map( A0 => mult_21_C249_n89, A1 => 
                           mult_21_C249_n1417, SL => mult_21_C249_n668, Z => 
                           mult_21_C249_n971);
   mult_21_C249_U430 : MUXB2DL port map( A0 => mult_21_C249_n89, A1 => 
                           mult_21_C249_n1417, SL => mult_21_C249_n667, Z => 
                           mult_21_C249_n970);
   mult_21_C249_U428 : MUXB2DL port map( A0 => mult_21_C249_n89, A1 => 
                           mult_21_C249_n1417, SL => mult_21_C249_n666, Z => 
                           mult_21_C249_n969);
   mult_21_C249_U426 : MUXB2DL port map( A0 => mult_21_C249_n89, A1 => 
                           mult_21_C249_n1417, SL => mult_21_C249_n665, Z => 
                           mult_21_C249_n968);
   mult_21_C249_U424 : MUXB2DL port map( A0 => mult_21_C249_n89, A1 => 
                           mult_21_C249_n1417, SL => mult_21_C249_n664, Z => 
                           mult_21_C249_n967);
   mult_21_C249_U421 : MUXB2DL port map( A0 => mult_21_C249_n94, A1 => 
                           mult_21_C249_n1419, SL => mult_21_C249_n663, Z => 
                           mult_21_C249_n966);
   mult_21_C249_U419 : MUXB2DL port map( A0 => mult_21_C249_n94, A1 => 
                           mult_21_C249_n1419, SL => mult_21_C249_n662, Z => 
                           mult_21_C249_n965);
   mult_21_C249_U417 : MUXB2DL port map( A0 => mult_21_C249_n94, A1 => 
                           mult_21_C249_n1419, SL => mult_21_C249_n661, Z => 
                           mult_21_C249_n964);
   mult_21_C249_U415 : MUXB2DL port map( A0 => mult_21_C249_n94, A1 => 
                           mult_21_C249_n1419, SL => mult_21_C249_n660, Z => 
                           mult_21_C249_n963);
   mult_21_C249_U413 : MUXB2DL port map( A0 => mult_21_C249_n94, A1 => 
                           mult_21_C249_n1419, SL => mult_21_C249_n659, Z => 
                           mult_21_C249_n962);
   mult_21_C249_U411 : MUXB2DL port map( A0 => mult_21_C249_n94, A1 => 
                           mult_21_C249_n1419, SL => mult_21_C249_n658, Z => 
                           mult_21_C249_n961);
   mult_21_C249_U408 : MUXB2DL port map( A0 => mult_21_C249_n99, A1 => 
                           mult_21_C249_n1422, SL => mult_21_C249_n657, Z => 
                           mult_21_C249_n960);
   mult_21_C249_U406 : MUXB2DL port map( A0 => mult_21_C249_n99, A1 => 
                           mult_21_C249_n1422, SL => mult_21_C249_n656, Z => 
                           mult_21_C249_n959);
   mult_21_C249_U404 : MUXB2DL port map( A0 => mult_21_C249_n99, A1 => 
                           mult_21_C249_n1422, SL => mult_21_C249_n655, Z => 
                           mult_21_C249_n958);
   mult_21_C249_U402 : MUXB2DL port map( A0 => mult_21_C249_n99, A1 => 
                           mult_21_C249_n1422, SL => mult_21_C249_n654, Z => 
                           mult_21_C249_n957);
   mult_21_C249_U399 : MUXB2DL port map( A0 => mult_21_C249_n104, A1 => 
                           mult_21_C249_n1423, SL => mult_21_C249_n653, Z => 
                           mult_21_C249_n956);
   mult_21_C249_U397 : MUXB2DL port map( A0 => mult_21_C249_n104, A1 => 
                           mult_21_C249_n1423, SL => mult_21_C249_n652, Z => 
                           mult_21_C249_n955);
   mult_21_C249_U395 : ADHALFDL port map( A => mult_21_C249_n1224, B => 
                           mult_21_C249_n953, CO => mult_21_C249_n650, S => 
                           mult_21_C249_n651);
   mult_21_C249_U394 : ADHALFDL port map( A => mult_21_C249_n650, B => 
                           mult_21_C249_n1223, CO => mult_21_C249_n648, S => 
                           mult_21_C249_n649);
   mult_21_C249_U393 : ADHALFDL port map( A => mult_21_C249_n1222, B => 
                           mult_21_C249_n952, CO => mult_21_C249_n646, S => 
                           mult_21_C249_n647);
   mult_21_C249_U392 : ADFULD1 port map( A => mult_21_C249_n1192, B => 
                           mult_21_C249_n1164, CI => mult_21_C249_n647, CO => 
                           mult_21_C249_n644, S => mult_21_C249_n645);
   mult_21_C249_U391 : ADHALFDL port map( A => mult_21_C249_n646, B => 
                           mult_21_C249_n1221, CO => mult_21_C249_n642, S => 
                           mult_21_C249_n643);
   mult_21_C249_U390 : ADFULD1 port map( A => mult_21_C249_n1163, B => 
                           mult_21_C249_n1191, CI => mult_21_C249_n643, CO => 
                           mult_21_C249_n640, S => mult_21_C249_n641);
   mult_21_C249_U389 : ADHALFDL port map( A => mult_21_C249_n1220, B => 
                           mult_21_C249_n951, CO => mult_21_C249_n638, S => 
                           mult_21_C249_n639);
   mult_21_C249_U388 : ADFULD1 port map( A => mult_21_C249_n1190, B => 
                           mult_21_C249_n1136, CI => mult_21_C249_n1162, CO => 
                           mult_21_C249_n636, S => mult_21_C249_n637);
   mult_21_C249_U387 : ADFULD1 port map( A => mult_21_C249_n642, B => 
                           mult_21_C249_n639, CI => mult_21_C249_n637, CO => 
                           mult_21_C249_n634, S => mult_21_C249_n635);
   mult_21_C249_U386 : ADHALFDL port map( A => mult_21_C249_n638, B => 
                           mult_21_C249_n1219, CO => mult_21_C249_n632, S => 
                           mult_21_C249_n633);
   mult_21_C249_U385 : ADFULD1 port map( A => mult_21_C249_n1135, B => 
                           mult_21_C249_n1189, CI => mult_21_C249_n1161, CO => 
                           mult_21_C249_n630, S => mult_21_C249_n631);
   mult_21_C249_U384 : ADFULD1 port map( A => mult_21_C249_n636, B => 
                           mult_21_C249_n633, CI => mult_21_C249_n631, CO => 
                           mult_21_C249_n628, S => mult_21_C249_n629);
   mult_21_C249_U383 : ADHALFDL port map( A => mult_21_C249_n1218, B => 
                           mult_21_C249_n950, CO => mult_21_C249_n626, S => 
                           mult_21_C249_n627);
   mult_21_C249_U382 : ADFULD1 port map( A => mult_21_C249_n1188, B => 
                           mult_21_C249_n1110, CI => mult_21_C249_n1134, CO => 
                           mult_21_C249_n624, S => mult_21_C249_n625);
   mult_21_C249_U381 : ADFULD1 port map( A => mult_21_C249_n627, B => 
                           mult_21_C249_n1160, CI => mult_21_C249_n632, CO => 
                           mult_21_C249_n622, S => mult_21_C249_n623);
   mult_21_C249_U380 : ADFULD1 port map( A => mult_21_C249_n625, B => 
                           mult_21_C249_n630, CI => mult_21_C249_n623, CO => 
                           mult_21_C249_n620, S => mult_21_C249_n621);
   mult_21_C249_U379 : ADHALFDL port map( A => mult_21_C249_n626, B => 
                           mult_21_C249_n1217, CO => mult_21_C249_n618, S => 
                           mult_21_C249_n619);
   mult_21_C249_U378 : ADFULD1 port map( A => mult_21_C249_n1109, B => 
                           mult_21_C249_n1133, CI => mult_21_C249_n1159, CO => 
                           mult_21_C249_n616, S => mult_21_C249_n617);
   mult_21_C249_U377 : ADFULD1 port map( A => mult_21_C249_n619, B => 
                           mult_21_C249_n1187, CI => mult_21_C249_n624, CO => 
                           mult_21_C249_n614, S => mult_21_C249_n615);
   mult_21_C249_U376 : ADFULD1 port map( A => mult_21_C249_n617, B => 
                           mult_21_C249_n622, CI => mult_21_C249_n615, CO => 
                           mult_21_C249_n612, S => mult_21_C249_n613);
   mult_21_C249_U375 : ADHALFDL port map( A => mult_21_C249_n1216, B => 
                           mult_21_C249_n949, CO => mult_21_C249_n610, S => 
                           mult_21_C249_n611);
   mult_21_C249_U374 : ADFULD1 port map( A => mult_21_C249_n1132, B => 
                           mult_21_C249_n1086, CI => mult_21_C249_n1186, CO => 
                           mult_21_C249_n608, S => mult_21_C249_n609);
   mult_21_C249_U373 : ADFULD1 port map( A => mult_21_C249_n1108, B => 
                           mult_21_C249_n1158, CI => mult_21_C249_n611, CO => 
                           mult_21_C249_n606, S => mult_21_C249_n607);
   mult_21_C249_U372 : ADFULD1 port map( A => mult_21_C249_n616, B => 
                           mult_21_C249_n618, CI => mult_21_C249_n609, CO => 
                           mult_21_C249_n604, S => mult_21_C249_n605);
   mult_21_C249_U371 : ADFULD1 port map( A => mult_21_C249_n614, B => 
                           mult_21_C249_n607, CI => mult_21_C249_n605, CO => 
                           mult_21_C249_n602, S => mult_21_C249_n603);
   mult_21_C249_U370 : ADHALFDL port map( A => mult_21_C249_n610, B => 
                           mult_21_C249_n1215, CO => mult_21_C249_n600, S => 
                           mult_21_C249_n601);
   mult_21_C249_U369 : ADFULD1 port map( A => mult_21_C249_n1085, B => 
                           mult_21_C249_n1131, CI => mult_21_C249_n1185, CO => 
                           mult_21_C249_n598, S => mult_21_C249_n599);
   mult_21_C249_U368 : ADFULD1 port map( A => mult_21_C249_n1107, B => 
                           mult_21_C249_n1157, CI => mult_21_C249_n601, CO => 
                           mult_21_C249_n596, S => mult_21_C249_n597);
   mult_21_C249_U367 : ADFULD1 port map( A => mult_21_C249_n606, B => 
                           mult_21_C249_n608, CI => mult_21_C249_n599, CO => 
                           mult_21_C249_n594, S => mult_21_C249_n595);
   mult_21_C249_U366 : ADFULD1 port map( A => mult_21_C249_n604, B => 
                           mult_21_C249_n597, CI => mult_21_C249_n595, CO => 
                           mult_21_C249_n592, S => mult_21_C249_n593);
   mult_21_C249_U365 : ADHALFDL port map( A => mult_21_C249_n1214, B => 
                           mult_21_C249_n948, CO => mult_21_C249_n590, S => 
                           mult_21_C249_n591);
   mult_21_C249_U364 : ADFULD1 port map( A => mult_21_C249_n1130, B => 
                           mult_21_C249_n1064, CI => mult_21_C249_n1184, CO => 
                           mult_21_C249_n588, S => mult_21_C249_n589);
   mult_21_C249_U363 : ADFULD1 port map( A => mult_21_C249_n1084, B => 
                           mult_21_C249_n1156, CI => mult_21_C249_n591, CO => 
                           mult_21_C249_n586, S => mult_21_C249_n587);
   mult_21_C249_U362 : ADFULD1 port map( A => mult_21_C249_n600, B => 
                           mult_21_C249_n1106, CI => mult_21_C249_n598, CO => 
                           mult_21_C249_n584, S => mult_21_C249_n585);
   mult_21_C249_U361 : ADFULD1 port map( A => mult_21_C249_n587, B => 
                           mult_21_C249_n589, CI => mult_21_C249_n596, CO => 
                           mult_21_C249_n582, S => mult_21_C249_n583);
   mult_21_C249_U360 : ADFULD1 port map( A => mult_21_C249_n585, B => 
                           mult_21_C249_n594, CI => mult_21_C249_n583, CO => 
                           mult_21_C249_n580, S => mult_21_C249_n581);
   mult_21_C249_U359 : ADHALFDL port map( A => mult_21_C249_n590, B => 
                           mult_21_C249_n1213, CO => mult_21_C249_n578, S => 
                           mult_21_C249_n579);
   mult_21_C249_U358 : ADFULD1 port map( A => mult_21_C249_n1183, B => 
                           mult_21_C249_n1105, CI => mult_21_C249_n1155, CO => 
                           mult_21_C249_n576, S => mult_21_C249_n577);
   mult_21_C249_U357 : ADFULD1 port map( A => mult_21_C249_n1063, B => 
                           mult_21_C249_n1129, CI => mult_21_C249_n1083, CO => 
                           mult_21_C249_n574, S => mult_21_C249_n575);
   mult_21_C249_U356 : ADFULD1 port map( A => mult_21_C249_n588, B => 
                           mult_21_C249_n579, CI => mult_21_C249_n586, CO => 
                           mult_21_C249_n572, S => mult_21_C249_n573);
   mult_21_C249_U355 : ADFULD1 port map( A => mult_21_C249_n577, B => 
                           mult_21_C249_n575, CI => mult_21_C249_n584, CO => 
                           mult_21_C249_n570, S => mult_21_C249_n571);
   mult_21_C249_U354 : ADFULD1 port map( A => mult_21_C249_n582, B => 
                           mult_21_C249_n573, CI => mult_21_C249_n571, CO => 
                           mult_21_C249_n568, S => mult_21_C249_n569);
   mult_21_C249_U353 : ADHALFDL port map( A => mult_21_C249_n1212, B => 
                           mult_21_C249_n947, CO => mult_21_C249_n566, S => 
                           mult_21_C249_n567);
   mult_21_C249_U352 : ADFULD1 port map( A => mult_21_C249_n1104, B => 
                           mult_21_C249_n1044, CI => mult_21_C249_n1182, CO => 
                           mult_21_C249_n564, S => mult_21_C249_n565);
   mult_21_C249_U351 : ADFULD1 port map( A => mult_21_C249_n1154, B => 
                           mult_21_C249_n1082, CI => mult_21_C249_n567, CO => 
                           mult_21_C249_n562, S => mult_21_C249_n563);
   mult_21_C249_U350 : ADFULD1 port map( A => mult_21_C249_n1062, B => 
                           mult_21_C249_n1128, CI => mult_21_C249_n578, CO => 
                           mult_21_C249_n560, S => mult_21_C249_n561);
   mult_21_C249_U349 : ADFULD1 port map( A => mult_21_C249_n574, B => 
                           mult_21_C249_n576, CI => mult_21_C249_n565, CO => 
                           mult_21_C249_n558, S => mult_21_C249_n559);
   mult_21_C249_U348 : ADFULD1 port map( A => mult_21_C249_n561, B => 
                           mult_21_C249_n563, CI => mult_21_C249_n572, CO => 
                           mult_21_C249_n556, S => mult_21_C249_n557);
   mult_21_C249_U347 : ADFULD1 port map( A => mult_21_C249_n570, B => 
                           mult_21_C249_n559, CI => mult_21_C249_n557, CO => 
                           mult_21_C249_n554, S => mult_21_C249_n555);
   mult_21_C249_U346 : ADHALFDL port map( A => mult_21_C249_n566, B => 
                           mult_21_C249_n1211, CO => mult_21_C249_n552, S => 
                           mult_21_C249_n553);
   mult_21_C249_U345 : ADFULD1 port map( A => mult_21_C249_n1043, B => 
                           mult_21_C249_n1103, CI => mult_21_C249_n1061, CO => 
                           mult_21_C249_n550, S => mult_21_C249_n551);
   mult_21_C249_U344 : ADFULD1 port map( A => mult_21_C249_n1181, B => 
                           mult_21_C249_n1081, CI => mult_21_C249_n1127, CO => 
                           mult_21_C249_n548, S => mult_21_C249_n549);
   mult_21_C249_U343 : ADFULD1 port map( A => mult_21_C249_n553, B => 
                           mult_21_C249_n1153, CI => mult_21_C249_n564, CO => 
                           mult_21_C249_n546, S => mult_21_C249_n547);
   mult_21_C249_U342 : ADFULD1 port map( A => mult_21_C249_n560, B => 
                           mult_21_C249_n562, CI => mult_21_C249_n549, CO => 
                           mult_21_C249_n544, S => mult_21_C249_n545);
   mult_21_C249_U341 : ADFULD1 port map( A => mult_21_C249_n547, B => 
                           mult_21_C249_n551, CI => mult_21_C249_n558, CO => 
                           mult_21_C249_n542, S => mult_21_C249_n543);
   mult_21_C249_U340 : ADFULD1 port map( A => mult_21_C249_n556, B => 
                           mult_21_C249_n545, CI => mult_21_C249_n543, CO => 
                           mult_21_C249_n540, S => mult_21_C249_n541);
   mult_21_C249_U339 : ADHALFDL port map( A => mult_21_C249_n1210, B => 
                           mult_21_C249_n946, CO => mult_21_C249_n538, S => 
                           mult_21_C249_n539);
   mult_21_C249_U338 : ADFULD1 port map( A => mult_21_C249_n1102, B => 
                           mult_21_C249_n1026, CI => mult_21_C249_n1180, CO => 
                           mult_21_C249_n536, S => mult_21_C249_n537);
   mult_21_C249_U337 : ADFULD1 port map( A => mult_21_C249_n1042, B => 
                           mult_21_C249_n1060, CI => mult_21_C249_n539, CO => 
                           mult_21_C249_n534, S => mult_21_C249_n535);
   mult_21_C249_U336 : ADFULD1 port map( A => mult_21_C249_n1080, B => 
                           mult_21_C249_n1152, CI => mult_21_C249_n1126, CO => 
                           mult_21_C249_n532, S => mult_21_C249_n533);
   mult_21_C249_U335 : ADFULD1 port map( A => mult_21_C249_n550, B => 
                           mult_21_C249_n552, CI => mult_21_C249_n548, CO => 
                           mult_21_C249_n530, S => mult_21_C249_n531);
   mult_21_C249_U334 : ADFULD1 port map( A => mult_21_C249_n533, B => 
                           mult_21_C249_n537, CI => mult_21_C249_n535, CO => 
                           mult_21_C249_n528, S => mult_21_C249_n529);
   mult_21_C249_U333 : ADFULD1 port map( A => mult_21_C249_n544, B => 
                           mult_21_C249_n546, CI => mult_21_C249_n531, CO => 
                           mult_21_C249_n526, S => mult_21_C249_n527);
   mult_21_C249_U332 : ADFULD1 port map( A => mult_21_C249_n542, B => 
                           mult_21_C249_n529, CI => mult_21_C249_n527, CO => 
                           mult_21_C249_n524, S => mult_21_C249_n525);
   mult_21_C249_U331 : ADHALFDL port map( A => mult_21_C249_n538, B => 
                           mult_21_C249_n1209, CO => mult_21_C249_n522, S => 
                           mult_21_C249_n523);
   mult_21_C249_U330 : ADFULD1 port map( A => mult_21_C249_n1179, B => 
                           mult_21_C249_n1079, CI => mult_21_C249_n1151, CO => 
                           mult_21_C249_n520, S => mult_21_C249_n521);
   mult_21_C249_U329 : ADFULD1 port map( A => mult_21_C249_n1025, B => 
                           mult_21_C249_n1041, CI => mult_21_C249_n1059, CO => 
                           mult_21_C249_n518, S => mult_21_C249_n519);
   mult_21_C249_U328 : ADFULD1 port map( A => mult_21_C249_n1101, B => 
                           mult_21_C249_n1125, CI => mult_21_C249_n523, CO => 
                           mult_21_C249_n516, S => mult_21_C249_n517);
   mult_21_C249_U327 : ADFULD1 port map( A => mult_21_C249_n534, B => 
                           mult_21_C249_n536, CI => mult_21_C249_n532, CO => 
                           mult_21_C249_n514, S => mult_21_C249_n515);
   mult_21_C249_U326 : ADFULD1 port map( A => mult_21_C249_n521, B => 
                           mult_21_C249_n519, CI => mult_21_C249_n517, CO => 
                           mult_21_C249_n512, S => mult_21_C249_n513);
   mult_21_C249_U325 : ADFULD1 port map( A => mult_21_C249_n528, B => 
                           mult_21_C249_n530, CI => mult_21_C249_n515, CO => 
                           mult_21_C249_n510, S => mult_21_C249_n511);
   mult_21_C249_U324 : ADFULD1 port map( A => mult_21_C249_n526, B => 
                           mult_21_C249_n513, CI => mult_21_C249_n511, CO => 
                           mult_21_C249_n508, S => mult_21_C249_n509);
   mult_21_C249_U323 : ADHALFDL port map( A => mult_21_C249_n1208, B => 
                           mult_21_C249_n945, CO => mult_21_C249_n506, S => 
                           mult_21_C249_n507);
   mult_21_C249_U322 : ADFULD1 port map( A => mult_21_C249_n1078, B => 
                           mult_21_C249_n1010, CI => mult_21_C249_n1024, CO => 
                           mult_21_C249_n504, S => mult_21_C249_n505);
   mult_21_C249_U321 : ADFULD1 port map( A => mult_21_C249_n1178, B => 
                           mult_21_C249_n1100, CI => mult_21_C249_n507, CO => 
                           mult_21_C249_n502, S => mult_21_C249_n503);
   mult_21_C249_U320 : ADFULD1 port map( A => mult_21_C249_n1040, B => 
                           mult_21_C249_n1150, CI => mult_21_C249_n1058, CO => 
                           mult_21_C249_n500, S => mult_21_C249_n501);
   mult_21_C249_U319 : ADFULD1 port map( A => mult_21_C249_n522, B => 
                           mult_21_C249_n1124, CI => mult_21_C249_n520, CO => 
                           mult_21_C249_n498, S => mult_21_C249_n499);
   mult_21_C249_U318 : ADFULD1 port map( A => mult_21_C249_n505, B => 
                           mult_21_C249_n518, CI => mult_21_C249_n501, CO => 
                           mult_21_C249_n496, S => mult_21_C249_n497);
   mult_21_C249_U317 : ADFULD1 port map( A => mult_21_C249_n516, B => 
                           mult_21_C249_n503, CI => mult_21_C249_n514, CO => 
                           mult_21_C249_n494, S => mult_21_C249_n495);
   mult_21_C249_U316 : ADFULD1 port map( A => mult_21_C249_n497, B => 
                           mult_21_C249_n499, CI => mult_21_C249_n512, CO => 
                           mult_21_C249_n492, S => mult_21_C249_n493);
   mult_21_C249_U315 : ADFULD1 port map( A => mult_21_C249_n510, B => 
                           mult_21_C249_n495, CI => mult_21_C249_n493, CO => 
                           mult_21_C249_n490, S => mult_21_C249_n491);
   mult_21_C249_U314 : ADHALFDL port map( A => mult_21_C249_n506, B => 
                           mult_21_C249_n1207, CO => mult_21_C249_n488, S => 
                           mult_21_C249_n489);
   mult_21_C249_U313 : ADFULD1 port map( A => mult_21_C249_n1009, B => 
                           mult_21_C249_n1077, CI => mult_21_C249_n1023, CO => 
                           mult_21_C249_n486, S => mult_21_C249_n487);
   mult_21_C249_U312 : ADFULD1 port map( A => mult_21_C249_n1177, B => 
                           mult_21_C249_n1099, CI => mult_21_C249_n1039, CO => 
                           mult_21_C249_n484, S => mult_21_C249_n485);
   mult_21_C249_U311 : ADFULD1 port map( A => mult_21_C249_n1057, B => 
                           mult_21_C249_n1149, CI => mult_21_C249_n1123, CO => 
                           mult_21_C249_n482, S => mult_21_C249_n483);
   mult_21_C249_U310 : ADFULD1 port map( A => mult_21_C249_n504, B => 
                           mult_21_C249_n489, CI => mult_21_C249_n502, CO => 
                           mult_21_C249_n480, S => mult_21_C249_n481);
   mult_21_C249_U309 : ADFULD1 port map( A => mult_21_C249_n483, B => 
                           mult_21_C249_n500, CI => mult_21_C249_n485, CO => 
                           mult_21_C249_n478, S => mult_21_C249_n479);
   mult_21_C249_U308 : ADFULD1 port map( A => mult_21_C249_n498, B => 
                           mult_21_C249_n487, CI => mult_21_C249_n496, CO => 
                           mult_21_C249_n476, S => mult_21_C249_n477);
   mult_21_C249_U307 : ADFULD1 port map( A => mult_21_C249_n479, B => 
                           mult_21_C249_n481, CI => mult_21_C249_n494, CO => 
                           mult_21_C249_n474, S => mult_21_C249_n475);
   mult_21_C249_U306 : ADFULD1 port map( A => mult_21_C249_n492, B => 
                           mult_21_C249_n477, CI => mult_21_C249_n475, CO => 
                           mult_21_C249_n472, S => mult_21_C249_n473);
   mult_21_C249_U305 : ADHALFDL port map( A => mult_21_C249_n1206, B => 
                           mult_21_C249_n944, CO => mult_21_C249_n470, S => 
                           mult_21_C249_n471);
   mult_21_C249_U304 : ADFULD1 port map( A => mult_21_C249_n1076, B => 
                           mult_21_C249_n996, CI => mult_21_C249_n1176, CO => 
                           mult_21_C249_n468, S => mult_21_C249_n469);
   mult_21_C249_U303 : ADFULD1 port map( A => mult_21_C249_n1008, B => 
                           mult_21_C249_n1038, CI => mult_21_C249_n471, CO => 
                           mult_21_C249_n466, S => mult_21_C249_n467);
   mult_21_C249_U302 : ADFULD1 port map( A => mult_21_C249_n1022, B => 
                           mult_21_C249_n1148, CI => mult_21_C249_n1056, CO => 
                           mult_21_C249_n464, S => mult_21_C249_n465);
   mult_21_C249_U301 : ADFULD1 port map( A => mult_21_C249_n1098, B => 
                           mult_21_C249_n1122, CI => mult_21_C249_n488, CO => 
                           mult_21_C249_n462, S => mult_21_C249_n463);
   mult_21_C249_U300 : ADFULD1 port map( A => mult_21_C249_n482, B => 
                           mult_21_C249_n486, CI => mult_21_C249_n484, CO => 
                           mult_21_C249_n460, S => mult_21_C249_n461);
   mult_21_C249_U299 : ADFULD1 port map( A => mult_21_C249_n465, B => 
                           mult_21_C249_n469, CI => mult_21_C249_n467, CO => 
                           mult_21_C249_n458, S => mult_21_C249_n459);
   mult_21_C249_U298 : ADFULD1 port map( A => mult_21_C249_n480, B => 
                           mult_21_C249_n463, CI => mult_21_C249_n478, CO => 
                           mult_21_C249_n456, S => mult_21_C249_n457);
   mult_21_C249_U297 : ADFULD1 port map( A => mult_21_C249_n459, B => 
                           mult_21_C249_n461, CI => mult_21_C249_n476, CO => 
                           mult_21_C249_n454, S => mult_21_C249_n455);
   mult_21_C249_U296 : ADFULD1 port map( A => mult_21_C249_n474, B => 
                           mult_21_C249_n457, CI => mult_21_C249_n455, CO => 
                           mult_21_C249_n452, S => mult_21_C249_n453);
   mult_21_C249_U295 : ADHALFDL port map( A => mult_21_C249_n470, B => 
                           mult_21_C249_n1205, CO => mult_21_C249_n450, S => 
                           mult_21_C249_n451);
   mult_21_C249_U294 : ADFULD1 port map( A => mult_21_C249_n1175, B => 
                           mult_21_C249_n1055, CI => mult_21_C249_n1147, CO => 
                           mult_21_C249_n448, S => mult_21_C249_n449);
   mult_21_C249_U293 : ADFULD1 port map( A => mult_21_C249_n1121, B => 
                           mult_21_C249_n1021, CI => mult_21_C249_n1097, CO => 
                           mult_21_C249_n446, S => mult_21_C249_n447);
   mult_21_C249_U292 : ADFULD1 port map( A => mult_21_C249_n995, B => 
                           mult_21_C249_n1075, CI => mult_21_C249_n1007, CO => 
                           mult_21_C249_n444, S => mult_21_C249_n445);
   mult_21_C249_U291 : ADFULD1 port map( A => mult_21_C249_n451, B => 
                           mult_21_C249_n1037, CI => mult_21_C249_n468, CO => 
                           mult_21_C249_n442, S => mult_21_C249_n443);
   mult_21_C249_U290 : ADFULD1 port map( A => mult_21_C249_n464, B => 
                           mult_21_C249_n466, CI => mult_21_C249_n462, CO => 
                           mult_21_C249_n440, S => mult_21_C249_n441);
   mult_21_C249_U289 : ADFULD1 port map( A => mult_21_C249_n449, B => 
                           mult_21_C249_n445, CI => mult_21_C249_n447, CO => 
                           mult_21_C249_n438, S => mult_21_C249_n439);
   mult_21_C249_U288 : ADFULD1 port map( A => mult_21_C249_n443, B => 
                           mult_21_C249_n460, CI => mult_21_C249_n458, CO => 
                           mult_21_C249_n436, S => mult_21_C249_n437);
   mult_21_C249_U287 : ADFULD1 port map( A => mult_21_C249_n439, B => 
                           mult_21_C249_n441, CI => mult_21_C249_n456, CO => 
                           mult_21_C249_n434, S => mult_21_C249_n435);
   mult_21_C249_U286 : ADFULD1 port map( A => mult_21_C249_n454, B => 
                           mult_21_C249_n437, CI => mult_21_C249_n435, CO => 
                           mult_21_C249_n432, S => mult_21_C249_n433);
   mult_21_C249_U285 : ADHALFDL port map( A => mult_21_C249_n1204, B => 
                           mult_21_C249_n943, CO => mult_21_C249_n430, S => 
                           mult_21_C249_n431);
   mult_21_C249_U284 : ADFULD1 port map( A => mult_21_C249_n1054, B => 
                           mult_21_C249_n984, CI => mult_21_C249_n994, CO => 
                           mult_21_C249_n428, S => mult_21_C249_n429);
   mult_21_C249_U283 : ADFULD1 port map( A => mult_21_C249_n1174, B => 
                           mult_21_C249_n1036, CI => mult_21_C249_n431, CO => 
                           mult_21_C249_n426, S => mult_21_C249_n427);
   mult_21_C249_U282 : ADFULD1 port map( A => mult_21_C249_n1006, B => 
                           mult_21_C249_n1146, CI => mult_21_C249_n1020, CO => 
                           mult_21_C249_n424, S => mult_21_C249_n425);
   mult_21_C249_U281 : ADFULD1 port map( A => mult_21_C249_n1074, B => 
                           mult_21_C249_n1120, CI => mult_21_C249_n1096, CO => 
                           mult_21_C249_n422, S => mult_21_C249_n423);
   mult_21_C249_U280 : ADFULD1 port map( A => mult_21_C249_n448, B => 
                           mult_21_C249_n450, CI => mult_21_C249_n446, CO => 
                           mult_21_C249_n420, S => mult_21_C249_n421);
   mult_21_C249_U279 : ADFULD1 port map( A => mult_21_C249_n429, B => 
                           mult_21_C249_n444, CI => mult_21_C249_n423, CO => 
                           mult_21_C249_n418, S => mult_21_C249_n419);
   mult_21_C249_U278 : ADFULD1 port map( A => mult_21_C249_n427, B => 
                           mult_21_C249_n425, CI => mult_21_C249_n442, CO => 
                           mult_21_C249_n416, S => mult_21_C249_n417);
   mult_21_C249_U277 : ADFULD1 port map( A => mult_21_C249_n421, B => 
                           mult_21_C249_n440, CI => mult_21_C249_n438, CO => 
                           mult_21_C249_n414, S => mult_21_C249_n415);
   mult_21_C249_U276 : ADFULD1 port map( A => mult_21_C249_n417, B => 
                           mult_21_C249_n419, CI => mult_21_C249_n436, CO => 
                           mult_21_C249_n412, S => mult_21_C249_n413);
   mult_21_C249_U275 : ADFULD1 port map( A => mult_21_C249_n434, B => 
                           mult_21_C249_n415, CI => mult_21_C249_n413, CO => 
                           mult_21_C249_n410, S => mult_21_C249_n411);
   mult_21_C249_U274 : ADHALFDL port map( A => mult_21_C249_n430, B => 
                           mult_21_C249_n1203, CO => mult_21_C249_n408, S => 
                           mult_21_C249_n409);
   mult_21_C249_U273 : ADFULD1 port map( A => mult_21_C249_n983, B => 
                           mult_21_C249_n1053, CI => mult_21_C249_n993, CO => 
                           mult_21_C249_n406, S => mult_21_C249_n407);
   mult_21_C249_U272 : ADFULD1 port map( A => mult_21_C249_n1173, B => 
                           mult_21_C249_n1035, CI => mult_21_C249_n1145, CO => 
                           mult_21_C249_n404, S => mult_21_C249_n405);
   mult_21_C249_U271 : ADFULD1 port map( A => mult_21_C249_n1005, B => 
                           mult_21_C249_n1119, CI => mult_21_C249_n1019, CO => 
                           mult_21_C249_n402, S => mult_21_C249_n403);
   mult_21_C249_U270 : ADFULD1 port map( A => mult_21_C249_n1073, B => 
                           mult_21_C249_n1095, CI => mult_21_C249_n409, CO => 
                           mult_21_C249_n400, S => mult_21_C249_n401);
   mult_21_C249_U269 : ADFULD1 port map( A => mult_21_C249_n426, B => 
                           mult_21_C249_n428, CI => mult_21_C249_n422, CO => 
                           mult_21_C249_n398, S => mult_21_C249_n399);
   mult_21_C249_U268 : ADFULD1 port map( A => mult_21_C249_n403, B => 
                           mult_21_C249_n424, CI => mult_21_C249_n405, CO => 
                           mult_21_C249_n396, S => mult_21_C249_n397);
   mult_21_C249_U267 : ADFULD1 port map( A => mult_21_C249_n401, B => 
                           mult_21_C249_n407, CI => mult_21_C249_n420, CO => 
                           mult_21_C249_n394, S => mult_21_C249_n395);
   mult_21_C249_U266 : ADFULD1 port map( A => mult_21_C249_n399, B => 
                           mult_21_C249_n418, CI => mult_21_C249_n416, CO => 
                           mult_21_C249_n392, S => mult_21_C249_n393);
   mult_21_C249_U265 : ADFULD1 port map( A => mult_21_C249_n395, B => 
                           mult_21_C249_n397, CI => mult_21_C249_n414, CO => 
                           mult_21_C249_n390, S => mult_21_C249_n391);
   mult_21_C249_U264 : ADFULD1 port map( A => mult_21_C249_n412, B => 
                           mult_21_C249_n393, CI => mult_21_C249_n391, CO => 
                           mult_21_C249_n388, S => mult_21_C249_n389);
   mult_21_C249_U263 : ADHALFDL port map( A => mult_21_C249_n1202, B => 
                           mult_21_C249_n942, CO => mult_21_C249_n386, S => 
                           mult_21_C249_n387);
   mult_21_C249_U262 : ADFULD1 port map( A => mult_21_C249_n1052, B => 
                           mult_21_C249_n974, CI => mult_21_C249_n1172, CO => 
                           mult_21_C249_n384, S => mult_21_C249_n385);
   mult_21_C249_U261 : ADFULD1 port map( A => mult_21_C249_n982, B => 
                           mult_21_C249_n1018, CI => mult_21_C249_n387, CO => 
                           mult_21_C249_n382, S => mult_21_C249_n383);
   mult_21_C249_U260 : ADFULD1 port map( A => mult_21_C249_n992, B => 
                           mult_21_C249_n1144, CI => mult_21_C249_n1118, CO => 
                           mult_21_C249_n380, S => mult_21_C249_n381);
   mult_21_C249_U259 : ADFULD1 port map( A => mult_21_C249_n1004, B => 
                           mult_21_C249_n1094, CI => mult_21_C249_n1034, CO => 
                           mult_21_C249_n378, S => mult_21_C249_n379);
   mult_21_C249_U258 : ADFULD1 port map( A => mult_21_C249_n408, B => 
                           mult_21_C249_n1072, CI => mult_21_C249_n406, CO => 
                           mult_21_C249_n376, S => mult_21_C249_n377);
   mult_21_C249_U257 : ADFULD1 port map( A => mult_21_C249_n402, B => 
                           mult_21_C249_n404, CI => mult_21_C249_n385, CO => 
                           mult_21_C249_n374, S => mult_21_C249_n375);
   mult_21_C249_U256 : ADFULD1 port map( A => mult_21_C249_n383, B => 
                           mult_21_C249_n379, CI => mult_21_C249_n381, CO => 
                           mult_21_C249_n372, S => mult_21_C249_n373);
   mult_21_C249_U255 : ADFULD1 port map( A => mult_21_C249_n398, B => 
                           mult_21_C249_n400, CI => mult_21_C249_n377, CO => 
                           mult_21_C249_n370, S => mult_21_C249_n371);
   mult_21_C249_U254 : ADFULD1 port map( A => mult_21_C249_n375, B => 
                           mult_21_C249_n396, CI => mult_21_C249_n373, CO => 
                           mult_21_C249_n368, S => mult_21_C249_n369);
   mult_21_C249_U253 : ADFULD1 port map( A => mult_21_C249_n371, B => 
                           mult_21_C249_n394, CI => mult_21_C249_n392, CO => 
                           mult_21_C249_n366, S => mult_21_C249_n367);
   mult_21_C249_U252 : ADFULD1 port map( A => mult_21_C249_n390, B => 
                           mult_21_C249_n369, CI => mult_21_C249_n367, CO => 
                           mult_21_C249_n364, S => mult_21_C249_n365);
   mult_21_C249_U251 : ADHALFDL port map( A => mult_21_C249_n386, B => 
                           mult_21_C249_n1201, CO => mult_21_C249_n362, S => 
                           mult_21_C249_n363);
   mult_21_C249_U250 : ADFULD1 port map( A => mult_21_C249_n1171, B => 
                           mult_21_C249_n1051, CI => mult_21_C249_n1143, CO => 
                           mult_21_C249_n360, S => mult_21_C249_n361);
   mult_21_C249_U249 : ADFULD1 port map( A => mult_21_C249_n973, B => 
                           mult_21_C249_n1003, CI => mult_21_C249_n981, CO => 
                           mult_21_C249_n358, S => mult_21_C249_n359);
   mult_21_C249_U248 : ADFULD1 port map( A => mult_21_C249_n991, B => 
                           mult_21_C249_n1117, CI => mult_21_C249_n1017, CO => 
                           mult_21_C249_n356, S => mult_21_C249_n357);
   mult_21_C249_U247 : ADFULD1 port map( A => mult_21_C249_n1033, B => 
                           mult_21_C249_n1093, CI => mult_21_C249_n1071, CO => 
                           mult_21_C249_n354, S => mult_21_C249_n355);
   mult_21_C249_U246 : ADFULD1 port map( A => mult_21_C249_n384, B => 
                           mult_21_C249_n363, CI => mult_21_C249_n382, CO => 
                           mult_21_C249_n352, S => mult_21_C249_n353);
   mult_21_C249_U245 : ADFULD1 port map( A => mult_21_C249_n378, B => 
                           mult_21_C249_n380, CI => mult_21_C249_n355, CO => 
                           mult_21_C249_n350, S => mult_21_C249_n351);
   mult_21_C249_U244 : ADFULD1 port map( A => mult_21_C249_n361, B => 
                           mult_21_C249_n357, CI => mult_21_C249_n359, CO => 
                           mult_21_C249_n348, S => mult_21_C249_n349);
   mult_21_C249_U243 : ADFULD1 port map( A => mult_21_C249_n374, B => 
                           mult_21_C249_n376, CI => mult_21_C249_n353, CO => 
                           mult_21_C249_n346, S => mult_21_C249_n347);
   mult_21_C249_U242 : ADFULD1 port map( A => mult_21_C249_n351, B => 
                           mult_21_C249_n372, CI => mult_21_C249_n349, CO => 
                           mult_21_C249_n344, S => mult_21_C249_n345);
   mult_21_C249_U241 : ADFULD1 port map( A => mult_21_C249_n347, B => 
                           mult_21_C249_n370, CI => mult_21_C249_n368, CO => 
                           mult_21_C249_n342, S => mult_21_C249_n343);
   mult_21_C249_U240 : ADFULD1 port map( A => mult_21_C249_n366, B => 
                           mult_21_C249_n345, CI => mult_21_C249_n343, CO => 
                           mult_21_C249_n340, S => mult_21_C249_n341);
   mult_21_C249_U239 : ADHALFDL port map( A => mult_21_C249_n1200, B => 
                           mult_21_C249_n941, CO => mult_21_C249_n338, S => 
                           mult_21_C249_n339);
   mult_21_C249_U238 : ADFULD1 port map( A => mult_21_C249_n1050, B => 
                           mult_21_C249_n966, CI => mult_21_C249_n972, CO => 
                           mult_21_C249_n336, S => mult_21_C249_n337);
   mult_21_C249_U237 : ADFULD1 port map( A => mult_21_C249_n980, B => 
                           mult_21_C249_n1032, CI => mult_21_C249_n339, CO => 
                           mult_21_C249_n334, S => mult_21_C249_n335);
   mult_21_C249_U236 : ADFULD1 port map( A => mult_21_C249_n990, B => 
                           mult_21_C249_n1170, CI => mult_21_C249_n1002, CO => 
                           mult_21_C249_n332, S => mult_21_C249_n333);
   mult_21_C249_U235 : ADFULD1 port map( A => mult_21_C249_n1016, B => 
                           mult_21_C249_n1142, CI => mult_21_C249_n1070, CO => 
                           mult_21_C249_n330, S => mult_21_C249_n331);
   mult_21_C249_U234 : ADFULD1 port map( A => mult_21_C249_n1092, B => 
                           mult_21_C249_n1116, CI => mult_21_C249_n362, CO => 
                           mult_21_C249_n328, S => mult_21_C249_n329);
   mult_21_C249_U233 : ADFULD1 port map( A => mult_21_C249_n354, B => 
                           mult_21_C249_n360, CI => mult_21_C249_n356, CO => 
                           mult_21_C249_n326, S => mult_21_C249_n327);
   mult_21_C249_U232 : ADFULD1 port map( A => mult_21_C249_n337, B => 
                           mult_21_C249_n358, CI => mult_21_C249_n331, CO => 
                           mult_21_C249_n324, S => mult_21_C249_n325);
   mult_21_C249_U231 : ADFULD1 port map( A => mult_21_C249_n333, B => 
                           mult_21_C249_n335, CI => mult_21_C249_n329, CO => 
                           mult_21_C249_n322, S => mult_21_C249_n323);
   mult_21_C249_U230 : ADFULD1 port map( A => mult_21_C249_n350, B => 
                           mult_21_C249_n352, CI => mult_21_C249_n348, CO => 
                           mult_21_C249_n320, S => mult_21_C249_n321);
   mult_21_C249_U229 : ADFULD1 port map( A => mult_21_C249_n325, B => 
                           mult_21_C249_n327, CI => mult_21_C249_n323, CO => 
                           mult_21_C249_n318, S => mult_21_C249_n319);
   mult_21_C249_U228 : ADFULD1 port map( A => mult_21_C249_n344, B => 
                           mult_21_C249_n346, CI => mult_21_C249_n321, CO => 
                           mult_21_C249_n316, S => mult_21_C249_n317);
   mult_21_C249_U227 : ADFULD1 port map( A => mult_21_C249_n342, B => 
                           mult_21_C249_n319, CI => mult_21_C249_n317, CO => 
                           mult_21_C249_n314, S => mult_21_C249_n315);
   mult_21_C249_U226 : ADHALFDL port map( A => mult_21_C249_n338, B => 
                           mult_21_C249_n1199, CO => mult_21_C249_n312, S => 
                           mult_21_C249_n313);
   mult_21_C249_U225 : ADFULD1 port map( A => mult_21_C249_n965, B => 
                           mult_21_C249_n1031, CI => mult_21_C249_n971, CO => 
                           mult_21_C249_n310, S => mult_21_C249_n311);
   mult_21_C249_U224 : ADFULD1 port map( A => mult_21_C249_n979, B => 
                           mult_21_C249_n1049, CI => mult_21_C249_n1169, CO => 
                           mult_21_C249_n308, S => mult_21_C249_n309);
   mult_21_C249_U223 : ADFULD1 port map( A => mult_21_C249_n1141, B => 
                           mult_21_C249_n1001, CI => mult_21_C249_n989, CO => 
                           mult_21_C249_n306, S => mult_21_C249_n307);
   mult_21_C249_U222 : ADFULD1 port map( A => mult_21_C249_n1015, B => 
                           mult_21_C249_n1115, CI => mult_21_C249_n1069, CO => 
                           mult_21_C249_n304, S => mult_21_C249_n305);
   mult_21_C249_U221 : ADFULD1 port map( A => mult_21_C249_n313, B => 
                           mult_21_C249_n1091, CI => mult_21_C249_n336, CO => 
                           mult_21_C249_n302, S => mult_21_C249_n303);
   mult_21_C249_U220 : ADFULD1 port map( A => mult_21_C249_n332, B => 
                           mult_21_C249_n330, CI => mult_21_C249_n334, CO => 
                           mult_21_C249_n300, S => mult_21_C249_n301);
   mult_21_C249_U219 : ADFULD1 port map( A => mult_21_C249_n305, B => 
                           mult_21_C249_n328, CI => mult_21_C249_n311, CO => 
                           mult_21_C249_n298, S => mult_21_C249_n299);
   mult_21_C249_U218 : ADFULD1 port map( A => mult_21_C249_n307, B => 
                           mult_21_C249_n309, CI => mult_21_C249_n326, CO => 
                           mult_21_C249_n296, S => mult_21_C249_n297);
   mult_21_C249_U217 : ADFULD1 port map( A => mult_21_C249_n324, B => 
                           mult_21_C249_n303, CI => mult_21_C249_n301, CO => 
                           mult_21_C249_n294, S => mult_21_C249_n295);
   mult_21_C249_U216 : ADFULD1 port map( A => mult_21_C249_n299, B => 
                           mult_21_C249_n322, CI => mult_21_C249_n320, CO => 
                           mult_21_C249_n292, S => mult_21_C249_n293);
   mult_21_C249_U215 : ADFULD1 port map( A => mult_21_C249_n318, B => 
                           mult_21_C249_n297, CI => mult_21_C249_n295, CO => 
                           mult_21_C249_n290, S => mult_21_C249_n291);
   mult_21_C249_U214 : ADFULD1 port map( A => mult_21_C249_n316, B => 
                           mult_21_C249_n293, CI => mult_21_C249_n291, CO => 
                           mult_21_C249_n288, S => mult_21_C249_n289);
   mult_21_C249_U213 : ADHALFDL port map( A => mult_21_C249_n1198, B => 
                           mult_21_C249_n940, CO => mult_21_C249_n286, S => 
                           mult_21_C249_n287);
   mult_21_C249_U212 : ADFULD1 port map( A => mult_21_C249_n1030, B => 
                           mult_21_C249_n960, CI => mult_21_C249_n1168, CO => 
                           mult_21_C249_n284, S => mult_21_C249_n285);
   mult_21_C249_U211 : ADFULD1 port map( A => mult_21_C249_n1140, B => 
                           mult_21_C249_n1000, CI => mult_21_C249_n287, CO => 
                           mult_21_C249_n282, S => mult_21_C249_n283);
   mult_21_C249_U210 : ADFULD1 port map( A => mult_21_C249_n964, B => 
                           mult_21_C249_n1114, CI => mult_21_C249_n970, CO => 
                           mult_21_C249_n280, S => mult_21_C249_n281);
   mult_21_C249_U209 : ADFULD1 port map( A => mult_21_C249_n978, B => 
                           mult_21_C249_n1090, CI => mult_21_C249_n988, CO => 
                           mult_21_C249_n278, S => mult_21_C249_n279);
   mult_21_C249_U208 : ADFULD1 port map( A => mult_21_C249_n1014, B => 
                           mult_21_C249_n1068, CI => mult_21_C249_n1048, CO => 
                           mult_21_C249_n276, S => mult_21_C249_n277);
   mult_21_C249_U207 : ADFULD1 port map( A => mult_21_C249_n304, B => 
                           mult_21_C249_n312, CI => mult_21_C249_n306, CO => 
                           mult_21_C249_n274, S => mult_21_C249_n275);
   mult_21_C249_U206 : ADFULD1 port map( A => mult_21_C249_n310, B => 
                           mult_21_C249_n308, CI => mult_21_C249_n285, CO => 
                           mult_21_C249_n272, S => mult_21_C249_n273);
   mult_21_C249_U205 : ADFULD1 port map( A => mult_21_C249_n283, B => 
                           mult_21_C249_n277, CI => mult_21_C249_n279, CO => 
                           mult_21_C249_n270, S => mult_21_C249_n271);
   mult_21_C249_U204 : ADFULD1 port map( A => mult_21_C249_n302, B => 
                           mult_21_C249_n281, CI => mult_21_C249_n300, CO => 
                           mult_21_C249_n268, S => mult_21_C249_n269);
   mult_21_C249_U203 : ADFULD1 port map( A => mult_21_C249_n275, B => 
                           mult_21_C249_n298, CI => mult_21_C249_n273, CO => 
                           mult_21_C249_n266, S => mult_21_C249_n267);
   mult_21_C249_U202 : ADFULD1 port map( A => mult_21_C249_n296, B => 
                           mult_21_C249_n271, CI => mult_21_C249_n269, CO => 
                           mult_21_C249_n264, S => mult_21_C249_n265);
   mult_21_C249_U201 : ADFULD1 port map( A => mult_21_C249_n267, B => 
                           mult_21_C249_n294, CI => mult_21_C249_n292, CO => 
                           mult_21_C249_n262, S => mult_21_C249_n263);
   mult_21_C249_U200 : ADFULD1 port map( A => mult_21_C249_n290, B => 
                           mult_21_C249_n265, CI => mult_21_C249_n263, CO => 
                           mult_21_C249_n260, S => mult_21_C249_n261);
   mult_21_C249_U199 : ADHALFDL port map( A => mult_21_C249_n286, B => 
                           mult_21_C249_n1197, CO => mult_21_C249_n258, S => 
                           mult_21_C249_n259);
   mult_21_C249_U198 : ADFULD1 port map( A => mult_21_C249_n1167, B => 
                           mult_21_C249_n1029, CI => mult_21_C249_n1139, CO => 
                           mult_21_C249_n256, S => mult_21_C249_n257);
   mult_21_C249_U197 : ADFULD1 port map( A => mult_21_C249_n1113, B => 
                           mult_21_C249_n987, CI => mult_21_C249_n1089, CO => 
                           mult_21_C249_n254, S => mult_21_C249_n255);
   mult_21_C249_U196 : ADFULD1 port map( A => mult_21_C249_n959, B => 
                           mult_21_C249_n969, CI => mult_21_C249_n963, CO => 
                           mult_21_C249_n252, S => mult_21_C249_n253);
   mult_21_C249_U195 : ADFULD1 port map( A => mult_21_C249_n977, B => 
                           mult_21_C249_n1067, CI => mult_21_C249_n999, CO => 
                           mult_21_C249_n250, S => mult_21_C249_n251);
   mult_21_C249_U194 : ADFULD1 port map( A => mult_21_C249_n1047, B => 
                           mult_21_C249_n1013, CI => mult_21_C249_n259, CO => 
                           mult_21_C249_n248, S => mult_21_C249_n249);
   mult_21_C249_U193 : ADFULD1 port map( A => mult_21_C249_n278, B => 
                           mult_21_C249_n284, CI => mult_21_C249_n282, CO => 
                           mult_21_C249_n246, S => mult_21_C249_n247);
   mult_21_C249_U192 : ADFULD1 port map( A => mult_21_C249_n280, B => 
                           mult_21_C249_n276, CI => mult_21_C249_n251, CO => 
                           mult_21_C249_n244, S => mult_21_C249_n245);
   mult_21_C249_U191 : ADFULD1 port map( A => mult_21_C249_n253, B => 
                           mult_21_C249_n255, CI => mult_21_C249_n257, CO => 
                           mult_21_C249_n242, S => mult_21_C249_n243);
   mult_21_C249_U190 : ADFULD1 port map( A => mult_21_C249_n274, B => 
                           mult_21_C249_n249, CI => mult_21_C249_n272, CO => 
                           mult_21_C249_n240, S => mult_21_C249_n241);
   mult_21_C249_U189 : ADFULD1 port map( A => mult_21_C249_n270, B => 
                           mult_21_C249_n247, CI => mult_21_C249_n245, CO => 
                           mult_21_C249_n238, S => mult_21_C249_n239);
   mult_21_C249_U188 : ADFULD1 port map( A => mult_21_C249_n268, B => 
                           mult_21_C249_n243, CI => mult_21_C249_n241, CO => 
                           mult_21_C249_n236, S => mult_21_C249_n237);
   mult_21_C249_U187 : ADFULD1 port map( A => mult_21_C249_n239, B => 
                           mult_21_C249_n266, CI => mult_21_C249_n264, CO => 
                           mult_21_C249_n234, S => mult_21_C249_n235);
   mult_21_C249_U186 : ADFULD1 port map( A => mult_21_C249_n262, B => 
                           mult_21_C249_n237, CI => mult_21_C249_n235, CO => 
                           mult_21_C249_n232, S => mult_21_C249_n233);
   mult_21_C249_U185 : ADHALFDL port map( A => mult_21_C249_n1196, B => 
                           mult_21_C249_n939, CO => mult_21_C249_n230, S => 
                           mult_21_C249_n231);
   mult_21_C249_U184 : ADFULD1 port map( A => mult_21_C249_n1028, B => 
                           mult_21_C249_n956, CI => mult_21_C249_n958, CO => 
                           mult_21_C249_n228, S => mult_21_C249_n229);
   mult_21_C249_U183 : ADFULD1 port map( A => mult_21_C249_n1166, B => 
                           mult_21_C249_n1012, CI => mult_21_C249_n231, CO => 
                           mult_21_C249_n226, S => mult_21_C249_n227);
   mult_21_C249_U182 : ADFULD1 port map( A => mult_21_C249_n962, B => 
                           mult_21_C249_n1138, CI => mult_21_C249_n968, CO => 
                           mult_21_C249_n224, S => mult_21_C249_n225);
   mult_21_C249_U181 : ADFULD1 port map( A => mult_21_C249_n986, B => 
                           mult_21_C249_n976, CI => mult_21_C249_n998, CO => 
                           mult_21_C249_n222, S => mult_21_C249_n223);
   mult_21_C249_U180 : ADFULD1 port map( A => mult_21_C249_n1046, B => 
                           mult_21_C249_n1112, CI => mult_21_C249_n1066, CO => 
                           mult_21_C249_n220, S => mult_21_C249_n221);
   mult_21_C249_U179 : ADFULD1 port map( A => mult_21_C249_n258, B => 
                           mult_21_C249_n1088, CI => mult_21_C249_n250, CO => 
                           mult_21_C249_n218, S => mult_21_C249_n219);
   mult_21_C249_U178 : ADFULD1 port map( A => mult_21_C249_n256, B => 
                           mult_21_C249_n252, CI => mult_21_C249_n254, CO => 
                           mult_21_C249_n216, S => mult_21_C249_n217);
   mult_21_C249_U177 : ADFULD1 port map( A => mult_21_C249_n221, B => 
                           mult_21_C249_n229, CI => mult_21_C249_n227, CO => 
                           mult_21_C249_n214, S => mult_21_C249_n215);
   mult_21_C249_U176 : ADFULD1 port map( A => mult_21_C249_n225, B => 
                           mult_21_C249_n223, CI => mult_21_C249_n248, CO => 
                           mult_21_C249_n212, S => mult_21_C249_n213);
   mult_21_C249_U175 : ADFULD1 port map( A => mult_21_C249_n244, B => 
                           mult_21_C249_n246, CI => mult_21_C249_n219, CO => 
                           mult_21_C249_n210, S => mult_21_C249_n211);
   mult_21_C249_U174 : ADFULD1 port map( A => mult_21_C249_n217, B => 
                           mult_21_C249_n242, CI => mult_21_C249_n215, CO => 
                           mult_21_C249_n208, S => mult_21_C249_n209);
   mult_21_C249_U173 : ADFULD1 port map( A => mult_21_C249_n240, B => 
                           mult_21_C249_n213, CI => mult_21_C249_n238, CO => 
                           mult_21_C249_n206, S => mult_21_C249_n207);
   mult_21_C249_U172 : ADFULD1 port map( A => mult_21_C249_n209, B => 
                           mult_21_C249_n211, CI => mult_21_C249_n236, CO => 
                           mult_21_C249_n204, S => mult_21_C249_n205);
   mult_21_C249_U171 : ADFULD1 port map( A => mult_21_C249_n234, B => 
                           mult_21_C249_n207, CI => mult_21_C249_n205, CO => 
                           mult_21_C249_n202, S => mult_21_C249_n203);
   mult_21_C249_U155 : ADHALFDL port map( A => mult_21_C249_n1226, B => N3042, 
                           CO => mult_21_C249_n186, S => N3361);
   mult_21_C249_U154 : ADHALFDL port map( A => mult_21_C249_n186, B => 
                           mult_21_C249_n1225, CO => mult_21_C249_n185, S => 
                           N3362);
   mult_21_C249_U153 : ADFULD1 port map( A => mult_21_C249_n651, B => 
                           mult_21_C249_n1194, CI => mult_21_C249_n185, CO => 
                           mult_21_C249_n184, S => N3363);
   mult_21_C249_U152 : ADFULD1 port map( A => mult_21_C249_n649, B => 
                           mult_21_C249_n1193, CI => mult_21_C249_n184, CO => 
                           mult_21_C249_n183, S => N3364);
   mult_21_C249_U151 : ADFULD1 port map( A => mult_21_C249_n645, B => 
                           mult_21_C249_n648, CI => mult_21_C249_n183, CO => 
                           mult_21_C249_n182, S => N3365);
   mult_21_C249_U150 : ADFULD1 port map( A => mult_21_C249_n641, B => 
                           mult_21_C249_n644, CI => mult_21_C249_n182, CO => 
                           mult_21_C249_n181, S => N3366);
   mult_21_C249_U149 : ADFULD1 port map( A => mult_21_C249_n635, B => 
                           mult_21_C249_n640, CI => mult_21_C249_n181, CO => 
                           mult_21_C249_n180, S => N3367);
   mult_21_C249_U148 : ADFULD1 port map( A => mult_21_C249_n629, B => 
                           mult_21_C249_n634, CI => mult_21_C249_n180, CO => 
                           mult_21_C249_n179, S => N3368);
   mult_21_C249_U147 : ADFULD1 port map( A => mult_21_C249_n621, B => 
                           mult_21_C249_n628, CI => mult_21_C249_n179, CO => 
                           mult_21_C249_n178, S => N3369);
   mult_21_C249_U146 : ADFULD1 port map( A => mult_21_C249_n613, B => 
                           mult_21_C249_n620, CI => mult_21_C249_n178, CO => 
                           mult_21_C249_n177, S => N3370);
   mult_21_C249_U145 : ADFULD1 port map( A => mult_21_C249_n603, B => 
                           mult_21_C249_n612, CI => mult_21_C249_n177, CO => 
                           mult_21_C249_n176, S => N3371);
   mult_21_C249_U144 : ADFULD1 port map( A => mult_21_C249_n593, B => 
                           mult_21_C249_n602, CI => mult_21_C249_n176, CO => 
                           mult_21_C249_n175, S => N3372);
   mult_21_C249_U143 : ADFULD1 port map( A => mult_21_C249_n581, B => 
                           mult_21_C249_n592, CI => mult_21_C249_n175, CO => 
                           mult_21_C249_n174, S => N3373);
   mult_21_C249_U142 : ADFULD1 port map( A => mult_21_C249_n569, B => 
                           mult_21_C249_n580, CI => mult_21_C249_n174, CO => 
                           mult_21_C249_n173, S => N3374);
   mult_21_C249_U141 : ADFULD1 port map( A => mult_21_C249_n555, B => 
                           mult_21_C249_n568, CI => mult_21_C249_n173, CO => 
                           mult_21_C249_n172, S => N3375);
   mult_21_C249_U140 : ADFULD1 port map( A => mult_21_C249_n541, B => 
                           mult_21_C249_n554, CI => mult_21_C249_n172, CO => 
                           mult_21_C249_n171, S => N3376);
   mult_21_C249_U139 : ADFULD1 port map( A => mult_21_C249_n525, B => 
                           mult_21_C249_n540, CI => mult_21_C249_n171, CO => 
                           mult_21_C249_n170, S => N3377);
   mult_21_C249_U138 : ADFULD1 port map( A => mult_21_C249_n509, B => 
                           mult_21_C249_n524, CI => mult_21_C249_n170, CO => 
                           mult_21_C249_n169, S => N3378);
   mult_21_C249_U137 : ADFULD1 port map( A => mult_21_C249_n491, B => 
                           mult_21_C249_n508, CI => mult_21_C249_n169, CO => 
                           mult_21_C249_n168, S => N3379);
   mult_21_C249_U136 : ADFULD1 port map( A => mult_21_C249_n473, B => 
                           mult_21_C249_n490, CI => mult_21_C249_n168, CO => 
                           mult_21_C249_n167, S => N3380);
   mult_21_C249_U135 : ADFULD1 port map( A => mult_21_C249_n453, B => 
                           mult_21_C249_n472, CI => mult_21_C249_n167, CO => 
                           mult_21_C249_n166, S => N3381);
   mult_21_C249_U134 : ADFULD1 port map( A => mult_21_C249_n433, B => 
                           mult_21_C249_n452, CI => mult_21_C249_n166, CO => 
                           mult_21_C249_n165, S => N3382);
   mult_21_C249_U133 : ADFULD1 port map( A => mult_21_C249_n411, B => 
                           mult_21_C249_n432, CI => mult_21_C249_n165, CO => 
                           mult_21_C249_n164, S => N3383);
   mult_21_C249_U132 : ADFULD1 port map( A => mult_21_C249_n389, B => 
                           mult_21_C249_n410, CI => mult_21_C249_n164, CO => 
                           mult_21_C249_n163, S => N3384);
   mult_21_C249_U131 : ADFULD1 port map( A => mult_21_C249_n365, B => 
                           mult_21_C249_n388, CI => mult_21_C249_n163, CO => 
                           mult_21_C249_n162, S => N3385);
   mult_21_C249_U130 : ADFULD1 port map( A => mult_21_C249_n341, B => 
                           mult_21_C249_n364, CI => mult_21_C249_n162, CO => 
                           mult_21_C249_n161, S => N3386);
   mult_21_C249_U129 : ADFULD1 port map( A => mult_21_C249_n315, B => 
                           mult_21_C249_n340, CI => mult_21_C249_n161, CO => 
                           mult_21_C249_n160, S => N3387);
   mult_21_C249_U128 : ADFULD1 port map( A => mult_21_C249_n289, B => 
                           mult_21_C249_n314, CI => mult_21_C249_n160, CO => 
                           mult_21_C249_n159, S => N3388);
   mult_21_C249_U127 : ADFULD1 port map( A => mult_21_C249_n261, B => 
                           mult_21_C249_n288, CI => mult_21_C249_n159, CO => 
                           mult_21_C249_n158, S => N3389);
   mult_21_C249_U126 : ADFULD1 port map( A => mult_21_C249_n233, B => 
                           mult_21_C249_n260, CI => mult_21_C249_n158, CO => 
                           mult_21_C249_n157, S => N3390);
   mult_21_C249_U125 : ADFULD1 port map( A => mult_21_C249_n203, B => 
                           mult_21_C249_n232, CI => mult_21_C249_n157, CO => 
                           mult_21_C249_n156, S => N3391);

end flat_filter_none_20;
