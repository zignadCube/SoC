
library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

package CONV_PACK_gp_custom is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_gp_custom;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_gp_custom.all;

architecture hier_filter_none_5 of gp_custom_DW_mult_tc_9 is

   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AO21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component MUXB2DL
      port( A0, A1, SL : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component EXOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n6, n8, n14, n22, n30, n38, n42, n45, n48, n50, n53, n56, n58, 
      n61, n63, n66, n69, n71, n73, n76, n78, n79, n81, n83, n84, n86, n88, n89
      , n91, n93, n94, n96, n98, n99, n101, n103, n104, n105, n106, n155, n156,
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n178, n179, n180, n181, 
      n182, n183, n184, n185, n187, n188, n189, n190, n194, n195, n197, n199, 
      n200, n201, n202, n204, n206, n207, n208, n209, n211, n214, n215, n216, 
      n217, n219, n221, n222, n223, n224, n225, n226, n227, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n246, n248, n249, n251, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n268, n270, n271, n273, n275, 
      n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, 
      n288, n289, n293, n294, n295, n296, n297, n301, n302, n303, n305, n310, 
      n312, n313, n314, n315, n318, n319, n322, n323, n324, n326, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, 
      n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
      n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, 
      n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, 
      n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, 
      n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, 
      n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, 
      n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, 
      n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, 
      n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, 
      n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, 
      n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, 
      n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, 
      n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, 
      n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, 
      n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, 
      n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, 
      n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, 
      n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, 
      n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, 
      n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, 
      n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, 
      n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, 
      n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, 
      n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, 
      n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, 
      n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, 
      n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, 
      n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, 
      n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, 
      n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, 
      n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, 
      n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, 
      n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, 
      n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, 
      n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, 
      n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, 
      n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, 
      n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, 
      n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, 
      n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002
      , n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, 
      n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, 
      n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, 
      n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, 
      n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
      n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
      n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, 
      n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, 
      n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
      n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, 
      n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, 
      n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, 
      n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, 
      n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, 
      n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, 
      n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, 
      n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, 
      n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, 
      n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, 
      n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, 
      n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, 
      n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, 
      n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, 
      n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, 
      n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, 
      n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, 
      n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, 
      n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, 
      n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, 
      n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, 
      n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, 
      n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, 
      n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, 
      n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, 
      n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, 
      n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, 
      n1363, n1364, n1365, n1366, n1367, n1368, n1517, n1518, n1519, n1520, 
      n1521, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, 
      n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, 
      n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, 
      n1552, n1553, n1554, n1555, n1556, n1557 : std_logic;

begin
   
   U125 : ADFULD1 port map( A => n345, B => n374, CI => n179, CO => n178, S => 
                           product(30));
   U126 : ADFULD1 port map( A => n375, B => n402, CI => n180, CO => n179, S => 
                           product(29));
   U127 : ADFULD1 port map( A => n403, B => n430, CI => n181, CO => n180, S => 
                           product(28));
   U128 : ADFULD1 port map( A => n431, B => n456, CI => n182, CO => n181, S => 
                           product(27));
   U129 : ADFULD1 port map( A => n457, B => n482, CI => n183, CO => n182, S => 
                           product(26));
   U130 : ADFULD1 port map( A => n483, B => n506, CI => n184, CO => n183, S => 
                           product(25));
   U131 : ADFULD1 port map( A => n507, B => n530, CI => n185, CO => n184, S => 
                           product(24));
   U132 : ADFULD1 port map( A => n531, B => n552, CI => n1523, CO => n185, S =>
                           product(23));
   U134 : EXOR2D1 port map( A1 => n195, A2 => n156, Z => product(22));
   U137 : OAI21D1 port map( A1 => n202, A2 => n189, B => n190, Z => n188);
   U146 : EXNOR2D1 port map( A1 => n200, A2 => n157, Z => product(21));
   U147 : AOI21D1 port map( A1 => n200, A2 => n1528, B => n197, Z => n195);
   U154 : EXNOR2D1 port map( A1 => n207, A2 => n158, Z => product(20));
   U155 : OAI21D1 port map( A1 => n214, A2 => n201, B => n202, Z => n200);
   U157 : AOI21D1 port map( A1 => n1527, A2 => n211, B => n204, Z => n202);
   U164 : EXOR2D1 port map( A1 => n214, A2 => n159, Z => product(19));
   U165 : OAI21D1 port map( A1 => n214, A2 => n208, B => n209, Z => n207);
   U174 : EXOR2D1 port map( A1 => n222, A2 => n160, Z => product(18));
   U176 : OAI21D1 port map( A1 => n233, A2 => n216, B => n217, Z => n215);
   U178 : AOI21D1 port map( A1 => n224, A2 => n1530, B => n219, Z => n217);
   U185 : EXOR2D1 port map( A1 => n227, A2 => n161, Z => product(17));
   U186 : AOI21D1 port map( A1 => n232, A2 => n223, B => n224, Z => n222);
   U188 : OAI21D1 port map( A1 => n225, A2 => n231, B => n226, Z => n224);
   U193 : EXNOR2D1 port map( A1 => n232, A2 => n162, Z => product(16));
   U194 : AOI21D1 port map( A1 => n232, A2 => n313, B => n229, Z => n227);
   U201 : EXNOR2D1 port map( A1 => n238, A2 => n163, Z => product(15));
   U203 : AOI21D1 port map( A1 => n242, A2 => n234, B => n235, Z => n233);
   U205 : OAI21D1 port map( A1 => n236, A2 => n240, B => n237, Z => n235);
   U210 : EXOR2D1 port map( A1 => n241, A2 => n164, Z => product(14));
   U211 : OAI21D1 port map( A1 => n241, A2 => n239, B => n240, Z => n238);
   U216 : EXOR2D1 port map( A1 => n249, A2 => n165, Z => product(13));
   U218 : OAI21D1 port map( A1 => n255, A2 => n243, B => n244, Z => n242);
   U220 : AOI21D1 port map( A1 => n1532, A2 => n251, B => n246, Z => n244);
   U227 : EXNOR2D1 port map( A1 => n254, A2 => n166, Z => product(12));
   U228 : AOI21D1 port map( A1 => n254, A2 => n1531, B => n251, Z => n249);
   U235 : EXNOR2D1 port map( A1 => n260, A2 => n167, Z => product(11));
   U237 : AOI21D1 port map( A1 => n256, A2 => n264, B => n257, Z => n255);
   U239 : OAI21D1 port map( A1 => n258, A2 => n262, B => n259, Z => n257);
   U244 : EXOR2D1 port map( A1 => n263, A2 => n168, Z => product(10));
   U245 : OAI21D1 port map( A1 => n263, A2 => n261, B => n262, Z => n260);
   U250 : EXOR2D1 port map( A1 => n271, A2 => n169, Z => product(9));
   U252 : OAI21D1 port map( A1 => n265, A2 => n277, B => n266, Z => n264);
   U254 : AOI21D1 port map( A1 => n1526, A2 => n273, B => n268, Z => n266);
   U261 : EXNOR2D1 port map( A1 => n276, A2 => n170, Z => product(8));
   U262 : AOI21D1 port map( A1 => n276, A2 => n1529, B => n273, Z => n271);
   U269 : EXNOR2D1 port map( A1 => n282, A2 => n171, Z => product(7));
   U271 : AOI21D1 port map( A1 => n278, A2 => n286, B => n279, Z => n277);
   U273 : OAI21D1 port map( A1 => n280, A2 => n284, B => n281, Z => n279);
   U278 : EXOR2D1 port map( A1 => n172, A2 => n285, Z => product(6));
   U279 : OAI21D1 port map( A1 => n285, A2 => n283, B => n284, Z => n282);
   U284 : EXOR2D1 port map( A1 => n173, A2 => n289, Z => product(5));
   U286 : OAI21D1 port map( A1 => n289, A2 => n287, B => n288, Z => n286);
   U291 : EXNOR2D1 port map( A1 => n174, A2 => n294, Z => product(4));
   U299 : EXOR2D1 port map( A1 => n297, A2 => n175, Z => product(3));
   U300 : OAI21D1 port map( A1 => n297, A2 => n295, B => n296, Z => n294);
   U305 : EXNOR2D1 port map( A1 => n176, A2 => n302, Z => product(2));
   U313 : EXOR2D1 port map( A1 => n303, A2 => n305, Z => product(1));
   U321 : EXOR3D1 port map( A1 => n346, A2 => n331, A3 => n330, Z => n329);
   U322 : EXOR3D1 port map( A1 => n332, A2 => n350, A3 => n348, Z => n330);
   U323 : EXOR3D1 port map( A1 => n352, A2 => n334, A3 => n333, Z => n331);
   U324 : EXOR3D1 port map( A1 => n354, A2 => n356, A3 => n335, Z => n332);
   U325 : EXOR3D1 port map( A1 => n337, A2 => n358, A3 => n336, Z => n333);
   U326 : EXOR3D1 port map( A1 => n339, A2 => n340, A3 => n360, Z => n334);
   U327 : EXOR3D1 port map( A1 => n342, A2 => n338, A3 => n341, Z => n335);
   U328 : EXOR3D1 port map( A1 => n366, A2 => n343, A3 => n362, Z => n336);
   U329 : EXOR3D1 port map( A1 => n368, A2 => n370, A3 => n364, Z => n337);
   U330 : EXOR3D1 port map( A1 => n1187, A2 => n1169, A3 => n372, Z => n338);
   U331 : EXOR3D1 port map( A1 => n1139, A2 => n1229, A3 => n1153, Z => n339);
   U332 : EXOR3D1 port map( A1 => n1103, A2 => n1117, A3 => n1109, Z => n340);
   U333 : EXOR3D1 port map( A1 => n1253, A2 => n1127, A3 => n1099, Z => n341);
   U334 : EXOR3D1 port map( A1 => n1097, A2 => n1279, A3 => n1207, Z => n342);
   U336 : ADFULD1 port map( A => n376, B => n349, CI => n347, CO => n344, S => 
                           n345);
   U337 : ADFULD1 port map( A => n351, B => n353, CI => n378, CO => n346, S => 
                           n347);
   U338 : ADFULD1 port map( A => n382, B => n355, CI => n380, CO => n348, S => 
                           n349);
   U339 : ADFULD1 port map( A => n359, B => n384, CI => n357, CO => n350, S => 
                           n351);
   U340 : ADFULD1 port map( A => n361, B => n388, CI => n386, CO => n352, S => 
                           n353);
   U341 : ADFULD1 port map( A => n365, B => n363, CI => n390, CO => n354, S => 
                           n355);
   U342 : ADFULD1 port map( A => n369, B => n371, CI => n367, CO => n356, S => 
                           n357);
   U343 : ADFULD1 port map( A => n398, B => n394, CI => n396, CO => n358, S => 
                           n359);
   U344 : ADFULD1 port map( A => n373, B => n400, CI => n392, CO => n360, S => 
                           n361);
   U345 : ADFULD1 port map( A => n1170, B => n1118, CI => n1140, CO => n362, S 
                           => n363);
   U346 : ADFULD1 port map( A => n1104, B => n1188, CI => n1110, CO => n364, S 
                           => n365);
   U347 : ADFULD1 port map( A => n1254, B => n1128, CI => n1230, CO => n366, S 
                           => n367);
   U348 : ADFULD1 port map( A => n1280, B => n1154, CI => n1208, CO => n368, S 
                           => n369);
   U349 : ADFULD1 port map( A => n1100, B => n1338, CI => n1308, CO => n370, S 
                           => n371);
   U351 : ADFULD1 port map( A => n404, B => n379, CI => n377, CO => n374, S => 
                           n375);
   U352 : ADFULD1 port map( A => n381, B => n408, CI => n406, CO => n376, S => 
                           n377);
   U353 : ADFULD1 port map( A => n410, B => n385, CI => n383, CO => n378, S => 
                           n379);
   U354 : ADFULD1 port map( A => n412, B => n389, CI => n387, CO => n380, S => 
                           n381);
   U355 : ADFULD1 port map( A => n391, B => n416, CI => n414, CO => n382, S => 
                           n383);
   U356 : ADFULD1 port map( A => n395, B => n397, CI => n399, CO => n384, S => 
                           n385);
   U357 : ADFULD1 port map( A => n418, B => n422, CI => n393, CO => n386, S => 
                           n387);
   U358 : ADFULD1 port map( A => n424, B => n426, CI => n420, CO => n388, S => 
                           n389);
   U359 : ADFULD1 port map( A => n428, B => n1189, CI => n401, CO => n390, S =>
                           n391);
   U360 : ADFULD1 port map( A => n1141, B => n1231, CI => n1171, CO => n392, S 
                           => n393);
   U361 : ADFULD1 port map( A => n1255, B => n1119, CI => n1111, CO => n394, S 
                           => n395);
   U362 : ADFULD1 port map( A => n1281, B => n1129, CI => n1105, CO => n396, S 
                           => n397);
   U363 : ADFULD1 port map( A => n1101, B => n1155, CI => n1209, CO => n398, S 
                           => n399);
   U365 : ADFULD1 port map( A => n432, B => n407, CI => n405, CO => n402, S => 
                           n403);
   U366 : ADFULD1 port map( A => n409, B => n436, CI => n434, CO => n404, S => 
                           n405);
   U367 : ADFULD1 port map( A => n438, B => n413, CI => n411, CO => n406, S => 
                           n407);
   U368 : ADFULD1 port map( A => n440, B => n417, CI => n415, CO => n408, S => 
                           n409);
   U369 : ADFULD1 port map( A => n444, B => n419, CI => n442, CO => n410, S => 
                           n411);
   U370 : ADFULD1 port map( A => n421, B => n423, CI => n425, CO => n412, S => 
                           n413);
   U371 : ADFULD1 port map( A => n448, B => n446, CI => n427, CO => n414, S => 
                           n415);
   U372 : ADFULD1 port map( A => n452, B => n429, CI => n450, CO => n416, S => 
                           n417);
   U373 : ADFULD1 port map( A => n1232, B => n1190, CI => n454, CO => n418, S 
                           => n419);
   U374 : ADFULD1 port map( A => n1142, B => n1256, CI => n1172, CO => n420, S 
                           => n421);
   U375 : ADFULD1 port map( A => n1112, B => n1130, CI => n1120, CO => n422, S 
                           => n423);
   U376 : ADFULD1 port map( A => n1282, B => n1156, CI => n1210, CO => n424, S 
                           => n425);
   U377 : ADFULD1 port map( A => n1106, B => n1340, CI => n1310, CO => n426, S 
                           => n427);
   U379 : ADFULD1 port map( A => n458, B => n435, CI => n433, CO => n430, S => 
                           n431);
   U380 : ADFULD1 port map( A => n437, B => n439, CI => n460, CO => n432, S => 
                           n433);
   U381 : ADFULD1 port map( A => n441, B => n464, CI => n462, CO => n434, S => 
                           n435);
   U382 : ADFULD1 port map( A => n466, B => n445, CI => n443, CO => n436, S => 
                           n437);
   U383 : ADFULD1 port map( A => n449, B => n451, CI => n468, CO => n438, S => 
                           n439);
   U384 : ADFULD1 port map( A => n453, B => n447, CI => n470, CO => n440, S => 
                           n441);
   U385 : ADFULD1 port map( A => n474, B => n472, CI => n476, CO => n442, S => 
                           n443);
   U386 : ADFULD1 port map( A => n455, B => n480, CI => n478, CO => n444, S => 
                           n445);
   U387 : ADFULD1 port map( A => n1131, B => n1191, CI => n1173, CO => n446, S 
                           => n447);
   U388 : ADFULD1 port map( A => n1113, B => n1233, CI => n1121, CO => n448, S 
                           => n449);
   U389 : ADFULD1 port map( A => n1283, B => n1143, CI => n1257, CO => n450, S 
                           => n451);
   U390 : ADFULD1 port map( A => n1107, B => n1157, CI => n1211, CO => n452, S 
                           => n453);
   U392 : ADFULD1 port map( A => n484, B => n461, CI => n459, CO => n456, S => 
                           n457);
   U393 : ADFULD1 port map( A => n486, B => n488, CI => n463, CO => n458, S => 
                           n459);
   U394 : ADFULD1 port map( A => n467, B => n469, CI => n465, CO => n460, S => 
                           n461);
   U395 : ADFULD1 port map( A => n492, B => n494, CI => n490, CO => n462, S => 
                           n463);
   U396 : ADFULD1 port map( A => n475, B => n477, CI => n471, CO => n464, S => 
                           n465);
   U397 : ADFULD1 port map( A => n479, B => n500, CI => n473, CO => n466, S => 
                           n467);
   U398 : ADFULD1 port map( A => n498, B => n502, CI => n496, CO => n468, S => 
                           n469);
   U399 : ADFULD1 port map( A => n504, B => n1192, CI => n481, CO => n470, S =>
                           n471);
   U400 : ADFULD1 port map( A => n1144, B => n1234, CI => n1158, CO => n472, S 
                           => n473);
   U401 : ADFULD1 port map( A => n1258, B => n1132, CI => n1122, CO => n474, S 
                           => n475);
   U402 : ADFULD1 port map( A => n1284, B => n1174, CI => n1212, CO => n476, S 
                           => n477);
   U403 : ADFULD1 port map( A => n1114, B => n1342, CI => n1312, CO => n478, S 
                           => n479);
   U405 : ADFULD1 port map( A => n508, B => n487, CI => n485, CO => n482, S => 
                           n483);
   U406 : ADFULD1 port map( A => n510, B => n512, CI => n489, CO => n484, S => 
                           n485);
   U407 : ADFULD1 port map( A => n493, B => n514, CI => n491, CO => n486, S => 
                           n487);
   U408 : ADFULD1 port map( A => n516, B => n518, CI => n495, CO => n488, S => 
                           n489);
   U409 : ADFULD1 port map( A => n501, B => n503, CI => n497, CO => n490, S => 
                           n491);
   U410 : ADFULD1 port map( A => n522, B => n524, CI => n499, CO => n492, S => 
                           n493);
   U411 : ADFULD1 port map( A => n526, B => n505, CI => n520, CO => n494, S => 
                           n495);
   U412 : ADFULD1 port map( A => n1235, B => n1259, CI => n528, CO => n496, S 
                           => n497);
   U413 : ADFULD1 port map( A => n1159, B => n1285, CI => n1193, CO => n498, S 
                           => n499);
   U414 : ADFULD1 port map( A => n1123, B => n1145, CI => n1133, CO => n500, S 
                           => n501);
   U415 : ADFULD1 port map( A => n1115, B => n1175, CI => n1213, CO => n502, S 
                           => n503);
   U417 : ADFULD1 port map( A => n532, B => n511, CI => n509, CO => n506, S => 
                           n507);
   U418 : ADFULD1 port map( A => n513, B => n536, CI => n534, CO => n508, S => 
                           n509);
   U419 : ADFULD1 port map( A => n517, B => n538, CI => n515, CO => n510, S => 
                           n511);
   U420 : ADFULD1 port map( A => n540, B => n542, CI => n519, CO => n512, S => 
                           n513);
   U421 : ADFULD1 port map( A => n525, B => n521, CI => n523, CO => n514, S => 
                           n515);
   U422 : ADFULD1 port map( A => n544, B => n546, CI => n527, CO => n516, S => 
                           n517);
   U423 : ADFULD1 port map( A => n529, B => n550, CI => n548, CO => n518, S => 
                           n519);
   U424 : ADFULD1 port map( A => n1194, B => n1260, CI => n1236, CO => n520, S 
                           => n521);
   U425 : ADFULD1 port map( A => n1134, B => n1286, CI => n1160, CO => n522, S 
                           => n523);
   U426 : ADFULD1 port map( A => n1124, B => n1176, CI => n1214, CO => n524, S 
                           => n525);
   U427 : ADFULD1 port map( A => n1146, B => n1344, CI => n1314, CO => n526, S 
                           => n527);
   U429 : ADFULD1 port map( A => n554, B => n535, CI => n533, CO => n530, S => 
                           n531);
   U430 : ADFULD1 port map( A => n556, B => n539, CI => n537, CO => n532, S => 
                           n533);
   U431 : ADFULD1 port map( A => n541, B => n560, CI => n558, CO => n534, S => 
                           n535);
   U432 : ADFULD1 port map( A => n562, B => n545, CI => n543, CO => n536, S => 
                           n537);
   U433 : ADFULD1 port map( A => n549, B => n564, CI => n547, CO => n538, S => 
                           n539);
   U434 : ADFULD1 port map( A => n566, B => n570, CI => n568, CO => n540, S => 
                           n541);
   U435 : ADFULD1 port map( A => n572, B => n1195, CI => n551, CO => n542, S =>
                           n543);
   U436 : ADFULD1 port map( A => n1135, B => n1237, CI => n1147, CO => n544, S 
                           => n545);
   U437 : ADFULD1 port map( A => n1287, B => n1161, CI => n1261, CO => n546, S 
                           => n547);
   U438 : ADFULD1 port map( A => n1125, B => n1177, CI => n1215, CO => n548, S 
                           => n549);
   U440 : ADFULD1 port map( A => n576, B => n557, CI => n555, CO => n552, S => 
                           n553);
   U441 : ADFULD1 port map( A => n559, B => n561, CI => n578, CO => n554, S => 
                           n555);
   U442 : ADFULD1 port map( A => n563, B => n582, CI => n580, CO => n556, S => 
                           n557);
   U443 : ADFULD1 port map( A => n565, B => n569, CI => n584, CO => n558, S => 
                           n559);
   U444 : ADFULD1 port map( A => n571, B => n586, CI => n567, CO => n560, S => 
                           n561);
   U445 : ADFULD1 port map( A => n590, B => n573, CI => n588, CO => n562, S => 
                           n563);
   U446 : ADFULD1 port map( A => n1196, B => n1238, CI => n592, CO => n564, S 
                           => n565);
   U447 : ADFULD1 port map( A => n1148, B => n1262, CI => n1162, CO => n566, S 
                           => n567);
   U448 : ADFULD1 port map( A => n1288, B => n1178, CI => n1216, CO => n568, S 
                           => n569);
   U449 : ADFULD1 port map( A => n1136, B => n1346, CI => n1316, CO => n570, S 
                           => n571);
   U451 : ADFULD1 port map( A => n596, B => n579, CI => n577, CO => n574, S => 
                           n575);
   U452 : ADFULD1 port map( A => n581, B => n583, CI => n598, CO => n576, S => 
                           n577);
   U453 : ADFULD1 port map( A => n585, B => n602, CI => n600, CO => n578, S => 
                           n579);
   U454 : ADFULD1 port map( A => n591, B => n589, CI => n604, CO => n580, S => 
                           n581);
   U455 : ADFULD1 port map( A => n606, B => n608, CI => n587, CO => n582, S => 
                           n583);
   U456 : ADFULD1 port map( A => n593, B => n612, CI => n610, CO => n584, S => 
                           n585);
   U457 : ADFULD1 port map( A => n1197, B => n1263, CI => n1239, CO => n586, S 
                           => n587);
   U458 : ADFULD1 port map( A => n1289, B => n1163, CI => n1149, CO => n588, S 
                           => n589);
   U459 : ADFULD1 port map( A => n1137, B => n1179, CI => n1217, CO => n590, S 
                           => n591);
   U461 : ADFULD1 port map( A => n616, B => n599, CI => n597, CO => n594, S => 
                           n595);
   U462 : ADFULD1 port map( A => n601, B => n603, CI => n618, CO => n596, S => 
                           n597);
   U463 : ADFULD1 port map( A => n622, B => n605, CI => n620, CO => n598, S => 
                           n599);
   U464 : ADFULD1 port map( A => n609, B => n611, CI => n607, CO => n600, S => 
                           n601);
   U465 : ADFULD1 port map( A => n626, B => n628, CI => n624, CO => n602, S => 
                           n603);
   U466 : ADFULD1 port map( A => n630, B => n1240, CI => n613, CO => n604, S =>
                           n605);
   U467 : ADFULD1 port map( A => n1150, B => n1264, CI => n1180, CO => n606, S 
                           => n607);
   U468 : ADFULD1 port map( A => n1290, B => n1198, CI => n1218, CO => n608, S 
                           => n609);
   U469 : ADFULD1 port map( A => n1164, B => n1348, CI => n1318, CO => n610, S 
                           => n611);
   U471 : ADFULD1 port map( A => n634, B => n619, CI => n617, CO => n614, S => 
                           n615);
   U472 : ADFULD1 port map( A => n621, B => n623, CI => n636, CO => n616, S => 
                           n617);
   U473 : ADFULD1 port map( A => n640, B => n625, CI => n638, CO => n618, S => 
                           n619);
   U474 : ADFULD1 port map( A => n627, B => n644, CI => n629, CO => n620, S => 
                           n621);
   U475 : ADFULD1 port map( A => n646, B => n631, CI => n642, CO => n622, S => 
                           n623);
   U476 : ADFULD1 port map( A => n1241, B => n1265, CI => n648, CO => n624, S 
                           => n625);
   U477 : ADFULD1 port map( A => n1291, B => n1181, CI => n1165, CO => n626, S 
                           => n627);
   U478 : ADFULD1 port map( A => n1151, B => n1199, CI => n1219, CO => n628, S 
                           => n629);
   U480 : ADFULD1 port map( A => n652, B => n637, CI => n635, CO => n632, S => 
                           n633);
   U481 : ADFULD1 port map( A => n639, B => n641, CI => n654, CO => n634, S => 
                           n635);
   U482 : ADFULD1 port map( A => n658, B => n645, CI => n656, CO => n636, S => 
                           n637);
   U483 : ADFULD1 port map( A => n647, B => n660, CI => n643, CO => n638, S => 
                           n639);
   U484 : ADFULD1 port map( A => n649, B => n664, CI => n662, CO => n640, S => 
                           n641);
   U485 : ADFULD1 port map( A => n1182, B => n1292, CI => n1242, CO => n642, S 
                           => n643);
   U486 : ADFULD1 port map( A => n1166, B => n1266, CI => n1220, CO => n644, S 
                           => n645);
   U487 : ADFULD1 port map( A => n1200, B => n1350, CI => n1320, CO => n646, S 
                           => n647);
   U489 : ADFULD1 port map( A => n668, B => n655, CI => n653, CO => n650, S => 
                           n651);
   U490 : ADFULD1 port map( A => n670, B => n659, CI => n657, CO => n652, S => 
                           n653);
   U491 : ADFULD1 port map( A => n663, B => n661, CI => n672, CO => n654, S => 
                           n655);
   U492 : ADFULD1 port map( A => n676, B => n678, CI => n674, CO => n656, S => 
                           n657);
   U493 : ADFULD1 port map( A => n680, B => n1293, CI => n665, CO => n658, S =>
                           n659);
   U494 : ADFULD1 port map( A => n1243, B => n1183, CI => n1267, CO => n660, S 
                           => n661);
   U495 : ADFULD1 port map( A => n1167, B => n1201, CI => n1221, CO => n662, S 
                           => n663);
   U497 : ADFULD1 port map( A => n684, B => n671, CI => n669, CO => n666, S => 
                           n667);
   U498 : ADFULD1 port map( A => n686, B => n688, CI => n673, CO => n668, S => 
                           n669);
   U499 : ADFULD1 port map( A => n677, B => n679, CI => n675, CO => n670, S => 
                           n671);
   U500 : ADFULD1 port map( A => n692, B => n681, CI => n690, CO => n672, S => 
                           n673);
   U501 : ADFULD1 port map( A => n1244, B => n1294, CI => n694, CO => n674, S 
                           => n675);
   U502 : ADFULD1 port map( A => n1184, B => n1268, CI => n1222, CO => n676, S 
                           => n677);
   U503 : ADFULD1 port map( A => n1202, B => n1352, CI => n1322, CO => n678, S 
                           => n679);
   U505 : ADFULD1 port map( A => n698, B => n687, CI => n685, CO => n682, S => 
                           n683);
   U506 : ADFULD1 port map( A => n700, B => n702, CI => n689, CO => n684, S => 
                           n685);
   U507 : ADFULD1 port map( A => n691, B => n704, CI => n693, CO => n686, S => 
                           n687);
   U508 : ADFULD1 port map( A => n695, B => n708, CI => n706, CO => n688, S => 
                           n689);
   U509 : ADFULD1 port map( A => n1203, B => n1295, CI => n1245, CO => n690, S 
                           => n691);
   U510 : ADFULD1 port map( A => n1185, B => n1269, CI => n1223, CO => n692, S 
                           => n693);
   U512 : ADFULD1 port map( A => n712, B => n701, CI => n699, CO => n696, S => 
                           n697);
   U513 : ADFULD1 port map( A => n703, B => n705, CI => n714, CO => n698, S => 
                           n699);
   U514 : ADFULD1 port map( A => n716, B => n718, CI => n707, CO => n700, S => 
                           n701);
   U515 : ADFULD1 port map( A => n720, B => n1270, CI => n709, CO => n702, S =>
                           n703);
   U516 : ADFULD1 port map( A => n1246, B => n1296, CI => n1224, CO => n704, S 
                           => n705);
   U517 : ADFULD1 port map( A => n1204, B => n1354, CI => n1324, CO => n706, S 
                           => n707);
   U519 : ADFULD1 port map( A => n724, B => n715, CI => n713, CO => n710, S => 
                           n711);
   U520 : ADFULD1 port map( A => n717, B => n719, CI => n726, CO => n712, S => 
                           n713);
   U521 : ADFULD1 port map( A => n730, B => n721, CI => n728, CO => n714, S => 
                           n715);
   U522 : ADFULD1 port map( A => n1247, B => n1271, CI => n732, CO => n716, S 
                           => n717);
   U523 : ADFULD1 port map( A => n1205, B => n1297, CI => n1225, CO => n718, S 
                           => n719);
   U525 : ADFULD1 port map( A => n736, B => n727, CI => n725, CO => n722, S => 
                           n723);
   U526 : ADFULD1 port map( A => n729, B => n731, CI => n738, CO => n724, S => 
                           n725);
   U527 : ADFULD1 port map( A => n733, B => n742, CI => n740, CO => n726, S => 
                           n727);
   U528 : ADFULD1 port map( A => n1272, B => n1298, CI => n1226, CO => n728, S 
                           => n729);
   U529 : ADFULD1 port map( A => n1248, B => n1356, CI => n1326, CO => n730, S 
                           => n731);
   U531 : ADFULD1 port map( A => n746, B => n739, CI => n737, CO => n734, S => 
                           n735);
   U532 : ADFULD1 port map( A => n748, B => n750, CI => n741, CO => n736, S => 
                           n737);
   U533 : ADFULD1 port map( A => n752, B => n1299, CI => n743, CO => n738, S =>
                           n739);
   U534 : ADFULD1 port map( A => n1273, B => n1249, CI => n1227, CO => n740, S 
                           => n741);
   U536 : ADFULD1 port map( A => n756, B => n749, CI => n747, CO => n744, S => 
                           n745);
   U537 : ADFULD1 port map( A => n758, B => n753, CI => n751, CO => n746, S => 
                           n747);
   U538 : ADFULD1 port map( A => n1274, B => n1300, CI => n760, CO => n748, S 
                           => n749);
   U539 : ADFULD1 port map( A => n1250, B => n1358, CI => n1328, CO => n750, S 
                           => n751);
   U541 : ADFULD1 port map( A => n764, B => n759, CI => n757, CO => n754, S => 
                           n755);
   U542 : ADFULD1 port map( A => n761, B => n768, CI => n766, CO => n756, S => 
                           n757);
   U543 : ADFULD1 port map( A => n1275, B => n1301, CI => n1251, CO => n758, S 
                           => n759);
   U545 : ADFULD1 port map( A => n767, B => n772, CI => n765, CO => n762, S => 
                           n763);
   U546 : ADFULD1 port map( A => n774, B => n1302, CI => n769, CO => n764, S =>
                           n765);
   U547 : ADFULD1 port map( A => n1276, B => n1360, CI => n1330, CO => n766, S 
                           => n767);
   U549 : ADFULD1 port map( A => n778, B => n775, CI => n773, CO => n770, S => 
                           n771);
   U550 : ADFULD1 port map( A => n1277, B => n1303, CI => n780, CO => n772, S 
                           => n773);
   U552 : ADFULD1 port map( A => n781, B => n784, CI => n779, CO => n776, S => 
                           n777);
   U553 : ADFULD1 port map( A => n1304, B => n1362, CI => n1332, CO => n778, S 
                           => n779);
   U555 : ADFULD1 port map( A => n788, B => n1305, CI => n785, CO => n782, S =>
                           n783);
   U557 : ADFULD1 port map( A => n1334, B => n1364, CI => n790, CO => n786, S 
                           => n787);
   U561 : NOR2M1D1 port map( A1 => n104, A2 => n105, Z => n1081);
   U562 : MUXB2DL port map( A0 => n104, A1 => n105, SL => n794, Z => n1097);
   U563 : MUXB2DL port map( A0 => n1553, A1 => b(0), SL => n106, Z => n794);
   U564 : MUXB2DL port map( A0 => n104, A1 => n105, SL => n795, Z => n1098);
   U565 : NAN2M1D1 port map( A1 => n106, A2 => n1556, Z => n795);
   U566 : NOR2M1D1 port map( A1 => n99, A2 => n101, Z => n1082);
   U567 : MUXB2DL port map( A0 => n99, A1 => n101, SL => n796, Z => n1099);
   U568 : MUXB2DL port map( A0 => n1551, A1 => b(2), SL => n103, Z => n796);
   U569 : MUXB2DL port map( A0 => n99, A1 => n101, SL => n797, Z => n1100);
   U570 : MUXB2DL port map( A0 => b(2), A1 => n1553, SL => n103, Z => n797);
   U571 : MUXB2DL port map( A0 => n99, A1 => n101, SL => n798, Z => n1101);
   U572 : MUXB2DL port map( A0 => n1553, A1 => b(0), SL => n103, Z => n798);
   U573 : MUXB2DL port map( A0 => n99, A1 => n101, SL => n799, Z => n1102);
   U574 : NAN2M1D1 port map( A1 => n103, A2 => n1556, Z => n799);
   U575 : NOR2M1D1 port map( A1 => n94, A2 => n96, Z => n1083);
   U576 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n800, Z => n1103);
   U577 : MUXB2DL port map( A0 => b(5), A1 => n1549, SL => n98, Z => n800);
   U578 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n801, Z => n1104);
   U579 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n98, Z => n801);
   U580 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n802, Z => n1105);
   U581 : MUXB2DL port map( A0 => n1551, A1 => b(2), SL => n98, Z => n802);
   U582 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n803, Z => n1106);
   U583 : MUXB2DL port map( A0 => b(2), A1 => n1554, SL => n98, Z => n803);
   U584 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n804, Z => n1107);
   U585 : MUXB2DL port map( A0 => n1553, A1 => b(0), SL => n98, Z => n804);
   U586 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n805, Z => n1108);
   U587 : NAN2M1D1 port map( A1 => n98, A2 => n1556, Z => n805);
   U588 : NOR2M1D1 port map( A1 => n89, A2 => n91, Z => n1084);
   U589 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n806, Z => n1109);
   U590 : MUXB2DL port map( A0 => b(7), A1 => n1545, SL => n93, Z => n806);
   U591 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n807, Z => n1110);
   U592 : MUXB2DL port map( A0 => b(6), A1 => n1547, SL => n93, Z => n807);
   U593 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n808, Z => n1111);
   U594 : MUXB2DL port map( A0 => b(5), A1 => n1549, SL => n93, Z => n808);
   U595 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n809, Z => n1112);
   U596 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n93, Z => n809);
   U597 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n810, Z => n1113);
   U598 : MUXB2DL port map( A0 => n1551, A1 => b(2), SL => n93, Z => n810);
   U599 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n811, Z => n1114);
   U600 : MUXB2DL port map( A0 => b(2), A1 => n1553, SL => n93, Z => n811);
   U601 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n812, Z => n1115);
   U602 : MUXB2DL port map( A0 => n1553, A1 => b(0), SL => n93, Z => n812);
   U603 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n813, Z => n1116);
   U604 : NAN2M1D1 port map( A1 => n93, A2 => b(0), Z => n813);
   U605 : NOR2M1D1 port map( A1 => n84, A2 => n86, Z => n1085);
   U606 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n814, Z => n1117);
   U607 : MUXB2DL port map( A0 => n1541, A1 => b(8), SL => n88, Z => n814);
   U608 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n815, Z => n1118);
   U609 : MUXB2DL port map( A0 => b(8), A1 => n1543, SL => n88, Z => n815);
   U610 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n816, Z => n1119);
   U611 : MUXB2DL port map( A0 => b(7), A1 => n1545, SL => n88, Z => n816);
   U612 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n817, Z => n1120);
   U613 : MUXB2DL port map( A0 => b(6), A1 => n1547, SL => n88, Z => n817);
   U614 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n818, Z => n1121);
   U615 : MUXB2DL port map( A0 => b(5), A1 => n1549, SL => n88, Z => n818);
   U616 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n819, Z => n1122);
   U617 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n88, Z => n819);
   U618 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n820, Z => n1123);
   U619 : MUXB2DL port map( A0 => n1551, A1 => b(2), SL => n88, Z => n820);
   U620 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n821, Z => n1124);
   U621 : MUXB2DL port map( A0 => b(2), A1 => n1554, SL => n88, Z => n821);
   U622 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n822, Z => n1125);
   U623 : MUXB2DL port map( A0 => n1553, A1 => b(0), SL => n88, Z => n822);
   U624 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n823, Z => n1126);
   U625 : NAN2M1D1 port map( A1 => n88, A2 => b(0), Z => n823);
   U626 : NOR2M1D1 port map( A1 => n79, A2 => n81, Z => n1086);
   U627 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n824, Z => n1127);
   U628 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n83, Z => n824);
   U629 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n825, Z => n1128);
   U630 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n83, Z => n825);
   U631 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n826, Z => n1129);
   U632 : MUXB2DL port map( A0 => n1541, A1 => b(8), SL => n83, Z => n826);
   U633 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n827, Z => n1130);
   U634 : MUXB2DL port map( A0 => b(8), A1 => n1543, SL => n83, Z => n827);
   U635 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n828, Z => n1131);
   U636 : MUXB2DL port map( A0 => b(7), A1 => n1545, SL => n83, Z => n828);
   U637 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n829, Z => n1132);
   U638 : MUXB2DL port map( A0 => b(6), A1 => n1547, SL => n83, Z => n829);
   U639 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n830, Z => n1133);
   U640 : MUXB2DL port map( A0 => b(5), A1 => n1549, SL => n83, Z => n830);
   U641 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n831, Z => n1134);
   U642 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n83, Z => n831);
   U643 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n832, Z => n1135);
   U644 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n83, Z => n832);
   U645 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n833, Z => n1136);
   U646 : MUXB2DL port map( A0 => b(2), A1 => n1554, SL => n83, Z => n833);
   U647 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n834, Z => n1137);
   U648 : MUXB2DL port map( A0 => n1553, A1 => b(0), SL => n83, Z => n834);
   U649 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n835, Z => n1138);
   U650 : NAN2M1D1 port map( A1 => n83, A2 => n1556, Z => n835);
   U651 : NOR2M1D1 port map( A1 => n73, A2 => n76, Z => n1087);
   U652 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n836, Z => n1139);
   U653 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n78, Z => n836);
   U654 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n837, Z => n1140);
   U655 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n78, Z => n837);
   U656 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n838, Z => n1141);
   U657 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n78, Z => n838);
   U658 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n839, Z => n1142);
   U659 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n78, Z => n839);
   U660 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n840, Z => n1143);
   U661 : MUXB2DL port map( A0 => n1541, A1 => b(8), SL => n78, Z => n840);
   U662 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n841, Z => n1144);
   U663 : MUXB2DL port map( A0 => b(8), A1 => n1543, SL => n78, Z => n841);
   U664 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n842, Z => n1145);
   U665 : MUXB2DL port map( A0 => b(7), A1 => n1545, SL => n78, Z => n842);
   U666 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n843, Z => n1146);
   U667 : MUXB2DL port map( A0 => b(6), A1 => n1547, SL => n78, Z => n843);
   U668 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n844, Z => n1147);
   U669 : MUXB2DL port map( A0 => b(5), A1 => n1549, SL => n78, Z => n844);
   U670 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n845, Z => n1148);
   U671 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n78, Z => n845);
   U672 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n846, Z => n1149);
   U673 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n78, Z => n846);
   U674 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n847, Z => n1150);
   U675 : MUXB2DL port map( A0 => b(2), A1 => n1554, SL => n78, Z => n847);
   U676 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n848, Z => n1151);
   U677 : MUXB2DL port map( A0 => n1553, A1 => n1556, SL => n78, Z => n848);
   U678 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n849, Z => n1152);
   U679 : NAN2M1D1 port map( A1 => n78, A2 => b(0), Z => n849);
   U680 : NOR2M1D1 port map( A1 => n66, A2 => n69, Z => n1088);
   U681 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n850, Z => n1153);
   U682 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n71, Z => n850);
   U683 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n851, Z => n1154);
   U684 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n71, Z => n851);
   U685 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n852, Z => n1155);
   U686 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n71, Z => n852);
   U687 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n853, Z => n1156);
   U688 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n71, Z => n853);
   U689 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n854, Z => n1157);
   U690 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n71, Z => n854);
   U691 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n855, Z => n1158);
   U692 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n71, Z => n855);
   U693 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n856, Z => n1159);
   U694 : MUXB2DL port map( A0 => n1541, A1 => b(8), SL => n71, Z => n856);
   U695 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n857, Z => n1160);
   U696 : MUXB2DL port map( A0 => b(8), A1 => n1543, SL => n71, Z => n857);
   U697 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n858, Z => n1161);
   U698 : MUXB2DL port map( A0 => b(7), A1 => n1545, SL => n71, Z => n858);
   U699 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n859, Z => n1162);
   U700 : MUXB2DL port map( A0 => b(6), A1 => n1547, SL => n71, Z => n859);
   U701 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n860, Z => n1163);
   U702 : MUXB2DL port map( A0 => n1547, A1 => n1549, SL => n71, Z => n860);
   U703 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n861, Z => n1164);
   U704 : MUXB2DL port map( A0 => n1549, A1 => n1551, SL => n71, Z => n861);
   U705 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n862, Z => n1165);
   U706 : MUXB2DL port map( A0 => n1551, A1 => b(2), SL => n71, Z => n862);
   U707 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n863, Z => n1166);
   U708 : MUXB2DL port map( A0 => b(2), A1 => n1554, SL => n71, Z => n863);
   U709 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n864, Z => n1167);
   U710 : MUXB2DL port map( A0 => n1553, A1 => b(0), SL => n71, Z => n864);
   U711 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n865, Z => n1168);
   U712 : NAN2M1D1 port map( A1 => n71, A2 => n1556, Z => n865);
   U713 : NOR2M1D1 port map( A1 => n58, A2 => n61, Z => n1089);
   U714 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n866, Z => n1169);
   U715 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n63, Z => n866);
   U716 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n867, Z => n1170);
   U717 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n63, Z => n867);
   U718 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n868, Z => n1171);
   U719 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n63, Z => n868);
   U720 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n869, Z => n1172);
   U721 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n63, Z => n869);
   U722 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n870, Z => n1173);
   U723 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n63, Z => n870);
   U724 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n871, Z => n1174);
   U725 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n63, Z => n871);
   U726 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n872, Z => n1175);
   U727 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n63, Z => n872);
   U728 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n873, Z => n1176);
   U729 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n63, Z => n873);
   U730 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n874, Z => n1177);
   U731 : MUXB2DL port map( A0 => n1541, A1 => b(8), SL => n63, Z => n874);
   U732 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n875, Z => n1178);
   U733 : MUXB2DL port map( A0 => b(8), A1 => n1543, SL => n63, Z => n875);
   U734 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n876, Z => n1179);
   U735 : MUXB2DL port map( A0 => b(7), A1 => n1545, SL => n63, Z => n876);
   U736 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n877, Z => n1180);
   U737 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n63, Z => n877);
   U738 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n878, Z => n1181);
   U739 : MUXB2DL port map( A0 => n1547, A1 => n1549, SL => n63, Z => n878);
   U740 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n879, Z => n1182);
   U741 : MUXB2DL port map( A0 => n1549, A1 => b(3), SL => n63, Z => n879);
   U742 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n880, Z => n1183);
   U743 : MUXB2DL port map( A0 => n1551, A1 => b(2), SL => n63, Z => n880);
   U744 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n881, Z => n1184);
   U745 : MUXB2DL port map( A0 => b(2), A1 => n1554, SL => n63, Z => n881);
   U746 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n882, Z => n1185);
   U747 : MUXB2DL port map( A0 => n1554, A1 => b(0), SL => n63, Z => n882);
   U748 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n883, Z => n1186);
   U749 : NAN2M1D1 port map( A1 => n63, A2 => n1556, Z => n883);
   U750 : NOR2M1D1 port map( A1 => n50, A2 => n53, Z => n1090);
   U751 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n884, Z => n1187);
   U752 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n56, Z => n884);
   U753 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n885, Z => n1188);
   U754 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n56, Z => n885);
   U755 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n886, Z => n1189);
   U756 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n56, Z => n886);
   U757 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n887, Z => n1190);
   U758 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n56, Z => n887);
   U759 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n888, Z => n1191);
   U760 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n56, Z => n888);
   U761 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n889, Z => n1192);
   U762 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n56, Z => n889);
   U763 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n890, Z => n1193);
   U764 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n56, Z => n890);
   U765 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n891, Z => n1194);
   U766 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n56, Z => n891);
   U767 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n892, Z => n1195);
   U768 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n56, Z => n892);
   U769 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n893, Z => n1196);
   U770 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n56, Z => n893);
   U771 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n894, Z => n1197);
   U772 : MUXB2DL port map( A0 => n1541, A1 => b(8), SL => n56, Z => n894);
   U773 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n895, Z => n1198);
   U774 : MUXB2DL port map( A0 => b(8), A1 => n1543, SL => n56, Z => n895);
   U775 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n896, Z => n1199);
   U776 : MUXB2DL port map( A0 => n1543, A1 => n1545, SL => n56, Z => n896);
   U777 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n897, Z => n1200);
   U778 : MUXB2DL port map( A0 => n1545, A1 => n1547, SL => n56, Z => n897);
   U779 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n898, Z => n1201);
   U780 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n56, Z => n898);
   U781 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n899, Z => n1202);
   U782 : MUXB2DL port map( A0 => n1549, A1 => n1551, SL => n56, Z => n899);
   U783 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n900, Z => n1203);
   U784 : MUXB2DL port map( A0 => n1551, A1 => b(2), SL => n56, Z => n900);
   U785 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n901, Z => n1204);
   U786 : MUXB2DL port map( A0 => b(2), A1 => n1554, SL => n56, Z => n901);
   U787 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n902, Z => n1205);
   U788 : MUXB2DL port map( A0 => n1554, A1 => n1556, SL => n56, Z => n902);
   U789 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n903, Z => n1206);
   U790 : NAN2M1D1 port map( A1 => n56, A2 => n1556, Z => n903);
   U791 : NOR2M1D1 port map( A1 => n42, A2 => n45, Z => n1091);
   U792 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n904, Z => n1207);
   U793 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n48, Z => n904);
   U794 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n905, Z => n1208);
   U795 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n48, Z => n905);
   U796 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n906, Z => n1209);
   U797 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n48, Z => n906);
   U798 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n907, Z => n1210);
   U799 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n48, Z => n907);
   U800 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n908, Z => n1211);
   U801 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n48, Z => n908);
   U802 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n909, Z => n1212);
   U803 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n48, Z => n909);
   U804 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n910, Z => n1213);
   U805 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n48, Z => n910);
   U806 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n911, Z => n1214);
   U807 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n48, Z => n911);
   U808 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n912, Z => n1215);
   U809 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n48, Z => n912);
   U810 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n913, Z => n1216);
   U811 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n48, Z => n913);
   U812 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n914, Z => n1217);
   U813 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n48, Z => n914);
   U814 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n915, Z => n1218);
   U815 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n48, Z => n915);
   U816 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n916, Z => n1219);
   U817 : MUXB2DL port map( A0 => n1541, A1 => b(8), SL => n48, Z => n916);
   U818 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n917, Z => n1220);
   U819 : MUXB2DL port map( A0 => b(8), A1 => n1543, SL => n48, Z => n917);
   U820 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n918, Z => n1221);
   U821 : MUXB2DL port map( A0 => b(7), A1 => n1545, SL => n48, Z => n918);
   U822 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n919, Z => n1222);
   U823 : MUXB2DL port map( A0 => n1545, A1 => n1547, SL => n48, Z => n919);
   U824 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n920, Z => n1223);
   U825 : MUXB2DL port map( A0 => n1547, A1 => b(4), SL => n48, Z => n920);
   U826 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n921, Z => n1224);
   U827 : MUXB2DL port map( A0 => b(4), A1 => n1551, SL => n48, Z => n921);
   U828 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n922, Z => n1225);
   U829 : MUXB2DL port map( A0 => n1551, A1 => b(2), SL => n48, Z => n922);
   U830 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n923, Z => n1226);
   U831 : MUXB2DL port map( A0 => b(2), A1 => n1554, SL => n48, Z => n923);
   U832 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n924, Z => n1227);
   U833 : MUXB2DL port map( A0 => n1554, A1 => n1556, SL => n48, Z => n924);
   U834 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n925, Z => n1228);
   U835 : NAN2M1D1 port map( A1 => n48, A2 => n1556, Z => n925);
   U836 : NOR2M1D1 port map( A1 => n1521, A2 => n38, Z => n1092);
   U837 : MUXB2DL port map( A0 => n1521, A1 => n38, SL => n926, Z => n1229);
   U838 : MUXB2DL port map( A0 => b(23), A1 => b(22), SL => n1518, Z => n926);
   U839 : MUXB2DL port map( A0 => n1521, A1 => n38, SL => n927, Z => n1230);
   U840 : MUXB2DL port map( A0 => b(22), A1 => b(21), SL => n1518, Z => n927);
   U841 : MUXB2DL port map( A0 => n1521, A1 => n38, SL => n928, Z => n1231);
   U842 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n1518, Z => n928);
   U843 : MUXB2DL port map( A0 => n1521, A1 => n38, SL => n929, Z => n1232);
   U844 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n1518, Z => n929);
   U845 : MUXB2DL port map( A0 => n1521, A1 => n38, SL => n930, Z => n1233);
   U846 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n1518, Z => n930);
   U847 : MUXB2DL port map( A0 => n1521, A1 => n38, SL => n931, Z => n1234);
   U848 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n1518, Z => n931);
   U849 : MUXB2DL port map( A0 => n1521, A1 => n38, SL => n932, Z => n1235);
   U850 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n1518, Z => n932);
   U851 : MUXB2DL port map( A0 => n1521, A1 => n38, SL => n933, Z => n1236);
   U852 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n1518, Z => n933);
   U853 : MUXB2DL port map( A0 => n1521, A1 => n38, SL => n934, Z => n1237);
   U854 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n1518, Z => n934);
   U855 : MUXB2DL port map( A0 => n1521, A1 => n38, SL => n935, Z => n1238);
   U856 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n1518, Z => n935);
   U857 : MUXB2DL port map( A0 => n1521, A1 => n38, SL => n936, Z => n1239);
   U858 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n1518, Z => n936);
   U859 : MUXB2DL port map( A0 => n1521, A1 => n38, SL => n937, Z => n1240);
   U860 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n1518, Z => n937);
   U861 : MUXB2DL port map( A0 => n1521, A1 => n38, SL => n938, Z => n1241);
   U862 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n1518, Z => n938);
   U863 : MUXB2DL port map( A0 => n1521, A1 => n38, SL => n939, Z => n1242);
   U864 : MUXB2DL port map( A0 => b(10), A1 => n1541, SL => n1518, Z => n939);
   U865 : MUXB2DL port map( A0 => n1521, A1 => n38, SL => n940, Z => n1243);
   U866 : MUXB2DL port map( A0 => n1541, A1 => b(8), SL => n1518, Z => n940);
   U867 : MUXB2DL port map( A0 => n1521, A1 => n38, SL => n941, Z => n1244);
   U868 : MUXB2DL port map( A0 => b(8), A1 => n1543, SL => n1518, Z => n941);
   U869 : MUXB2DL port map( A0 => n1521, A1 => n38, SL => n942, Z => n1245);
   U870 : MUXB2DL port map( A0 => b(7), A1 => n1545, SL => n1518, Z => n942);
   U871 : MUXB2DL port map( A0 => n1521, A1 => n38, SL => n943, Z => n1246);
   U872 : MUXB2DL port map( A0 => b(6), A1 => n1547, SL => n1518, Z => n943);
   U873 : MUXB2DL port map( A0 => n1521, A1 => n38, SL => n944, Z => n1247);
   U874 : MUXB2DL port map( A0 => b(5), A1 => n1549, SL => n1518, Z => n944);
   U875 : MUXB2DL port map( A0 => n1521, A1 => n38, SL => n945, Z => n1248);
   U876 : MUXB2DL port map( A0 => b(4), A1 => n1551, SL => n1518, Z => n945);
   U877 : MUXB2DL port map( A0 => n1521, A1 => n38, SL => n946, Z => n1249);
   U878 : MUXB2DL port map( A0 => n1551, A1 => b(2), SL => n1518, Z => n946);
   U879 : MUXB2DL port map( A0 => n1521, A1 => n38, SL => n947, Z => n1250);
   U880 : MUXB2DL port map( A0 => b(2), A1 => n1554, SL => n1518, Z => n947);
   U881 : MUXB2DL port map( A0 => n1521, A1 => n38, SL => n948, Z => n1251);
   U882 : MUXB2DL port map( A0 => n1553, A1 => n1556, SL => n1518, Z => n948);
   U883 : MUXB2DL port map( A0 => n1521, A1 => n38, SL => n949, Z => n1252);
   U884 : NAN2M1D1 port map( A1 => n1518, A2 => n1556, Z => n949);
   U886 : MUXB2DL port map( A0 => n1538, A1 => n30, SL => n950, Z => n1253);
   U887 : MUXB2DL port map( A0 => b(25), A1 => b(24), SL => n1517, Z => n950);
   U888 : MUXB2DL port map( A0 => n1538, A1 => n30, SL => n951, Z => n1254);
   U889 : MUXB2DL port map( A0 => b(24), A1 => b(23), SL => n1517, Z => n951);
   U890 : MUXB2DL port map( A0 => n1538, A1 => n30, SL => n952, Z => n1255);
   U891 : MUXB2DL port map( A0 => b(23), A1 => b(22), SL => n1517, Z => n952);
   U892 : MUXB2DL port map( A0 => n1538, A1 => n30, SL => n953, Z => n1256);
   U893 : MUXB2DL port map( A0 => b(22), A1 => b(21), SL => n1517, Z => n953);
   U894 : MUXB2DL port map( A0 => n1538, A1 => n30, SL => n954, Z => n1257);
   U895 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n1517, Z => n954);
   U896 : MUXB2DL port map( A0 => n1538, A1 => n30, SL => n955, Z => n1258);
   U897 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n1517, Z => n955);
   U898 : MUXB2DL port map( A0 => n1538, A1 => n30, SL => n956, Z => n1259);
   U899 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n1517, Z => n956);
   U900 : MUXB2DL port map( A0 => n1538, A1 => n30, SL => n957, Z => n1260);
   U901 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n1517, Z => n957);
   U902 : MUXB2DL port map( A0 => n1538, A1 => n30, SL => n958, Z => n1261);
   U903 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n1517, Z => n958);
   U904 : MUXB2DL port map( A0 => n1538, A1 => n30, SL => n959, Z => n1262);
   U905 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n1517, Z => n959);
   U906 : MUXB2DL port map( A0 => n1538, A1 => n30, SL => n960, Z => n1263);
   U907 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n1517, Z => n960);
   U908 : MUXB2DL port map( A0 => n1538, A1 => n30, SL => n961, Z => n1264);
   U909 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n1517, Z => n961);
   U910 : MUXB2DL port map( A0 => n1538, A1 => n30, SL => n962, Z => n1265);
   U911 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n1517, Z => n962);
   U912 : MUXB2DL port map( A0 => n1538, A1 => n30, SL => n963, Z => n1266);
   U913 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n1517, Z => n963);
   U914 : MUXB2DL port map( A0 => n1538, A1 => n30, SL => n964, Z => n1267);
   U915 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n1517, Z => n964);
   U916 : MUXB2DL port map( A0 => n1538, A1 => n30, SL => n965, Z => n1268);
   U917 : MUXB2DL port map( A0 => b(10), A1 => n1541, SL => n1517, Z => n965);
   U918 : MUXB2DL port map( A0 => n1538, A1 => n30, SL => n966, Z => n1269);
   U919 : MUXB2DL port map( A0 => n1541, A1 => b(8), SL => n1517, Z => n966);
   U920 : MUXB2DL port map( A0 => n1538, A1 => n30, SL => n967, Z => n1270);
   U921 : MUXB2DL port map( A0 => b(8), A1 => n1543, SL => n1517, Z => n967);
   U922 : MUXB2DL port map( A0 => n1538, A1 => n30, SL => n968, Z => n1271);
   U923 : MUXB2DL port map( A0 => b(7), A1 => n1545, SL => n1517, Z => n968);
   U924 : MUXB2DL port map( A0 => n1538, A1 => n30, SL => n969, Z => n1272);
   U925 : MUXB2DL port map( A0 => b(6), A1 => n1547, SL => n1517, Z => n969);
   U926 : MUXB2DL port map( A0 => n1538, A1 => n30, SL => n970, Z => n1273);
   U927 : MUXB2DL port map( A0 => b(5), A1 => n1549, SL => n1517, Z => n970);
   U928 : MUXB2DL port map( A0 => n1538, A1 => n30, SL => n971, Z => n1274);
   U929 : MUXB2DL port map( A0 => b(4), A1 => n1551, SL => n1517, Z => n971);
   U930 : MUXB2DL port map( A0 => n1538, A1 => n30, SL => n972, Z => n1275);
   U931 : MUXB2DL port map( A0 => n1551, A1 => b(2), SL => n1517, Z => n972);
   U932 : MUXB2DL port map( A0 => n1538, A1 => n30, SL => n973, Z => n1276);
   U933 : MUXB2DL port map( A0 => b(2), A1 => n1554, SL => n1517, Z => n973);
   U934 : MUXB2DL port map( A0 => n1538, A1 => n30, SL => n974, Z => n1277);
   U935 : MUXB2DL port map( A0 => n1553, A1 => n1556, SL => n1517, Z => n974);
   U936 : MUXB2DL port map( A0 => n1538, A1 => n30, SL => n975, Z => n1278);
   U937 : NAN2M1D1 port map( A1 => n1517, A2 => n1556, Z => n975);
   U938 : NOR2M1D1 port map( A1 => n1520, A2 => n22, Z => n1094);
   U939 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n976, Z => n1279);
   U940 : MUXB2DL port map( A0 => b(27), A1 => b(26), SL => n1539, Z => n976);
   U941 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n977, Z => n1280);
   U942 : MUXB2DL port map( A0 => b(26), A1 => b(25), SL => n1539, Z => n977);
   U943 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n978, Z => n1281);
   U944 : MUXB2DL port map( A0 => b(25), A1 => b(24), SL => n1539, Z => n978);
   U945 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n979, Z => n1282);
   U946 : MUXB2DL port map( A0 => b(24), A1 => b(23), SL => n1539, Z => n979);
   U947 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n980, Z => n1283);
   U948 : MUXB2DL port map( A0 => b(23), A1 => b(22), SL => n1539, Z => n980);
   U949 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n981, Z => n1284);
   U950 : MUXB2DL port map( A0 => b(22), A1 => b(21), SL => n1539, Z => n981);
   U951 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n982, Z => n1285);
   U952 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n1539, Z => n982);
   U953 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n983, Z => n1286);
   U954 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n1539, Z => n983);
   U955 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n984, Z => n1287);
   U956 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n1539, Z => n984);
   U957 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n985, Z => n1288);
   U958 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n1539, Z => n985);
   U959 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n986, Z => n1289);
   U960 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n1539, Z => n986);
   U961 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n987, Z => n1290);
   U962 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n1539, Z => n987);
   U963 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n988, Z => n1291);
   U964 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n1539, Z => n988);
   U965 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n989, Z => n1292);
   U966 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n1539, Z => n989);
   U967 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n990, Z => n1293);
   U968 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n1539, Z => n990);
   U969 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n991, Z => n1294);
   U970 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n1539, Z => n991);
   U971 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n992, Z => n1295);
   U972 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n1539, Z => n992);
   U973 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n993, Z => n1296);
   U974 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n1539, Z => n993);
   U975 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n994, Z => n1297);
   U976 : MUXB2DL port map( A0 => n1541, A1 => b(8), SL => n1539, Z => n994);
   U977 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n995, Z => n1298);
   U978 : MUXB2DL port map( A0 => b(8), A1 => n1543, SL => n1539, Z => n995);
   U979 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n996, Z => n1299);
   U980 : MUXB2DL port map( A0 => b(7), A1 => n1545, SL => n1539, Z => n996);
   U981 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n997, Z => n1300);
   U982 : MUXB2DL port map( A0 => b(6), A1 => n1547, SL => n1539, Z => n997);
   U983 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n998, Z => n1301);
   U984 : MUXB2DL port map( A0 => b(5), A1 => n1549, SL => n1539, Z => n998);
   U985 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n999, Z => n1302);
   U986 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n1539, Z => n999);
   U987 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n1000, Z => n1303);
   U988 : MUXB2DL port map( A0 => n1551, A1 => b(2), SL => n1539, Z => n1000);
   U989 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n1001, Z => n1304);
   U990 : MUXB2DL port map( A0 => b(2), A1 => n1554, SL => n1539, Z => n1001);
   U991 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n1002, Z => n1305);
   U992 : MUXB2DL port map( A0 => n1553, A1 => n1556, SL => n1539, Z => n1002);
   U993 : MUXB2DL port map( A0 => n1520, A1 => n22, SL => n1003, Z => n1306);
   U994 : NAN2M1D1 port map( A1 => n1539, A2 => n1556, Z => n1003);
   U995 : NOR2M1D1 port map( A1 => n1519, A2 => n14, Z => n1095);
   U996 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1004, Z => n1307);
   U997 : MUXB2DL port map( A0 => b(29), A1 => b(28), SL => n1540, Z => n1004);
   U998 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1005, Z => n1308);
   U999 : MUXB2DL port map( A0 => b(28), A1 => b(27), SL => n1540, Z => n1005);
   U1000 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1006, Z => n1309);
   U1001 : MUXB2DL port map( A0 => b(27), A1 => b(26), SL => n1540, Z => n1006)
                           ;
   U1002 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1007, Z => n1310);
   U1003 : MUXB2DL port map( A0 => b(26), A1 => b(25), SL => n1540, Z => n1007)
                           ;
   U1004 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1008, Z => n1311);
   U1005 : MUXB2DL port map( A0 => b(25), A1 => b(24), SL => n1540, Z => n1008)
                           ;
   U1006 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1009, Z => n1312);
   U1007 : MUXB2DL port map( A0 => b(24), A1 => b(23), SL => n1540, Z => n1009)
                           ;
   U1008 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1010, Z => n1313);
   U1009 : MUXB2DL port map( A0 => b(23), A1 => b(22), SL => n1540, Z => n1010)
                           ;
   U1010 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1011, Z => n1314);
   U1011 : MUXB2DL port map( A0 => b(22), A1 => b(21), SL => n1540, Z => n1011)
                           ;
   U1012 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1012, Z => n1315);
   U1013 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n1540, Z => n1012)
                           ;
   U1014 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1013, Z => n1316);
   U1015 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n1540, Z => n1013)
                           ;
   U1016 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1014, Z => n1317);
   U1017 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n1540, Z => n1014)
                           ;
   U1018 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1015, Z => n1318);
   U1019 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n1540, Z => n1015)
                           ;
   U1020 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1016, Z => n1319);
   U1021 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n1540, Z => n1016)
                           ;
   U1022 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1017, Z => n1320);
   U1023 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n1540, Z => n1017)
                           ;
   U1024 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1018, Z => n1321);
   U1025 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n1540, Z => n1018)
                           ;
   U1026 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1019, Z => n1322);
   U1027 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n1540, Z => n1019)
                           ;
   U1028 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1020, Z => n1323);
   U1029 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n1540, Z => n1020)
                           ;
   U1030 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1021, Z => n1324);
   U1031 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n1540, Z => n1021)
                           ;
   U1032 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1022, Z => n1325);
   U1033 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n1540, Z => n1022)
                           ;
   U1034 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1023, Z => n1326);
   U1035 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n1540, Z => n1023);
   U1036 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1024, Z => n1327);
   U1037 : MUXB2DL port map( A0 => n1541, A1 => b(8), SL => n1540, Z => n1024);
   U1038 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1025, Z => n1328);
   U1039 : MUXB2DL port map( A0 => b(8), A1 => n1543, SL => n1540, Z => n1025);
   U1040 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1026, Z => n1329);
   U1041 : MUXB2DL port map( A0 => n1543, A1 => n1545, SL => n1540, Z => n1026)
                           ;
   U1042 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1027, Z => n1330);
   U1043 : MUXB2DL port map( A0 => b(6), A1 => n1547, SL => n1540, Z => n1027);
   U1044 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1028, Z => n1331);
   U1045 : MUXB2DL port map( A0 => b(5), A1 => n1549, SL => n1540, Z => n1028);
   U1046 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1029, Z => n1332);
   U1047 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n1540, Z => n1029);
   U1048 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1030, Z => n1333);
   U1049 : MUXB2DL port map( A0 => n1551, A1 => b(2), SL => n1540, Z => n1030);
   U1050 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1031, Z => n1334);
   U1051 : MUXB2DL port map( A0 => b(2), A1 => n1554, SL => n1540, Z => n1031);
   U1052 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1032, Z => n1335);
   U1053 : MUXB2DL port map( A0 => n1553, A1 => b(0), SL => n1540, Z => n1032);
   U1054 : MUXB2DL port map( A0 => n1519, A1 => n14, SL => n1033, Z => n1336);
   U1055 : NAN2M1D1 port map( A1 => n1540, A2 => n1556, Z => n1033);
   U1056 : NOR2M1D1 port map( A1 => n3, A2 => n6, Z => n1096);
   U1057 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1034, Z => n1337);
   U1058 : MUXB2DL port map( A0 => b(31), A1 => b(30), SL => n8, Z => n1034);
   U1059 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1035, Z => n1338);
   U1060 : MUXB2DL port map( A0 => b(30), A1 => b(29), SL => n8, Z => n1035);
   U1061 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1036, Z => n1339);
   U1062 : MUXB2DL port map( A0 => b(29), A1 => b(28), SL => n8, Z => n1036);
   U1063 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1037, Z => n1340);
   U1064 : MUXB2DL port map( A0 => b(28), A1 => b(27), SL => n8, Z => n1037);
   U1065 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1038, Z => n1341);
   U1066 : MUXB2DL port map( A0 => b(27), A1 => b(26), SL => n8, Z => n1038);
   U1067 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1039, Z => n1342);
   U1068 : MUXB2DL port map( A0 => b(26), A1 => b(25), SL => n8, Z => n1039);
   U1069 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1040, Z => n1343);
   U1070 : MUXB2DL port map( A0 => b(25), A1 => b(24), SL => n8, Z => n1040);
   U1071 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1041, Z => n1344);
   U1072 : MUXB2DL port map( A0 => b(24), A1 => b(23), SL => n8, Z => n1041);
   U1073 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1042, Z => n1345);
   U1074 : MUXB2DL port map( A0 => b(23), A1 => b(22), SL => n8, Z => n1042);
   U1075 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1043, Z => n1346);
   U1076 : MUXB2DL port map( A0 => b(22), A1 => b(21), SL => n8, Z => n1043);
   U1077 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1044, Z => n1347);
   U1078 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n8, Z => n1044);
   U1079 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1045, Z => n1348);
   U1080 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n8, Z => n1045);
   U1081 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1046, Z => n1349);
   U1082 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n8, Z => n1046);
   U1083 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1047, Z => n1350);
   U1084 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n8, Z => n1047);
   U1085 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1048, Z => n1351);
   U1086 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n8, Z => n1048);
   U1087 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1049, Z => n1352);
   U1088 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n8, Z => n1049);
   U1089 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1050, Z => n1353);
   U1090 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n8, Z => n1050);
   U1091 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1051, Z => n1354);
   U1092 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n8, Z => n1051);
   U1093 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1052, Z => n1355);
   U1094 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n8, Z => n1052);
   U1095 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1053, Z => n1356);
   U1096 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n8, Z => n1053);
   U1097 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1054, Z => n1357);
   U1098 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n8, Z => n1054);
   U1099 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1055, Z => n1358);
   U1100 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n8, Z => n1055);
   U1101 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1056, Z => n1359);
   U1102 : MUXB2DL port map( A0 => n1541, A1 => b(8), SL => n8, Z => n1056);
   U1103 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1057, Z => n1360);
   U1104 : MUXB2DL port map( A0 => b(8), A1 => n1543, SL => n8, Z => n1057);
   U1105 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1058, Z => n1361);
   U1106 : MUXB2DL port map( A0 => b(7), A1 => n1545, SL => n8, Z => n1058);
   U1107 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1059, Z => n1362);
   U1108 : MUXB2DL port map( A0 => b(6), A1 => n1547, SL => n8, Z => n1059);
   U1109 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1060, Z => n1363);
   U1110 : MUXB2DL port map( A0 => b(5), A1 => n1549, SL => n8, Z => n1060);
   U1111 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1061, Z => n1364);
   U1112 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n8, Z => n1061);
   U1113 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1062, Z => n1365);
   U1114 : MUXB2DL port map( A0 => n1551, A1 => b(2), SL => n8, Z => n1062);
   U1115 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1063, Z => n1366);
   U1116 : MUXB2DL port map( A0 => b(2), A1 => n1554, SL => n8, Z => n1063);
   U1117 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1064, Z => n1367);
   U1118 : MUXB2DL port map( A0 => n1553, A1 => b(0), SL => n8, Z => n1064);
   U1119 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1065, Z => n1368);
   U1120 : NAN2M1D1 port map( A1 => n8, A2 => b(0), Z => n1065);
   U1121 : OAI21D1 port map( A1 => a(29), A2 => a(30), B => n1066, Z => n104);
   U1123 : EXNOR2D1 port map( A1 => a(29), A2 => a(30), Z => n106);
   U1125 : OAI21D1 port map( A1 => a(27), A2 => a(28), B => n1067, Z => n99);
   U1127 : EXNOR2D1 port map( A1 => a(27), A2 => a(28), Z => n103);
   U1129 : OAI21D1 port map( A1 => a(25), A2 => a(26), B => n1068, Z => n94);
   U1131 : EXNOR2D1 port map( A1 => a(25), A2 => a(26), Z => n98);
   U1135 : EXNOR2D1 port map( A1 => a(23), A2 => a(24), Z => n93);
   U1186 : ADHALFDL port map( A => n1278, B => n1093, CO => n780, S => n781);
   U1187 : EXNOR2D1 port map( A1 => a(5), A2 => a(6), Z => n1517);
   U1188 : EXNOR2D1 port map( A1 => a(7), A2 => a(8), Z => n1518);
   U1189 : OAI21D1 port map( A1 => a(1), A2 => a(2), B => n1080, Z => n1519);
   U1190 : OAI21D1 port map( A1 => a(3), A2 => a(4), B => n1079, Z => n1520);
   U1191 : OAI21D1 port map( A1 => a(7), A2 => a(8), B => n1077, Z => n1521);
   U1192 : AND2D1 port map( A1 => n1524, A2 => n305, Z => product(0));
   U1193 : AO21D1 port map( A1 => n215, A2 => n187, B => n188, Z => n1523);
   U1194 : OR2D1 port map( A1 => n1368, A2 => n1096, Z => n1524);
   U1195 : OA21M20D1 port map( A1 => n1525, A2 => n197, B => n194, Z => n190);
   U1196 : INVD1 port map( A => n215, Z => n214);
   U1197 : INVD1 port map( A => n233, Z => n232);
   U1198 : NAN2D1 port map( A1 => n313, A2 => n231, Z => n162);
   U1199 : INVD1 port map( A => n242, Z => n241);
   U1200 : INVD1 port map( A => n255, Z => n254);
   U1201 : INVD1 port map( A => n230, Z => n313);
   U1202 : INVD1 port map( A => n231, Z => n229);
   U1203 : INVD1 port map( A => n264, Z => n263);
   U1204 : NAN2D1 port map( A1 => n223, A2 => n1530, Z => n216);
   U1205 : INVD1 port map( A => n221, Z => n219);
   U1206 : NAN2D1 port map( A1 => n1532, A2 => n1531, Z => n243);
   U1207 : INVD1 port map( A => n248, Z => n246);
   U1208 : NAN2D1 port map( A1 => n1526, A2 => n1529, Z => n265);
   U1209 : INVD1 port map( A => n270, Z => n268);
   U1210 : NOR2D1 port map( A1 => n258, A2 => n261, Z => n256);
   U1211 : NOR2D1 port map( A1 => n236, A2 => n239, Z => n234);
   U1212 : NOR2D1 port map( A1 => n189, A2 => n201, Z => n187);
   U1213 : INVD1 port map( A => n209, Z => n211);
   U1214 : INVD1 port map( A => n206, Z => n204);
   U1215 : INVD1 port map( A => n275, Z => n273);
   U1216 : OR2D1 port map( A1 => n553, A2 => n574, Z => n1525);
   U1217 : NAN2D1 port map( A1 => n1525, A2 => n1528, Z => n189);
   U1218 : INVD1 port map( A => n199, Z => n197);
   U1219 : NAN2D1 port map( A1 => n667, A2 => n682, Z => n231);
   U1220 : INVD1 port map( A => n253, Z => n251);
   U1221 : NOR2D1 port map( A1 => n225, A2 => n230, Z => n223);
   U1222 : NAN2D1 port map( A1 => n1527, A2 => n310, Z => n201);
   U1223 : NOR2D1 port map( A1 => n683, A2 => n696, Z => n236);
   U1224 : NAN2D1 port map( A1 => n553, A2 => n574, Z => n194);
   U1225 : NOR2D1 port map( A1 => n667, A2 => n682, Z => n230);
   U1226 : INVD1 port map( A => n208, Z => n310);
   U1227 : NAN2D1 port map( A1 => n683, A2 => n696, Z => n237);
   U1228 : NAN2D1 port map( A1 => n1525, A2 => n194, Z => n156);
   U1229 : NAN2D1 port map( A1 => n1528, A2 => n199, Z => n157);
   U1230 : NAN2D1 port map( A1 => n1527, A2 => n206, Z => n158);
   U1231 : NAN2D1 port map( A1 => n310, A2 => n209, Z => n159);
   U1232 : NAN2D1 port map( A1 => n312, A2 => n226, Z => n161);
   U1233 : INVD1 port map( A => n225, Z => n312);
   U1234 : NAN2D1 port map( A1 => n1530, A2 => n221, Z => n160);
   U1235 : NAN2D1 port map( A1 => n314, A2 => n237, Z => n163);
   U1236 : INVD1 port map( A => n236, Z => n314);
   U1237 : NAN2D1 port map( A1 => n1532, A2 => n248, Z => n165);
   U1238 : NAN2D1 port map( A1 => n315, A2 => n240, Z => n164);
   U1239 : INVD1 port map( A => n239, Z => n315);
   U1240 : NAN2D1 port map( A1 => n1531, A2 => n253, Z => n166);
   U1241 : NAN2D1 port map( A1 => n318, A2 => n259, Z => n167);
   U1242 : INVD1 port map( A => n258, Z => n318);
   U1243 : NAN2D1 port map( A1 => n319, A2 => n262, Z => n168);
   U1244 : INVD1 port map( A => n261, Z => n319);
   U1245 : INVD1 port map( A => n277, Z => n276);
   U1246 : NAN2D1 port map( A1 => n1526, A2 => n270, Z => n169);
   U1247 : NAN2D1 port map( A1 => n1529, A2 => n275, Z => n170);
   U1248 : INVD1 port map( A => n286, Z => n285);
   U1249 : OR2D1 port map( A1 => n755, A2 => n762, Z => n1526);
   U1250 : NAN2D1 port map( A1 => n755, A2 => n762, Z => n270);
   U1251 : NOR2D1 port map( A1 => n280, A2 => n283, Z => n278);
   U1252 : OA21M20D1 port map( A1 => n1533, A2 => n294, B => n293, Z => n289);
   U1253 : NOR2D1 port map( A1 => n651, A2 => n666, Z => n225);
   U1254 : OA21M20D1 port map( A1 => n1534, A2 => n302, B => n301, Z => n297);
   U1255 : OR2D1 port map( A1 => n595, A2 => n614, Z => n1527);
   U1256 : NOR2D1 port map( A1 => n771, A2 => n776, Z => n280);
   U1257 : NOR2D1 port map( A1 => n745, A2 => n754, Z => n261);
   U1258 : NOR2D1 port map( A1 => n735, A2 => n744, Z => n258);
   U1259 : NAN2D1 port map( A1 => n763, A2 => n770, Z => n275);
   U1260 : OR2D1 port map( A1 => n575, A2 => n594, Z => n1528);
   U1261 : NAN2D1 port map( A1 => n575, A2 => n594, Z => n199);
   U1262 : NAN2D1 port map( A1 => n723, A2 => n734, Z => n253);
   U1263 : NAN2D1 port map( A1 => n651, A2 => n666, Z => n226);
   U1264 : OR2D1 port map( A1 => n763, A2 => n770, Z => n1529);
   U1265 : NAN2D1 port map( A1 => n595, A2 => n614, Z => n206);
   U1266 : OR2D1 port map( A1 => n633, A2 => n650, Z => n1530);
   U1267 : NAN2D1 port map( A1 => n745, A2 => n754, Z => n262);
   U1268 : OR2D1 port map( A1 => n723, A2 => n734, Z => n1531);
   U1269 : OR2D1 port map( A1 => n711, A2 => n722, Z => n1532);
   U1270 : NAN2D1 port map( A1 => n771, A2 => n776, Z => n281);
   U1271 : NAN2D1 port map( A1 => n615, A2 => n632, Z => n209);
   U1272 : NAN2D1 port map( A1 => n735, A2 => n744, Z => n259);
   U1273 : NOR2D1 port map( A1 => n697, A2 => n710, Z => n239);
   U1274 : NOR2D1 port map( A1 => n615, A2 => n632, Z => n208);
   U1275 : NAN2D1 port map( A1 => n633, A2 => n650, Z => n221);
   U1276 : NAN2D1 port map( A1 => n711, A2 => n722, Z => n248);
   U1277 : NAN2D1 port map( A1 => n697, A2 => n710, Z => n240);
   U1278 : NAN2D1 port map( A1 => n322, A2 => n281, Z => n171);
   U1279 : INVD1 port map( A => n280, Z => n322);
   U1280 : NAN2D1 port map( A1 => n323, A2 => n284, Z => n172);
   U1281 : INVD1 port map( A => n283, Z => n323);
   U1282 : NAN2D1 port map( A1 => n324, A2 => n288, Z => n173);
   U1283 : INVD1 port map( A => n287, Z => n324);
   U1284 : NAN2D1 port map( A1 => n1533, A2 => n293, Z => n174);
   U1285 : NAN2D1 port map( A1 => n326, A2 => n296, Z => n175);
   U1286 : INVD1 port map( A => n295, Z => n326);
   U1287 : NAN2D1 port map( A1 => n1534, A2 => n301, Z => n176);
   U1288 : EXOR2D1 port map( A1 => n178, A2 => n155, Z => product(31));
   U1289 : EXOR2D1 port map( A1 => n329, A2 => n344, Z => n155);
   U1290 : OR2D1 port map( A1 => n787, A2 => n789, Z => n1533);
   U1291 : OR2D1 port map( A1 => n793, A2 => n1366, Z => n1534);
   U1292 : NOR2D1 port map( A1 => n777, A2 => n782, Z => n283);
   U1293 : NAN2D1 port map( A1 => n787, A2 => n789, Z => n293);
   U1294 : NAN2D1 port map( A1 => n793, A2 => n1366, Z => n301);
   U1295 : NAN2D1 port map( A1 => n777, A2 => n782, Z => n284);
   U1296 : NOR2D1 port map( A1 => n783, A2 => n786, Z => n287);
   U1297 : NOR2D1 port map( A1 => n791, A2 => n792, Z => n295);
   U1298 : NAN2D1 port map( A1 => n783, A2 => n786, Z => n288);
   U1299 : NAN2D1 port map( A1 => n791, A2 => n792, Z => n296);
   U1300 : NAN2D1 port map( A1 => n1368, A2 => n1096, Z => n305);
   U1301 : NOR2D1 port map( A1 => n303, A2 => n305, Z => n302);
   U1302 : ADHALFDL port map( A => n1329, B => n1359, CO => n760, S => n761);
   U1303 : INVD1 port map( A => n1535, Z => n1540);
   U1304 : ADHALFDL port map( A => n1335, B => n1365, CO => n790, S => n791);
   U1305 : ADHALFDL port map( A => n1336, B => n1095, CO => n792, S => n793);
   U1306 : NOR2D1 port map( A1 => n1537, A2 => n30, Z => n1093);
   U1307 : INVD1 port map( A => n1536, Z => n1539);
   U1308 : ADHALFDL port map( A => n1331, B => n1361, CO => n774, S => n775);
   U1309 : ADHALFDL port map( A => n1252, B => n1092, CO => n768, S => n769);
   U1310 : ADHALFDL port map( A => n1333, B => n1363, CO => n784, S => n785);
   U1311 : ADHALFDL port map( A => n1306, B => n1094, CO => n788, S => n789);
   U1312 : INVD1 port map( A => n1537, Z => n1538);
   U1313 : INVD1 port map( A => n1546, Z => n1545);
   U1314 : INVD1 port map( A => n1542, Z => n1541);
   U1315 : INVD1 port map( A => n1548, Z => n1547);
   U1316 : INVD1 port map( A => n1555, Z => n1554);
   U1317 : INVD1 port map( A => n1544, Z => n1543);
   U1318 : INVD1 port map( A => n1552, Z => n1551);
   U1319 : INVD1 port map( A => n1550, Z => n1549);
   U1320 : INVD1 port map( A => n1555, Z => n1553);
   U1321 : INVD1 port map( A => n1557, Z => n1556);
   U1322 : ADHALFDL port map( A => n1206, B => n1090, CO => n732, S => n733);
   U1323 : ADHALFDL port map( A => n1168, B => n1088, CO => n680, S => n681);
   U1324 : ADHALFDL port map( A => n1152, B => n1087, CO => n648, S => n649);
   U1325 : ADHALFDL port map( A => n1228, B => n1091, CO => n752, S => n753);
   U1326 : ADHALFDL port map( A => n1186, B => n1089, CO => n708, S => n709);
   U1327 : ADHALFDL port map( A => n1138, B => n1086, CO => n612, S => n613);
   U1328 : INVD1 port map( A => n1367, Z => n303);
   U1329 : ADHALFDL port map( A => n1126, B => n1085, CO => n572, S => n573);
   U1330 : ADHALFDL port map( A => n1116, B => n1084, CO => n528, S => n529);
   U1331 : ADHALFDL port map( A => n1108, B => n1083, CO => n480, S => n481);
   U1332 : ADHALFDL port map( A => n1102, B => n1082, CO => n428, S => n429);
   U1333 : EXOR2D1 port map( A1 => n1307, A2 => n1337, Z => n343);
   U1334 : ADHALFDL port map( A => n1098, B => n1081, CO => n372, S => n373);
   U1335 : EXOR2D1 port map( A1 => a(1), A2 => a(2), Z => n1535);
   U1336 : ADHALFDL port map( A => n1323, B => n1353, CO => n694, S => n695);
   U1337 : EXOR2D1 port map( A1 => a(3), A2 => a(4), Z => n1536);
   U1338 : ADHALFDL port map( A => n1317, B => n1347, CO => n592, S => n593);
   U1339 : ADHALFDL port map( A => n1327, B => n1357, CO => n742, S => n743);
   U1340 : ADHALFDL port map( A => n1319, B => n1349, CO => n630, S => n631);
   U1341 : ADHALFDL port map( A => n1321, B => n1351, CO => n664, S => n665);
   U1342 : ADHALFDL port map( A => n1325, B => n1355, CO => n720, S => n721);
   U1343 : OA21D1 port map( A1 => a(5), A2 => a(6), B => n1078, Z => n1537);
   U1344 : INVD1 port map( A => b(6), Z => n1546);
   U1345 : INVD1 port map( A => b(7), Z => n1544);
   U1346 : INVD1 port map( A => a(3), Z => n1080);
   U1347 : EXNOR2D1 port map( A1 => a(11), A2 => a(12), Z => n56);
   U1348 : INVD1 port map( A => b(9), Z => n1542);
   U1349 : INVD1 port map( A => a(7), Z => n1078);
   U1350 : INVD1 port map( A => b(5), Z => n1548);
   U1351 : INVD1 port map( A => b(1), Z => n1555);
   U1352 : NAN2D1 port map( A1 => a(0), A2 => n6, Z => n3);
   U1353 : INVD1 port map( A => a(1), Z => n6);
   U1354 : INVD1 port map( A => a(9), Z => n1077);
   U1355 : INVD1 port map( A => b(3), Z => n1552);
   U1356 : INVD1 port map( A => b(4), Z => n1550);
   U1357 : EXNOR2D1 port map( A1 => a(13), A2 => a(14), Z => n63);
   U1358 : EXNOR2D1 port map( A1 => a(15), A2 => a(16), Z => n71);
   U1359 : INVD1 port map( A => b(0), Z => n1557);
   U1360 : INVD1 port map( A => a(5), Z => n1079);
   U1361 : EXNOR2D1 port map( A1 => a(9), A2 => a(10), Z => n48);
   U1362 : EXNOR2D1 port map( A1 => a(17), A2 => a(18), Z => n78);
   U1363 : AO21D1 port map( A1 => a(1), A2 => a(2), B => n1080, Z => n14);
   U1364 : AO21D1 port map( A1 => a(5), A2 => a(6), B => n1078, Z => n30);
   U1365 : EXNOR2D1 port map( A1 => a(19), A2 => a(20), Z => n83);
   U1366 : INVD1 port map( A => a(0), Z => n8);
   U1367 : AO21D1 port map( A1 => a(11), A2 => a(12), B => n1075, Z => n53);
   U1368 : INVD1 port map( A => a(13), Z => n1075);
   U1369 : ADHALFDL port map( A => n1315, B => n1345, CO => n550, S => n551);
   U1370 : AO21D1 port map( A1 => a(3), A2 => a(4), B => n1079, Z => n22);
   U1371 : AO21D1 port map( A1 => a(7), A2 => a(8), B => n1077, Z => n38);
   U1372 : OAI21D1 port map( A1 => a(11), A2 => a(12), B => n1075, Z => n50);
   U1373 : AO21D1 port map( A1 => a(13), A2 => a(14), B => n1074, Z => n61);
   U1374 : AO21D1 port map( A1 => a(15), A2 => a(16), B => n1073, Z => n69);
   U1375 : INVD1 port map( A => a(15), Z => n1074);
   U1376 : OAI21D1 port map( A1 => a(13), A2 => a(14), B => n1074, Z => n58);
   U1377 : INVD1 port map( A => a(17), Z => n1073);
   U1378 : OAI21D1 port map( A1 => a(15), A2 => a(16), B => n1073, Z => n66);
   U1379 : AO21D1 port map( A1 => a(9), A2 => a(10), B => n1076, Z => n45);
   U1380 : INVD1 port map( A => a(11), Z => n1076);
   U1381 : OAI21D1 port map( A1 => a(17), A2 => a(18), B => n1072, Z => n73);
   U1382 : INVD1 port map( A => a(19), Z => n1072);
   U1383 : OAI21D1 port map( A1 => a(9), A2 => a(10), B => n1076, Z => n42);
   U1384 : AO21D1 port map( A1 => a(17), A2 => a(18), B => n1072, Z => n76);
   U1385 : EXNOR2D1 port map( A1 => a(21), A2 => a(22), Z => n88);
   U1386 : OAI21D1 port map( A1 => a(19), A2 => a(20), B => n1071, Z => n79);
   U1387 : INVD1 port map( A => a(21), Z => n1071);
   U1388 : AO21D1 port map( A1 => a(19), A2 => a(20), B => n1071, Z => n81);
   U1389 : OAI21D1 port map( A1 => a(21), A2 => a(22), B => n1070, Z => n84);
   U1390 : INVD1 port map( A => a(23), Z => n1070);
   U1391 : AO21D1 port map( A1 => a(21), A2 => a(22), B => n1070, Z => n86);
   U1392 : ADHALFDL port map( A => n1313, B => n1343, CO => n504, S => n505);
   U1393 : OAI21D1 port map( A1 => a(23), A2 => a(24), B => n1069, Z => n89);
   U1394 : ADHALFDL port map( A => n1311, B => n1341, CO => n454, S => n455);
   U1395 : INVD1 port map( A => a(25), Z => n1069);
   U1396 : AO21D1 port map( A1 => a(23), A2 => a(24), B => n1069, Z => n91);
   U1397 : ADHALFDL port map( A => n1309, B => n1339, CO => n400, S => n401);
   U1398 : AO21D1 port map( A1 => a(25), A2 => a(26), B => n1068, Z => n96);
   U1399 : INVD1 port map( A => a(27), Z => n1068);
   U1400 : AO21D1 port map( A1 => a(27), A2 => a(28), B => n1067, Z => n101);
   U1401 : INVD1 port map( A => a(29), Z => n1067);
   U1402 : AO21D1 port map( A1 => a(29), A2 => a(30), B => n1066, Z => n105);
   U1403 : INVD1 port map( A => a(31), Z => n1066);

end hier_filter_none_5;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_gp_custom.all;

architecture hier_filter_none_5 of gp_custom_DW_mult_tc_8 is

   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AO21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component MUXB2DL
      port( A0, A1, SL : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component EXOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n6, n8, n14, n22, n30, n38, n42, n45, n48, n50, n53, n56, n58, 
      n61, n63, n66, n69, n71, n73, n76, n78, n79, n81, n83, n84, n86, n88, n89
      , n91, n93, n94, n96, n98, n99, n101, n103, n104, n105, n106, n155, n156,
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n178, n179, n180, n181, 
      n182, n183, n184, n185, n187, n188, n189, n190, n194, n195, n197, n199, 
      n200, n201, n202, n204, n206, n207, n208, n209, n211, n214, n215, n216, 
      n217, n219, n221, n222, n223, n224, n225, n226, n227, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n246, n248, n249, n251, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n268, n270, n271, n273, n275, 
      n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, 
      n288, n289, n293, n294, n295, n296, n297, n301, n302, n303, n305, n310, 
      n312, n313, n314, n315, n318, n319, n322, n323, n324, n326, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, 
      n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
      n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, 
      n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, 
      n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, 
      n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, 
      n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, 
      n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, 
      n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, 
      n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, 
      n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, 
      n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, 
      n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, 
      n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, 
      n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, 
      n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, 
      n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, 
      n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, 
      n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, 
      n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, 
      n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, 
      n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, 
      n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, 
      n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, 
      n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, 
      n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, 
      n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, 
      n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, 
      n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, 
      n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, 
      n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, 
      n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, 
      n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, 
      n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, 
      n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, 
      n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, 
      n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, 
      n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, 
      n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, 
      n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, 
      n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002
      , n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, 
      n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, 
      n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, 
      n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, 
      n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
      n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
      n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, 
      n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, 
      n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
      n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, 
      n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, 
      n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, 
      n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, 
      n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, 
      n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, 
      n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, 
      n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, 
      n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, 
      n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, 
      n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, 
      n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, 
      n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, 
      n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, 
      n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, 
      n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, 
      n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, 
      n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, 
      n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, 
      n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, 
      n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, 
      n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, 
      n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, 
      n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, 
      n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, 
      n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, 
      n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, 
      n1363, n1364, n1365, n1366, n1367, n1368, n1517, n1518, n1519, n1521, 
      n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, 
      n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, 
      n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, 
      n1552, n1553, n1554, n1555, n1556, n1557 : std_logic;

begin
   
   U125 : ADFULD1 port map( A => n345, B => n374, CI => n179, CO => n178, S => 
                           product(30));
   U126 : ADFULD1 port map( A => n375, B => n402, CI => n180, CO => n179, S => 
                           product(29));
   U127 : ADFULD1 port map( A => n403, B => n430, CI => n181, CO => n180, S => 
                           product(28));
   U128 : ADFULD1 port map( A => n431, B => n456, CI => n182, CO => n181, S => 
                           product(27));
   U129 : ADFULD1 port map( A => n457, B => n482, CI => n183, CO => n182, S => 
                           product(26));
   U130 : ADFULD1 port map( A => n483, B => n506, CI => n184, CO => n183, S => 
                           product(25));
   U131 : ADFULD1 port map( A => n507, B => n530, CI => n185, CO => n184, S => 
                           product(24));
   U132 : ADFULD1 port map( A => n531, B => n552, CI => n1521, CO => n185, S =>
                           product(23));
   U134 : EXOR2D1 port map( A1 => n195, A2 => n156, Z => product(22));
   U137 : OAI21D1 port map( A1 => n202, A2 => n189, B => n190, Z => n188);
   U146 : EXNOR2D1 port map( A1 => n200, A2 => n157, Z => product(21));
   U147 : AOI21D1 port map( A1 => n200, A2 => n1526, B => n197, Z => n195);
   U154 : EXNOR2D1 port map( A1 => n207, A2 => n158, Z => product(20));
   U155 : OAI21D1 port map( A1 => n214, A2 => n201, B => n202, Z => n200);
   U157 : AOI21D1 port map( A1 => n1525, A2 => n211, B => n204, Z => n202);
   U164 : EXOR2D1 port map( A1 => n214, A2 => n159, Z => product(19));
   U165 : OAI21D1 port map( A1 => n214, A2 => n208, B => n209, Z => n207);
   U174 : EXOR2D1 port map( A1 => n222, A2 => n160, Z => product(18));
   U176 : OAI21D1 port map( A1 => n233, A2 => n216, B => n217, Z => n215);
   U178 : AOI21D1 port map( A1 => n224, A2 => n1528, B => n219, Z => n217);
   U185 : EXOR2D1 port map( A1 => n227, A2 => n161, Z => product(17));
   U186 : AOI21D1 port map( A1 => n232, A2 => n223, B => n224, Z => n222);
   U188 : OAI21D1 port map( A1 => n225, A2 => n231, B => n226, Z => n224);
   U193 : EXNOR2D1 port map( A1 => n232, A2 => n162, Z => product(16));
   U194 : AOI21D1 port map( A1 => n232, A2 => n313, B => n229, Z => n227);
   U201 : EXNOR2D1 port map( A1 => n238, A2 => n163, Z => product(15));
   U203 : AOI21D1 port map( A1 => n242, A2 => n234, B => n235, Z => n233);
   U205 : OAI21D1 port map( A1 => n236, A2 => n240, B => n237, Z => n235);
   U210 : EXOR2D1 port map( A1 => n241, A2 => n164, Z => product(14));
   U211 : OAI21D1 port map( A1 => n241, A2 => n239, B => n240, Z => n238);
   U216 : EXOR2D1 port map( A1 => n249, A2 => n165, Z => product(13));
   U218 : OAI21D1 port map( A1 => n255, A2 => n243, B => n244, Z => n242);
   U220 : AOI21D1 port map( A1 => n1530, A2 => n251, B => n246, Z => n244);
   U227 : EXNOR2D1 port map( A1 => n254, A2 => n166, Z => product(12));
   U228 : AOI21D1 port map( A1 => n254, A2 => n1529, B => n251, Z => n249);
   U235 : EXNOR2D1 port map( A1 => n260, A2 => n167, Z => product(11));
   U237 : AOI21D1 port map( A1 => n256, A2 => n264, B => n257, Z => n255);
   U239 : OAI21D1 port map( A1 => n258, A2 => n262, B => n259, Z => n257);
   U244 : EXOR2D1 port map( A1 => n263, A2 => n168, Z => product(10));
   U245 : OAI21D1 port map( A1 => n263, A2 => n261, B => n262, Z => n260);
   U250 : EXOR2D1 port map( A1 => n271, A2 => n169, Z => product(9));
   U252 : OAI21D1 port map( A1 => n265, A2 => n277, B => n266, Z => n264);
   U254 : AOI21D1 port map( A1 => n1524, A2 => n273, B => n268, Z => n266);
   U261 : EXNOR2D1 port map( A1 => n276, A2 => n170, Z => product(8));
   U262 : AOI21D1 port map( A1 => n276, A2 => n1527, B => n273, Z => n271);
   U269 : EXNOR2D1 port map( A1 => n282, A2 => n171, Z => product(7));
   U271 : AOI21D1 port map( A1 => n278, A2 => n286, B => n279, Z => n277);
   U273 : OAI21D1 port map( A1 => n280, A2 => n284, B => n281, Z => n279);
   U278 : EXOR2D1 port map( A1 => n172, A2 => n285, Z => product(6));
   U279 : OAI21D1 port map( A1 => n285, A2 => n283, B => n284, Z => n282);
   U284 : EXOR2D1 port map( A1 => n173, A2 => n289, Z => product(5));
   U286 : OAI21D1 port map( A1 => n289, A2 => n287, B => n288, Z => n286);
   U291 : EXNOR2D1 port map( A1 => n174, A2 => n294, Z => product(4));
   U299 : EXOR2D1 port map( A1 => n297, A2 => n175, Z => product(3));
   U300 : OAI21D1 port map( A1 => n297, A2 => n295, B => n296, Z => n294);
   U305 : EXNOR2D1 port map( A1 => n176, A2 => n302, Z => product(2));
   U313 : EXOR2D1 port map( A1 => n303, A2 => n305, Z => product(1));
   U321 : EXOR3D1 port map( A1 => n346, A2 => n331, A3 => n330, Z => n329);
   U322 : EXOR3D1 port map( A1 => n332, A2 => n350, A3 => n348, Z => n330);
   U323 : EXOR3D1 port map( A1 => n352, A2 => n334, A3 => n333, Z => n331);
   U324 : EXOR3D1 port map( A1 => n354, A2 => n356, A3 => n335, Z => n332);
   U325 : EXOR3D1 port map( A1 => n337, A2 => n358, A3 => n336, Z => n333);
   U326 : EXOR3D1 port map( A1 => n339, A2 => n340, A3 => n360, Z => n334);
   U327 : EXOR3D1 port map( A1 => n342, A2 => n338, A3 => n341, Z => n335);
   U328 : EXOR3D1 port map( A1 => n366, A2 => n343, A3 => n362, Z => n336);
   U329 : EXOR3D1 port map( A1 => n368, A2 => n370, A3 => n364, Z => n337);
   U330 : EXOR3D1 port map( A1 => n1187, A2 => n1169, A3 => n372, Z => n338);
   U331 : EXOR3D1 port map( A1 => n1139, A2 => n1229, A3 => n1153, Z => n339);
   U332 : EXOR3D1 port map( A1 => n1103, A2 => n1117, A3 => n1109, Z => n340);
   U333 : EXOR3D1 port map( A1 => n1253, A2 => n1127, A3 => n1099, Z => n341);
   U334 : EXOR3D1 port map( A1 => n1097, A2 => n1279, A3 => n1207, Z => n342);
   U336 : ADFULD1 port map( A => n376, B => n349, CI => n347, CO => n344, S => 
                           n345);
   U337 : ADFULD1 port map( A => n351, B => n353, CI => n378, CO => n346, S => 
                           n347);
   U338 : ADFULD1 port map( A => n382, B => n355, CI => n380, CO => n348, S => 
                           n349);
   U339 : ADFULD1 port map( A => n359, B => n384, CI => n357, CO => n350, S => 
                           n351);
   U340 : ADFULD1 port map( A => n361, B => n388, CI => n386, CO => n352, S => 
                           n353);
   U341 : ADFULD1 port map( A => n365, B => n363, CI => n390, CO => n354, S => 
                           n355);
   U342 : ADFULD1 port map( A => n369, B => n371, CI => n367, CO => n356, S => 
                           n357);
   U343 : ADFULD1 port map( A => n398, B => n394, CI => n396, CO => n358, S => 
                           n359);
   U344 : ADFULD1 port map( A => n373, B => n400, CI => n392, CO => n360, S => 
                           n361);
   U345 : ADFULD1 port map( A => n1170, B => n1118, CI => n1140, CO => n362, S 
                           => n363);
   U346 : ADFULD1 port map( A => n1104, B => n1188, CI => n1110, CO => n364, S 
                           => n365);
   U347 : ADFULD1 port map( A => n1254, B => n1128, CI => n1230, CO => n366, S 
                           => n367);
   U348 : ADFULD1 port map( A => n1280, B => n1154, CI => n1208, CO => n368, S 
                           => n369);
   U349 : ADFULD1 port map( A => n1100, B => n1338, CI => n1308, CO => n370, S 
                           => n371);
   U351 : ADFULD1 port map( A => n404, B => n379, CI => n377, CO => n374, S => 
                           n375);
   U352 : ADFULD1 port map( A => n381, B => n408, CI => n406, CO => n376, S => 
                           n377);
   U353 : ADFULD1 port map( A => n410, B => n385, CI => n383, CO => n378, S => 
                           n379);
   U354 : ADFULD1 port map( A => n412, B => n389, CI => n387, CO => n380, S => 
                           n381);
   U355 : ADFULD1 port map( A => n391, B => n416, CI => n414, CO => n382, S => 
                           n383);
   U356 : ADFULD1 port map( A => n395, B => n397, CI => n399, CO => n384, S => 
                           n385);
   U357 : ADFULD1 port map( A => n418, B => n422, CI => n393, CO => n386, S => 
                           n387);
   U358 : ADFULD1 port map( A => n424, B => n426, CI => n420, CO => n388, S => 
                           n389);
   U359 : ADFULD1 port map( A => n428, B => n1189, CI => n401, CO => n390, S =>
                           n391);
   U360 : ADFULD1 port map( A => n1141, B => n1231, CI => n1171, CO => n392, S 
                           => n393);
   U361 : ADFULD1 port map( A => n1255, B => n1119, CI => n1111, CO => n394, S 
                           => n395);
   U362 : ADFULD1 port map( A => n1281, B => n1129, CI => n1105, CO => n396, S 
                           => n397);
   U363 : ADFULD1 port map( A => n1101, B => n1155, CI => n1209, CO => n398, S 
                           => n399);
   U365 : ADFULD1 port map( A => n432, B => n407, CI => n405, CO => n402, S => 
                           n403);
   U366 : ADFULD1 port map( A => n409, B => n436, CI => n434, CO => n404, S => 
                           n405);
   U367 : ADFULD1 port map( A => n438, B => n413, CI => n411, CO => n406, S => 
                           n407);
   U368 : ADFULD1 port map( A => n440, B => n417, CI => n415, CO => n408, S => 
                           n409);
   U369 : ADFULD1 port map( A => n444, B => n419, CI => n442, CO => n410, S => 
                           n411);
   U370 : ADFULD1 port map( A => n421, B => n423, CI => n425, CO => n412, S => 
                           n413);
   U371 : ADFULD1 port map( A => n448, B => n446, CI => n427, CO => n414, S => 
                           n415);
   U372 : ADFULD1 port map( A => n452, B => n429, CI => n450, CO => n416, S => 
                           n417);
   U373 : ADFULD1 port map( A => n1232, B => n1190, CI => n454, CO => n418, S 
                           => n419);
   U374 : ADFULD1 port map( A => n1142, B => n1256, CI => n1172, CO => n420, S 
                           => n421);
   U375 : ADFULD1 port map( A => n1112, B => n1130, CI => n1120, CO => n422, S 
                           => n423);
   U376 : ADFULD1 port map( A => n1282, B => n1156, CI => n1210, CO => n424, S 
                           => n425);
   U377 : ADFULD1 port map( A => n1106, B => n1340, CI => n1310, CO => n426, S 
                           => n427);
   U379 : ADFULD1 port map( A => n458, B => n435, CI => n433, CO => n430, S => 
                           n431);
   U380 : ADFULD1 port map( A => n437, B => n439, CI => n460, CO => n432, S => 
                           n433);
   U381 : ADFULD1 port map( A => n441, B => n464, CI => n462, CO => n434, S => 
                           n435);
   U382 : ADFULD1 port map( A => n466, B => n445, CI => n443, CO => n436, S => 
                           n437);
   U383 : ADFULD1 port map( A => n449, B => n451, CI => n468, CO => n438, S => 
                           n439);
   U384 : ADFULD1 port map( A => n453, B => n447, CI => n470, CO => n440, S => 
                           n441);
   U385 : ADFULD1 port map( A => n474, B => n472, CI => n476, CO => n442, S => 
                           n443);
   U386 : ADFULD1 port map( A => n455, B => n480, CI => n478, CO => n444, S => 
                           n445);
   U387 : ADFULD1 port map( A => n1131, B => n1191, CI => n1173, CO => n446, S 
                           => n447);
   U388 : ADFULD1 port map( A => n1113, B => n1233, CI => n1121, CO => n448, S 
                           => n449);
   U389 : ADFULD1 port map( A => n1283, B => n1143, CI => n1257, CO => n450, S 
                           => n451);
   U390 : ADFULD1 port map( A => n1107, B => n1157, CI => n1211, CO => n452, S 
                           => n453);
   U392 : ADFULD1 port map( A => n484, B => n461, CI => n459, CO => n456, S => 
                           n457);
   U393 : ADFULD1 port map( A => n486, B => n488, CI => n463, CO => n458, S => 
                           n459);
   U394 : ADFULD1 port map( A => n467, B => n469, CI => n465, CO => n460, S => 
                           n461);
   U395 : ADFULD1 port map( A => n492, B => n494, CI => n490, CO => n462, S => 
                           n463);
   U396 : ADFULD1 port map( A => n475, B => n477, CI => n471, CO => n464, S => 
                           n465);
   U397 : ADFULD1 port map( A => n479, B => n500, CI => n473, CO => n466, S => 
                           n467);
   U398 : ADFULD1 port map( A => n498, B => n502, CI => n496, CO => n468, S => 
                           n469);
   U399 : ADFULD1 port map( A => n504, B => n1192, CI => n481, CO => n470, S =>
                           n471);
   U400 : ADFULD1 port map( A => n1144, B => n1234, CI => n1158, CO => n472, S 
                           => n473);
   U401 : ADFULD1 port map( A => n1258, B => n1132, CI => n1122, CO => n474, S 
                           => n475);
   U402 : ADFULD1 port map( A => n1284, B => n1174, CI => n1212, CO => n476, S 
                           => n477);
   U403 : ADFULD1 port map( A => n1114, B => n1342, CI => n1312, CO => n478, S 
                           => n479);
   U405 : ADFULD1 port map( A => n508, B => n487, CI => n485, CO => n482, S => 
                           n483);
   U406 : ADFULD1 port map( A => n510, B => n512, CI => n489, CO => n484, S => 
                           n485);
   U407 : ADFULD1 port map( A => n493, B => n514, CI => n491, CO => n486, S => 
                           n487);
   U408 : ADFULD1 port map( A => n516, B => n518, CI => n495, CO => n488, S => 
                           n489);
   U409 : ADFULD1 port map( A => n501, B => n503, CI => n497, CO => n490, S => 
                           n491);
   U410 : ADFULD1 port map( A => n522, B => n524, CI => n499, CO => n492, S => 
                           n493);
   U411 : ADFULD1 port map( A => n526, B => n505, CI => n520, CO => n494, S => 
                           n495);
   U412 : ADFULD1 port map( A => n1235, B => n1259, CI => n528, CO => n496, S 
                           => n497);
   U413 : ADFULD1 port map( A => n1159, B => n1285, CI => n1193, CO => n498, S 
                           => n499);
   U414 : ADFULD1 port map( A => n1123, B => n1145, CI => n1133, CO => n500, S 
                           => n501);
   U415 : ADFULD1 port map( A => n1115, B => n1175, CI => n1213, CO => n502, S 
                           => n503);
   U417 : ADFULD1 port map( A => n532, B => n511, CI => n509, CO => n506, S => 
                           n507);
   U418 : ADFULD1 port map( A => n513, B => n536, CI => n534, CO => n508, S => 
                           n509);
   U419 : ADFULD1 port map( A => n517, B => n538, CI => n515, CO => n510, S => 
                           n511);
   U420 : ADFULD1 port map( A => n540, B => n542, CI => n519, CO => n512, S => 
                           n513);
   U421 : ADFULD1 port map( A => n525, B => n521, CI => n523, CO => n514, S => 
                           n515);
   U422 : ADFULD1 port map( A => n544, B => n546, CI => n527, CO => n516, S => 
                           n517);
   U423 : ADFULD1 port map( A => n529, B => n550, CI => n548, CO => n518, S => 
                           n519);
   U424 : ADFULD1 port map( A => n1194, B => n1260, CI => n1236, CO => n520, S 
                           => n521);
   U425 : ADFULD1 port map( A => n1134, B => n1286, CI => n1160, CO => n522, S 
                           => n523);
   U426 : ADFULD1 port map( A => n1124, B => n1176, CI => n1214, CO => n524, S 
                           => n525);
   U427 : ADFULD1 port map( A => n1146, B => n1344, CI => n1314, CO => n526, S 
                           => n527);
   U429 : ADFULD1 port map( A => n554, B => n535, CI => n533, CO => n530, S => 
                           n531);
   U430 : ADFULD1 port map( A => n556, B => n539, CI => n537, CO => n532, S => 
                           n533);
   U431 : ADFULD1 port map( A => n541, B => n560, CI => n558, CO => n534, S => 
                           n535);
   U432 : ADFULD1 port map( A => n562, B => n545, CI => n543, CO => n536, S => 
                           n537);
   U433 : ADFULD1 port map( A => n549, B => n564, CI => n547, CO => n538, S => 
                           n539);
   U434 : ADFULD1 port map( A => n566, B => n570, CI => n568, CO => n540, S => 
                           n541);
   U435 : ADFULD1 port map( A => n572, B => n1195, CI => n551, CO => n542, S =>
                           n543);
   U436 : ADFULD1 port map( A => n1135, B => n1237, CI => n1147, CO => n544, S 
                           => n545);
   U437 : ADFULD1 port map( A => n1287, B => n1161, CI => n1261, CO => n546, S 
                           => n547);
   U438 : ADFULD1 port map( A => n1125, B => n1177, CI => n1215, CO => n548, S 
                           => n549);
   U440 : ADFULD1 port map( A => n576, B => n557, CI => n555, CO => n552, S => 
                           n553);
   U441 : ADFULD1 port map( A => n559, B => n561, CI => n578, CO => n554, S => 
                           n555);
   U442 : ADFULD1 port map( A => n563, B => n582, CI => n580, CO => n556, S => 
                           n557);
   U443 : ADFULD1 port map( A => n565, B => n569, CI => n584, CO => n558, S => 
                           n559);
   U444 : ADFULD1 port map( A => n571, B => n586, CI => n567, CO => n560, S => 
                           n561);
   U445 : ADFULD1 port map( A => n590, B => n573, CI => n588, CO => n562, S => 
                           n563);
   U446 : ADFULD1 port map( A => n1196, B => n1238, CI => n592, CO => n564, S 
                           => n565);
   U447 : ADFULD1 port map( A => n1148, B => n1262, CI => n1162, CO => n566, S 
                           => n567);
   U448 : ADFULD1 port map( A => n1288, B => n1178, CI => n1216, CO => n568, S 
                           => n569);
   U449 : ADFULD1 port map( A => n1136, B => n1346, CI => n1316, CO => n570, S 
                           => n571);
   U451 : ADFULD1 port map( A => n596, B => n579, CI => n577, CO => n574, S => 
                           n575);
   U452 : ADFULD1 port map( A => n581, B => n583, CI => n598, CO => n576, S => 
                           n577);
   U453 : ADFULD1 port map( A => n585, B => n602, CI => n600, CO => n578, S => 
                           n579);
   U454 : ADFULD1 port map( A => n591, B => n589, CI => n604, CO => n580, S => 
                           n581);
   U455 : ADFULD1 port map( A => n606, B => n608, CI => n587, CO => n582, S => 
                           n583);
   U456 : ADFULD1 port map( A => n593, B => n612, CI => n610, CO => n584, S => 
                           n585);
   U457 : ADFULD1 port map( A => n1197, B => n1263, CI => n1239, CO => n586, S 
                           => n587);
   U458 : ADFULD1 port map( A => n1289, B => n1163, CI => n1149, CO => n588, S 
                           => n589);
   U459 : ADFULD1 port map( A => n1137, B => n1179, CI => n1217, CO => n590, S 
                           => n591);
   U461 : ADFULD1 port map( A => n616, B => n599, CI => n597, CO => n594, S => 
                           n595);
   U462 : ADFULD1 port map( A => n601, B => n603, CI => n618, CO => n596, S => 
                           n597);
   U463 : ADFULD1 port map( A => n622, B => n605, CI => n620, CO => n598, S => 
                           n599);
   U464 : ADFULD1 port map( A => n609, B => n611, CI => n607, CO => n600, S => 
                           n601);
   U465 : ADFULD1 port map( A => n626, B => n628, CI => n624, CO => n602, S => 
                           n603);
   U466 : ADFULD1 port map( A => n630, B => n1240, CI => n613, CO => n604, S =>
                           n605);
   U467 : ADFULD1 port map( A => n1150, B => n1264, CI => n1180, CO => n606, S 
                           => n607);
   U468 : ADFULD1 port map( A => n1290, B => n1198, CI => n1218, CO => n608, S 
                           => n609);
   U469 : ADFULD1 port map( A => n1164, B => n1348, CI => n1318, CO => n610, S 
                           => n611);
   U471 : ADFULD1 port map( A => n634, B => n619, CI => n617, CO => n614, S => 
                           n615);
   U472 : ADFULD1 port map( A => n621, B => n623, CI => n636, CO => n616, S => 
                           n617);
   U473 : ADFULD1 port map( A => n640, B => n625, CI => n638, CO => n618, S => 
                           n619);
   U474 : ADFULD1 port map( A => n627, B => n644, CI => n629, CO => n620, S => 
                           n621);
   U475 : ADFULD1 port map( A => n646, B => n631, CI => n642, CO => n622, S => 
                           n623);
   U476 : ADFULD1 port map( A => n1241, B => n1265, CI => n648, CO => n624, S 
                           => n625);
   U477 : ADFULD1 port map( A => n1291, B => n1181, CI => n1165, CO => n626, S 
                           => n627);
   U478 : ADFULD1 port map( A => n1151, B => n1199, CI => n1219, CO => n628, S 
                           => n629);
   U480 : ADFULD1 port map( A => n652, B => n637, CI => n635, CO => n632, S => 
                           n633);
   U481 : ADFULD1 port map( A => n639, B => n641, CI => n654, CO => n634, S => 
                           n635);
   U482 : ADFULD1 port map( A => n658, B => n645, CI => n656, CO => n636, S => 
                           n637);
   U483 : ADFULD1 port map( A => n647, B => n660, CI => n643, CO => n638, S => 
                           n639);
   U484 : ADFULD1 port map( A => n649, B => n664, CI => n662, CO => n640, S => 
                           n641);
   U485 : ADFULD1 port map( A => n1182, B => n1292, CI => n1242, CO => n642, S 
                           => n643);
   U486 : ADFULD1 port map( A => n1166, B => n1266, CI => n1220, CO => n644, S 
                           => n645);
   U487 : ADFULD1 port map( A => n1200, B => n1350, CI => n1320, CO => n646, S 
                           => n647);
   U489 : ADFULD1 port map( A => n668, B => n655, CI => n653, CO => n650, S => 
                           n651);
   U490 : ADFULD1 port map( A => n670, B => n659, CI => n657, CO => n652, S => 
                           n653);
   U491 : ADFULD1 port map( A => n663, B => n661, CI => n672, CO => n654, S => 
                           n655);
   U492 : ADFULD1 port map( A => n676, B => n678, CI => n674, CO => n656, S => 
                           n657);
   U493 : ADFULD1 port map( A => n680, B => n1293, CI => n665, CO => n658, S =>
                           n659);
   U494 : ADFULD1 port map( A => n1243, B => n1183, CI => n1267, CO => n660, S 
                           => n661);
   U495 : ADFULD1 port map( A => n1167, B => n1201, CI => n1221, CO => n662, S 
                           => n663);
   U497 : ADFULD1 port map( A => n684, B => n671, CI => n669, CO => n666, S => 
                           n667);
   U498 : ADFULD1 port map( A => n686, B => n688, CI => n673, CO => n668, S => 
                           n669);
   U499 : ADFULD1 port map( A => n677, B => n679, CI => n675, CO => n670, S => 
                           n671);
   U500 : ADFULD1 port map( A => n692, B => n681, CI => n690, CO => n672, S => 
                           n673);
   U501 : ADFULD1 port map( A => n1244, B => n1294, CI => n694, CO => n674, S 
                           => n675);
   U502 : ADFULD1 port map( A => n1184, B => n1268, CI => n1222, CO => n676, S 
                           => n677);
   U503 : ADFULD1 port map( A => n1202, B => n1352, CI => n1322, CO => n678, S 
                           => n679);
   U505 : ADFULD1 port map( A => n698, B => n687, CI => n685, CO => n682, S => 
                           n683);
   U506 : ADFULD1 port map( A => n700, B => n702, CI => n689, CO => n684, S => 
                           n685);
   U507 : ADFULD1 port map( A => n691, B => n704, CI => n693, CO => n686, S => 
                           n687);
   U508 : ADFULD1 port map( A => n695, B => n708, CI => n706, CO => n688, S => 
                           n689);
   U509 : ADFULD1 port map( A => n1203, B => n1295, CI => n1245, CO => n690, S 
                           => n691);
   U510 : ADFULD1 port map( A => n1185, B => n1269, CI => n1223, CO => n692, S 
                           => n693);
   U512 : ADFULD1 port map( A => n712, B => n701, CI => n699, CO => n696, S => 
                           n697);
   U513 : ADFULD1 port map( A => n703, B => n705, CI => n714, CO => n698, S => 
                           n699);
   U514 : ADFULD1 port map( A => n716, B => n718, CI => n707, CO => n700, S => 
                           n701);
   U515 : ADFULD1 port map( A => n720, B => n1270, CI => n709, CO => n702, S =>
                           n703);
   U516 : ADFULD1 port map( A => n1246, B => n1296, CI => n1224, CO => n704, S 
                           => n705);
   U517 : ADFULD1 port map( A => n1204, B => n1354, CI => n1324, CO => n706, S 
                           => n707);
   U519 : ADFULD1 port map( A => n724, B => n715, CI => n713, CO => n710, S => 
                           n711);
   U520 : ADFULD1 port map( A => n717, B => n719, CI => n726, CO => n712, S => 
                           n713);
   U521 : ADFULD1 port map( A => n730, B => n721, CI => n728, CO => n714, S => 
                           n715);
   U522 : ADFULD1 port map( A => n1247, B => n1271, CI => n732, CO => n716, S 
                           => n717);
   U523 : ADFULD1 port map( A => n1205, B => n1297, CI => n1225, CO => n718, S 
                           => n719);
   U525 : ADFULD1 port map( A => n736, B => n727, CI => n725, CO => n722, S => 
                           n723);
   U526 : ADFULD1 port map( A => n729, B => n731, CI => n738, CO => n724, S => 
                           n725);
   U527 : ADFULD1 port map( A => n733, B => n742, CI => n740, CO => n726, S => 
                           n727);
   U528 : ADFULD1 port map( A => n1272, B => n1298, CI => n1226, CO => n728, S 
                           => n729);
   U529 : ADFULD1 port map( A => n1248, B => n1356, CI => n1326, CO => n730, S 
                           => n731);
   U531 : ADFULD1 port map( A => n746, B => n739, CI => n737, CO => n734, S => 
                           n735);
   U532 : ADFULD1 port map( A => n748, B => n750, CI => n741, CO => n736, S => 
                           n737);
   U533 : ADFULD1 port map( A => n752, B => n1299, CI => n743, CO => n738, S =>
                           n739);
   U534 : ADFULD1 port map( A => n1273, B => n1249, CI => n1227, CO => n740, S 
                           => n741);
   U536 : ADFULD1 port map( A => n756, B => n749, CI => n747, CO => n744, S => 
                           n745);
   U537 : ADFULD1 port map( A => n758, B => n753, CI => n751, CO => n746, S => 
                           n747);
   U538 : ADFULD1 port map( A => n1274, B => n1300, CI => n760, CO => n748, S 
                           => n749);
   U539 : ADFULD1 port map( A => n1250, B => n1358, CI => n1328, CO => n750, S 
                           => n751);
   U541 : ADFULD1 port map( A => n764, B => n759, CI => n757, CO => n754, S => 
                           n755);
   U542 : ADFULD1 port map( A => n761, B => n768, CI => n766, CO => n756, S => 
                           n757);
   U543 : ADFULD1 port map( A => n1275, B => n1301, CI => n1251, CO => n758, S 
                           => n759);
   U545 : ADFULD1 port map( A => n767, B => n772, CI => n765, CO => n762, S => 
                           n763);
   U546 : ADFULD1 port map( A => n774, B => n1302, CI => n769, CO => n764, S =>
                           n765);
   U547 : ADFULD1 port map( A => n1276, B => n1360, CI => n1330, CO => n766, S 
                           => n767);
   U549 : ADFULD1 port map( A => n778, B => n775, CI => n773, CO => n770, S => 
                           n771);
   U550 : ADFULD1 port map( A => n1277, B => n1303, CI => n780, CO => n772, S 
                           => n773);
   U552 : ADFULD1 port map( A => n781, B => n784, CI => n779, CO => n776, S => 
                           n777);
   U553 : ADFULD1 port map( A => n1304, B => n1362, CI => n1332, CO => n778, S 
                           => n779);
   U555 : ADFULD1 port map( A => n788, B => n1305, CI => n785, CO => n782, S =>
                           n783);
   U557 : ADFULD1 port map( A => n1334, B => n1364, CI => n790, CO => n786, S 
                           => n787);
   U561 : NOR2M1D1 port map( A1 => n104, A2 => n105, Z => n1081);
   U562 : MUXB2DL port map( A0 => n104, A1 => n105, SL => n794, Z => n1097);
   U563 : MUXB2DL port map( A0 => b(1), A1 => n1556, SL => n106, Z => n794);
   U564 : MUXB2DL port map( A0 => n104, A1 => n105, SL => n795, Z => n1098);
   U565 : NAN2M1D1 port map( A1 => n106, A2 => b(0), Z => n795);
   U566 : NOR2M1D1 port map( A1 => n99, A2 => n101, Z => n1082);
   U567 : MUXB2DL port map( A0 => n99, A1 => n101, SL => n796, Z => n1099);
   U568 : MUXB2DL port map( A0 => b(3), A1 => n1554, SL => n103, Z => n796);
   U569 : MUXB2DL port map( A0 => n99, A1 => n101, SL => n797, Z => n1100);
   U570 : MUXB2DL port map( A0 => n1553, A1 => b(1), SL => n103, Z => n797);
   U571 : MUXB2DL port map( A0 => n99, A1 => n101, SL => n798, Z => n1101);
   U572 : MUXB2DL port map( A0 => b(1), A1 => n1556, SL => n103, Z => n798);
   U573 : MUXB2DL port map( A0 => n99, A1 => n101, SL => n799, Z => n1102);
   U574 : NAN2M1D1 port map( A1 => n103, A2 => b(0), Z => n799);
   U575 : NOR2M1D1 port map( A1 => n94, A2 => n96, Z => n1083);
   U576 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n800, Z => n1103);
   U577 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n98, Z => n800);
   U578 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n801, Z => n1104);
   U579 : MUXB2DL port map( A0 => n1549, A1 => n1551, SL => n98, Z => n801);
   U580 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n802, Z => n1105);
   U581 : MUXB2DL port map( A0 => b(3), A1 => n1554, SL => n98, Z => n802);
   U582 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n803, Z => n1106);
   U583 : MUXB2DL port map( A0 => n1553, A1 => b(1), SL => n98, Z => n803);
   U584 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n804, Z => n1107);
   U585 : MUXB2DL port map( A0 => b(1), A1 => n1556, SL => n98, Z => n804);
   U586 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n805, Z => n1108);
   U587 : NAN2M1D1 port map( A1 => n98, A2 => b(0), Z => n805);
   U588 : NOR2M1D1 port map( A1 => n89, A2 => n91, Z => n1084);
   U589 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n806, Z => n1109);
   U590 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n93, Z => n806);
   U591 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n807, Z => n1110);
   U592 : MUXB2DL port map( A0 => b(6), A1 => n1547, SL => n93, Z => n807);
   U593 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n808, Z => n1111);
   U594 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n93, Z => n808);
   U595 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n809, Z => n1112);
   U596 : MUXB2DL port map( A0 => n1549, A1 => n1551, SL => n93, Z => n809);
   U597 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n810, Z => n1113);
   U598 : MUXB2DL port map( A0 => b(3), A1 => n1554, SL => n93, Z => n810);
   U599 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n811, Z => n1114);
   U600 : MUXB2DL port map( A0 => n1553, A1 => b(1), SL => n93, Z => n811);
   U601 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n812, Z => n1115);
   U602 : MUXB2DL port map( A0 => b(1), A1 => n1556, SL => n93, Z => n812);
   U603 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n813, Z => n1116);
   U604 : NAN2M1D1 port map( A1 => n93, A2 => n1556, Z => n813);
   U605 : NOR2M1D1 port map( A1 => n84, A2 => n86, Z => n1085);
   U606 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n814, Z => n1117);
   U607 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n88, Z => n814);
   U608 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n815, Z => n1118);
   U609 : MUXB2DL port map( A0 => n1545, A1 => b(7), SL => n88, Z => n815);
   U610 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n816, Z => n1119);
   U611 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n88, Z => n816);
   U612 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n817, Z => n1120);
   U613 : MUXB2DL port map( A0 => b(6), A1 => n1547, SL => n88, Z => n817);
   U614 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n818, Z => n1121);
   U615 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n88, Z => n818);
   U616 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n819, Z => n1122);
   U617 : MUXB2DL port map( A0 => n1549, A1 => n1551, SL => n88, Z => n819);
   U618 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n820, Z => n1123);
   U619 : MUXB2DL port map( A0 => b(3), A1 => n1554, SL => n88, Z => n820);
   U620 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n821, Z => n1124);
   U621 : MUXB2DL port map( A0 => n1553, A1 => b(1), SL => n88, Z => n821);
   U622 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n822, Z => n1125);
   U623 : MUXB2DL port map( A0 => b(1), A1 => n1556, SL => n88, Z => n822);
   U624 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n823, Z => n1126);
   U625 : NAN2M1D1 port map( A1 => n88, A2 => n1556, Z => n823);
   U626 : NOR2M1D1 port map( A1 => n79, A2 => n81, Z => n1086);
   U627 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n824, Z => n1127);
   U628 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n83, Z => n824);
   U629 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n825, Z => n1128);
   U630 : MUXB2DL port map( A0 => n1543, A1 => b(9), SL => n83, Z => n825);
   U631 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n826, Z => n1129);
   U632 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n83, Z => n826);
   U633 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n827, Z => n1130);
   U634 : MUXB2DL port map( A0 => n1545, A1 => b(7), SL => n83, Z => n827);
   U635 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n828, Z => n1131);
   U636 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n83, Z => n828);
   U637 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n829, Z => n1132);
   U638 : MUXB2DL port map( A0 => b(6), A1 => n1547, SL => n83, Z => n829);
   U639 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n830, Z => n1133);
   U640 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n83, Z => n830);
   U641 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n831, Z => n1134);
   U642 : MUXB2DL port map( A0 => n1549, A1 => n1551, SL => n83, Z => n831);
   U643 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n832, Z => n1135);
   U644 : MUXB2DL port map( A0 => n1551, A1 => n1554, SL => n83, Z => n832);
   U645 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n833, Z => n1136);
   U646 : MUXB2DL port map( A0 => n1554, A1 => b(1), SL => n83, Z => n833);
   U647 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n834, Z => n1137);
   U648 : MUXB2DL port map( A0 => b(1), A1 => n1556, SL => n83, Z => n834);
   U649 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n835, Z => n1138);
   U650 : NAN2M1D1 port map( A1 => n83, A2 => b(0), Z => n835);
   U651 : NOR2M1D1 port map( A1 => n73, A2 => n76, Z => n1087);
   U652 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n836, Z => n1139);
   U653 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n78, Z => n836);
   U654 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n837, Z => n1140);
   U655 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n78, Z => n837);
   U656 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n838, Z => n1141);
   U657 : MUXB2DL port map( A0 => b(11), A1 => n1543, SL => n78, Z => n838);
   U658 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n839, Z => n1142);
   U659 : MUXB2DL port map( A0 => n1543, A1 => b(9), SL => n78, Z => n839);
   U660 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n840, Z => n1143);
   U661 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n78, Z => n840);
   U662 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n841, Z => n1144);
   U663 : MUXB2DL port map( A0 => n1545, A1 => b(7), SL => n78, Z => n841);
   U664 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n842, Z => n1145);
   U665 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n78, Z => n842);
   U666 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n843, Z => n1146);
   U667 : MUXB2DL port map( A0 => b(6), A1 => n1547, SL => n78, Z => n843);
   U668 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n844, Z => n1147);
   U669 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n78, Z => n844);
   U670 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n845, Z => n1148);
   U671 : MUXB2DL port map( A0 => n1549, A1 => n1551, SL => n78, Z => n845);
   U672 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n846, Z => n1149);
   U673 : MUXB2DL port map( A0 => n1551, A1 => n1554, SL => n78, Z => n846);
   U674 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n847, Z => n1150);
   U675 : MUXB2DL port map( A0 => n1554, A1 => b(1), SL => n78, Z => n847);
   U676 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n848, Z => n1151);
   U677 : MUXB2DL port map( A0 => b(1), A1 => n1556, SL => n78, Z => n848);
   U678 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n849, Z => n1152);
   U679 : NAN2M1D1 port map( A1 => n78, A2 => n1556, Z => n849);
   U680 : NOR2M1D1 port map( A1 => n66, A2 => n69, Z => n1088);
   U681 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n850, Z => n1153);
   U682 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n71, Z => n850);
   U683 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n851, Z => n1154);
   U684 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n71, Z => n851);
   U685 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n852, Z => n1155);
   U686 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n71, Z => n852);
   U687 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n853, Z => n1156);
   U688 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n71, Z => n853);
   U689 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n854, Z => n1157);
   U690 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n71, Z => n854);
   U691 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n855, Z => n1158);
   U692 : MUXB2DL port map( A0 => n1543, A1 => b(9), SL => n71, Z => n855);
   U693 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n856, Z => n1159);
   U694 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n71, Z => n856);
   U695 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n857, Z => n1160);
   U696 : MUXB2DL port map( A0 => n1545, A1 => b(7), SL => n71, Z => n857);
   U697 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n858, Z => n1161);
   U698 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n71, Z => n858);
   U699 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n859, Z => n1162);
   U700 : MUXB2DL port map( A0 => b(6), A1 => n1547, SL => n71, Z => n859);
   U701 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n860, Z => n1163);
   U702 : MUXB2DL port map( A0 => n1547, A1 => n1549, SL => n71, Z => n860);
   U703 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n861, Z => n1164);
   U704 : MUXB2DL port map( A0 => b(4), A1 => n1551, SL => n71, Z => n861);
   U705 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n862, Z => n1165);
   U706 : MUXB2DL port map( A0 => n1551, A1 => n1554, SL => n71, Z => n862);
   U707 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n863, Z => n1166);
   U708 : MUXB2DL port map( A0 => n1553, A1 => b(1), SL => n71, Z => n863);
   U709 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n864, Z => n1167);
   U710 : MUXB2DL port map( A0 => b(1), A1 => n1556, SL => n71, Z => n864);
   U711 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n865, Z => n1168);
   U712 : NAN2M1D1 port map( A1 => n71, A2 => n1556, Z => n865);
   U713 : NOR2M1D1 port map( A1 => n58, A2 => n61, Z => n1089);
   U714 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n866, Z => n1169);
   U715 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n63, Z => n866);
   U716 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n867, Z => n1170);
   U717 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n63, Z => n867);
   U718 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n868, Z => n1171);
   U719 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n63, Z => n868);
   U720 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n869, Z => n1172);
   U721 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n63, Z => n869);
   U722 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n870, Z => n1173);
   U723 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n63, Z => n870);
   U724 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n871, Z => n1174);
   U725 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n63, Z => n871);
   U726 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n872, Z => n1175);
   U727 : MUXB2DL port map( A0 => b(11), A1 => n1543, SL => n63, Z => n872);
   U728 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n873, Z => n1176);
   U729 : MUXB2DL port map( A0 => n1543, A1 => b(9), SL => n63, Z => n873);
   U730 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n874, Z => n1177);
   U731 : MUXB2DL port map( A0 => b(9), A1 => n1545, SL => n63, Z => n874);
   U732 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n875, Z => n1178);
   U733 : MUXB2DL port map( A0 => n1545, A1 => b(7), SL => n63, Z => n875);
   U734 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n876, Z => n1179);
   U735 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n63, Z => n876);
   U736 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n877, Z => n1180);
   U737 : MUXB2DL port map( A0 => b(6), A1 => n1547, SL => n63, Z => n877);
   U738 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n878, Z => n1181);
   U739 : MUXB2DL port map( A0 => n1547, A1 => b(4), SL => n63, Z => n878);
   U740 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n879, Z => n1182);
   U741 : MUXB2DL port map( A0 => n1549, A1 => n1551, SL => n63, Z => n879);
   U742 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n880, Z => n1183);
   U743 : MUXB2DL port map( A0 => b(3), A1 => n1554, SL => n63, Z => n880);
   U744 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n881, Z => n1184);
   U745 : MUXB2DL port map( A0 => n1553, A1 => b(1), SL => n63, Z => n881);
   U746 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n882, Z => n1185);
   U747 : MUXB2DL port map( A0 => b(1), A1 => n1556, SL => n63, Z => n882);
   U748 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n883, Z => n1186);
   U749 : NAN2M1D1 port map( A1 => n63, A2 => b(0), Z => n883);
   U750 : NOR2M1D1 port map( A1 => n50, A2 => n53, Z => n1090);
   U751 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n884, Z => n1187);
   U752 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n56, Z => n884);
   U753 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n885, Z => n1188);
   U754 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n56, Z => n885);
   U755 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n886, Z => n1189);
   U756 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n56, Z => n886);
   U757 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n887, Z => n1190);
   U758 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n56, Z => n887);
   U759 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n888, Z => n1191);
   U760 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n56, Z => n888);
   U761 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n889, Z => n1192);
   U762 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n56, Z => n889);
   U763 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n890, Z => n1193);
   U764 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n56, Z => n890);
   U765 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n891, Z => n1194);
   U766 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n56, Z => n891);
   U767 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n892, Z => n1195);
   U768 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n56, Z => n892);
   U769 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n893, Z => n1196);
   U770 : MUXB2DL port map( A0 => n1543, A1 => b(9), SL => n56, Z => n893);
   U771 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n894, Z => n1197);
   U772 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n56, Z => n894);
   U773 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n895, Z => n1198);
   U774 : MUXB2DL port map( A0 => n1545, A1 => b(7), SL => n56, Z => n895);
   U775 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n896, Z => n1199);
   U776 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n56, Z => n896);
   U777 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n897, Z => n1200);
   U778 : MUXB2DL port map( A0 => b(6), A1 => n1547, SL => n56, Z => n897);
   U779 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n898, Z => n1201);
   U780 : MUXB2DL port map( A0 => b(5), A1 => n1549, SL => n56, Z => n898);
   U781 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n899, Z => n1202);
   U782 : MUXB2DL port map( A0 => n1549, A1 => n1551, SL => n56, Z => n899);
   U783 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n900, Z => n1203);
   U784 : MUXB2DL port map( A0 => n1551, A1 => n1553, SL => n56, Z => n900);
   U785 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n901, Z => n1204);
   U786 : MUXB2DL port map( A0 => n1553, A1 => b(1), SL => n56, Z => n901);
   U787 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n902, Z => n1205);
   U788 : MUXB2DL port map( A0 => b(1), A1 => b(0), SL => n56, Z => n902);
   U789 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n903, Z => n1206);
   U790 : NAN2M1D1 port map( A1 => n56, A2 => n1556, Z => n903);
   U791 : NOR2M1D1 port map( A1 => n42, A2 => n45, Z => n1091);
   U792 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n904, Z => n1207);
   U793 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n48, Z => n904);
   U794 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n905, Z => n1208);
   U795 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n48, Z => n905);
   U796 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n906, Z => n1209);
   U797 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n48, Z => n906);
   U798 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n907, Z => n1210);
   U799 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n48, Z => n907);
   U800 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n908, Z => n1211);
   U801 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n48, Z => n908);
   U802 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n909, Z => n1212);
   U803 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n48, Z => n909);
   U804 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n910, Z => n1213);
   U805 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n48, Z => n910);
   U806 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n911, Z => n1214);
   U807 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n48, Z => n911);
   U808 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n912, Z => n1215);
   U809 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n48, Z => n912);
   U810 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n913, Z => n1216);
   U811 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n48, Z => n913);
   U812 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n914, Z => n1217);
   U813 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n48, Z => n914);
   U814 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n915, Z => n1218);
   U815 : MUXB2DL port map( A0 => n1543, A1 => b(9), SL => n48, Z => n915);
   U816 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n916, Z => n1219);
   U817 : MUXB2DL port map( A0 => b(9), A1 => n1545, SL => n48, Z => n916);
   U818 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n917, Z => n1220);
   U819 : MUXB2DL port map( A0 => n1545, A1 => b(7), SL => n48, Z => n917);
   U820 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n918, Z => n1221);
   U821 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n48, Z => n918);
   U822 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n919, Z => n1222);
   U823 : MUXB2DL port map( A0 => b(6), A1 => n1547, SL => n48, Z => n919);
   U824 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n920, Z => n1223);
   U825 : MUXB2DL port map( A0 => b(5), A1 => n1549, SL => n48, Z => n920);
   U826 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n921, Z => n1224);
   U827 : MUXB2DL port map( A0 => n1549, A1 => b(3), SL => n48, Z => n921);
   U828 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n922, Z => n1225);
   U829 : MUXB2DL port map( A0 => b(3), A1 => n1554, SL => n48, Z => n922);
   U830 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n923, Z => n1226);
   U831 : MUXB2DL port map( A0 => n1553, A1 => b(1), SL => n48, Z => n923);
   U832 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n924, Z => n1227);
   U833 : MUXB2DL port map( A0 => b(1), A1 => b(0), SL => n48, Z => n924);
   U834 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n925, Z => n1228);
   U835 : NAN2M1D1 port map( A1 => n48, A2 => b(0), Z => n925);
   U836 : NOR2M1D1 port map( A1 => n1519, A2 => n38, Z => n1092);
   U837 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n926, Z => n1229);
   U838 : MUXB2DL port map( A0 => b(23), A1 => b(22), SL => n1538, Z => n926);
   U839 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n927, Z => n1230);
   U840 : MUXB2DL port map( A0 => b(22), A1 => b(21), SL => n1538, Z => n927);
   U841 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n928, Z => n1231);
   U842 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n1538, Z => n928);
   U843 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n929, Z => n1232);
   U844 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n1538, Z => n929);
   U845 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n930, Z => n1233);
   U846 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n1538, Z => n930);
   U847 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n931, Z => n1234);
   U848 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n1538, Z => n931);
   U849 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n932, Z => n1235);
   U850 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n1538, Z => n932);
   U851 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n933, Z => n1236);
   U852 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n1538, Z => n933);
   U853 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n934, Z => n1237);
   U854 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n1538, Z => n934);
   U855 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n935, Z => n1238);
   U856 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n1538, Z => n935);
   U857 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n936, Z => n1239);
   U858 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n1538, Z => n936);
   U859 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n937, Z => n1240);
   U860 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n1538, Z => n937);
   U861 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n938, Z => n1241);
   U862 : MUXB2DL port map( A0 => b(11), A1 => n1543, SL => n1538, Z => n938);
   U863 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n939, Z => n1242);
   U864 : MUXB2DL port map( A0 => n1543, A1 => b(9), SL => n1538, Z => n939);
   U865 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n940, Z => n1243);
   U866 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n1538, Z => n940);
   U867 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n941, Z => n1244);
   U868 : MUXB2DL port map( A0 => n1545, A1 => b(7), SL => n1538, Z => n941);
   U869 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n942, Z => n1245);
   U870 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n1538, Z => n942);
   U871 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n943, Z => n1246);
   U872 : MUXB2DL port map( A0 => b(6), A1 => n1547, SL => n1538, Z => n943);
   U873 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n944, Z => n1247);
   U874 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n1538, Z => n944);
   U875 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n945, Z => n1248);
   U876 : MUXB2DL port map( A0 => n1549, A1 => b(3), SL => n1538, Z => n945);
   U877 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n946, Z => n1249);
   U878 : MUXB2DL port map( A0 => b(3), A1 => n1553, SL => n1538, Z => n946);
   U879 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n947, Z => n1250);
   U880 : MUXB2DL port map( A0 => n1553, A1 => b(1), SL => n1538, Z => n947);
   U881 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n948, Z => n1251);
   U882 : MUXB2DL port map( A0 => b(1), A1 => b(0), SL => n1538, Z => n948);
   U883 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n949, Z => n1252);
   U884 : NAN2M1D1 port map( A1 => n1538, A2 => b(0), Z => n949);
   U886 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n950, Z => n1253);
   U887 : MUXB2DL port map( A0 => b(25), A1 => b(24), SL => n1539, Z => n950);
   U888 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n951, Z => n1254);
   U889 : MUXB2DL port map( A0 => b(24), A1 => b(23), SL => n1539, Z => n951);
   U890 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n952, Z => n1255);
   U891 : MUXB2DL port map( A0 => b(23), A1 => b(22), SL => n1539, Z => n952);
   U892 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n953, Z => n1256);
   U893 : MUXB2DL port map( A0 => b(22), A1 => b(21), SL => n1539, Z => n953);
   U894 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n954, Z => n1257);
   U895 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n1539, Z => n954);
   U896 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n955, Z => n1258);
   U897 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n1539, Z => n955);
   U898 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n956, Z => n1259);
   U899 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n1539, Z => n956);
   U900 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n957, Z => n1260);
   U901 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n1539, Z => n957);
   U902 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n958, Z => n1261);
   U903 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n1539, Z => n958);
   U904 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n959, Z => n1262);
   U905 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n1539, Z => n959);
   U906 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n960, Z => n1263);
   U907 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n1539, Z => n960);
   U908 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n961, Z => n1264);
   U909 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n1539, Z => n961);
   U910 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n962, Z => n1265);
   U911 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n1539, Z => n962);
   U912 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n963, Z => n1266);
   U913 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n1539, Z => n963);
   U914 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n964, Z => n1267);
   U915 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n1539, Z => n964);
   U916 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n965, Z => n1268);
   U917 : MUXB2DL port map( A0 => n1543, A1 => b(9), SL => n1539, Z => n965);
   U918 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n966, Z => n1269);
   U919 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n1539, Z => n966);
   U920 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n967, Z => n1270);
   U921 : MUXB2DL port map( A0 => n1545, A1 => b(7), SL => n1539, Z => n967);
   U922 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n968, Z => n1271);
   U923 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n1539, Z => n968);
   U924 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n969, Z => n1272);
   U925 : MUXB2DL port map( A0 => b(6), A1 => n1547, SL => n1539, Z => n969);
   U926 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n970, Z => n1273);
   U927 : MUXB2DL port map( A0 => b(5), A1 => n1549, SL => n1539, Z => n970);
   U928 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n971, Z => n1274);
   U929 : MUXB2DL port map( A0 => n1549, A1 => b(3), SL => n1539, Z => n971);
   U930 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n972, Z => n1275);
   U931 : MUXB2DL port map( A0 => b(3), A1 => n1553, SL => n1539, Z => n972);
   U932 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n973, Z => n1276);
   U933 : MUXB2DL port map( A0 => n1553, A1 => b(1), SL => n1539, Z => n973);
   U934 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n974, Z => n1277);
   U935 : MUXB2DL port map( A0 => b(1), A1 => b(0), SL => n1539, Z => n974);
   U936 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n975, Z => n1278);
   U937 : NAN2M1D1 port map( A1 => n1539, A2 => b(0), Z => n975);
   U938 : NOR2M1D1 port map( A1 => n1518, A2 => n22, Z => n1094);
   U939 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n976, Z => n1279);
   U940 : MUXB2DL port map( A0 => b(27), A1 => b(26), SL => n1541, Z => n976);
   U941 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n977, Z => n1280);
   U942 : MUXB2DL port map( A0 => b(26), A1 => b(25), SL => n1541, Z => n977);
   U943 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n978, Z => n1281);
   U944 : MUXB2DL port map( A0 => b(25), A1 => b(24), SL => n1541, Z => n978);
   U945 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n979, Z => n1282);
   U946 : MUXB2DL port map( A0 => b(24), A1 => b(23), SL => n1541, Z => n979);
   U947 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n980, Z => n1283);
   U948 : MUXB2DL port map( A0 => b(23), A1 => b(22), SL => n1541, Z => n980);
   U949 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n981, Z => n1284);
   U950 : MUXB2DL port map( A0 => b(22), A1 => b(21), SL => n1541, Z => n981);
   U951 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n982, Z => n1285);
   U952 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n1541, Z => n982);
   U953 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n983, Z => n1286);
   U954 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n1541, Z => n983);
   U955 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n984, Z => n1287);
   U956 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n1541, Z => n984);
   U957 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n985, Z => n1288);
   U958 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n1541, Z => n985);
   U959 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n986, Z => n1289);
   U960 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n1541, Z => n986);
   U961 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n987, Z => n1290);
   U962 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n1541, Z => n987);
   U963 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n988, Z => n1291);
   U964 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n1541, Z => n988);
   U965 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n989, Z => n1292);
   U966 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n1541, Z => n989);
   U967 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n990, Z => n1293);
   U968 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n1541, Z => n990);
   U969 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n991, Z => n1294);
   U970 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n1541, Z => n991);
   U971 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n992, Z => n1295);
   U972 : MUXB2DL port map( A0 => b(11), A1 => n1543, SL => n1541, Z => n992);
   U973 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n993, Z => n1296);
   U974 : MUXB2DL port map( A0 => n1543, A1 => b(9), SL => n1541, Z => n993);
   U975 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n994, Z => n1297);
   U976 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n1541, Z => n994);
   U977 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n995, Z => n1298);
   U978 : MUXB2DL port map( A0 => n1545, A1 => b(7), SL => n1541, Z => n995);
   U979 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n996, Z => n1299);
   U980 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n1541, Z => n996);
   U981 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n997, Z => n1300);
   U982 : MUXB2DL port map( A0 => b(6), A1 => n1547, SL => n1541, Z => n997);
   U983 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n998, Z => n1301);
   U984 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n1541, Z => n998);
   U985 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n999, Z => n1302);
   U986 : MUXB2DL port map( A0 => n1549, A1 => n1551, SL => n1541, Z => n999);
   U987 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n1000, Z => n1303);
   U988 : MUXB2DL port map( A0 => b(3), A1 => n1554, SL => n1541, Z => n1000);
   U989 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n1001, Z => n1304);
   U990 : MUXB2DL port map( A0 => n1553, A1 => b(1), SL => n1541, Z => n1001);
   U991 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n1002, Z => n1305);
   U992 : MUXB2DL port map( A0 => b(1), A1 => n1556, SL => n1541, Z => n1002);
   U993 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n1003, Z => n1306);
   U994 : NAN2M1D1 port map( A1 => n1541, A2 => b(0), Z => n1003);
   U995 : NOR2M1D1 port map( A1 => n1517, A2 => n14, Z => n1095);
   U996 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1004, Z => n1307);
   U997 : MUXB2DL port map( A0 => b(29), A1 => b(28), SL => n1542, Z => n1004);
   U998 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1005, Z => n1308);
   U999 : MUXB2DL port map( A0 => b(28), A1 => b(27), SL => n1542, Z => n1005);
   U1000 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1006, Z => n1309);
   U1001 : MUXB2DL port map( A0 => b(27), A1 => b(26), SL => n1542, Z => n1006)
                           ;
   U1002 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1007, Z => n1310);
   U1003 : MUXB2DL port map( A0 => b(26), A1 => b(25), SL => n1542, Z => n1007)
                           ;
   U1004 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1008, Z => n1311);
   U1005 : MUXB2DL port map( A0 => b(25), A1 => b(24), SL => n1542, Z => n1008)
                           ;
   U1006 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1009, Z => n1312);
   U1007 : MUXB2DL port map( A0 => b(24), A1 => b(23), SL => n1542, Z => n1009)
                           ;
   U1008 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1010, Z => n1313);
   U1009 : MUXB2DL port map( A0 => b(23), A1 => b(22), SL => n1542, Z => n1010)
                           ;
   U1010 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1011, Z => n1314);
   U1011 : MUXB2DL port map( A0 => b(22), A1 => b(21), SL => n1542, Z => n1011)
                           ;
   U1012 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1012, Z => n1315);
   U1013 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n1542, Z => n1012)
                           ;
   U1014 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1013, Z => n1316);
   U1015 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n1542, Z => n1013)
                           ;
   U1016 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1014, Z => n1317);
   U1017 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n1542, Z => n1014)
                           ;
   U1018 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1015, Z => n1318);
   U1019 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n1542, Z => n1015)
                           ;
   U1020 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1016, Z => n1319);
   U1021 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n1542, Z => n1016)
                           ;
   U1022 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1017, Z => n1320);
   U1023 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n1542, Z => n1017)
                           ;
   U1024 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1018, Z => n1321);
   U1025 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n1542, Z => n1018)
                           ;
   U1026 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1019, Z => n1322);
   U1027 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n1542, Z => n1019)
                           ;
   U1028 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1020, Z => n1323);
   U1029 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n1542, Z => n1020)
                           ;
   U1030 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1021, Z => n1324);
   U1031 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n1542, Z => n1021)
                           ;
   U1032 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1022, Z => n1325);
   U1033 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n1542, Z => n1022)
                           ;
   U1034 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1023, Z => n1326);
   U1035 : MUXB2DL port map( A0 => n1543, A1 => b(9), SL => n1542, Z => n1023);
   U1036 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1024, Z => n1327);
   U1037 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n1542, Z => n1024);
   U1038 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1025, Z => n1328);
   U1039 : MUXB2DL port map( A0 => n1545, A1 => b(7), SL => n1542, Z => n1025);
   U1040 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1026, Z => n1329);
   U1041 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n1542, Z => n1026);
   U1042 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1027, Z => n1330);
   U1043 : MUXB2DL port map( A0 => b(6), A1 => n1547, SL => n1542, Z => n1027);
   U1044 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1028, Z => n1331);
   U1045 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n1542, Z => n1028);
   U1046 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1029, Z => n1332);
   U1047 : MUXB2DL port map( A0 => n1549, A1 => n1551, SL => n1542, Z => n1029)
                           ;
   U1048 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1030, Z => n1333);
   U1049 : MUXB2DL port map( A0 => b(3), A1 => n1554, SL => n1542, Z => n1030);
   U1050 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1031, Z => n1334);
   U1051 : MUXB2DL port map( A0 => n1553, A1 => b(1), SL => n1542, Z => n1031);
   U1052 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1032, Z => n1335);
   U1053 : MUXB2DL port map( A0 => b(1), A1 => n1556, SL => n1542, Z => n1032);
   U1054 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1033, Z => n1336);
   U1055 : NAN2M1D1 port map( A1 => n1542, A2 => b(0), Z => n1033);
   U1056 : NOR2M1D1 port map( A1 => n3, A2 => n6, Z => n1096);
   U1057 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1034, Z => n1337);
   U1058 : MUXB2DL port map( A0 => b(31), A1 => b(30), SL => n8, Z => n1034);
   U1059 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1035, Z => n1338);
   U1060 : MUXB2DL port map( A0 => b(30), A1 => b(29), SL => n8, Z => n1035);
   U1061 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1036, Z => n1339);
   U1062 : MUXB2DL port map( A0 => b(29), A1 => b(28), SL => n8, Z => n1036);
   U1063 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1037, Z => n1340);
   U1064 : MUXB2DL port map( A0 => b(28), A1 => b(27), SL => n8, Z => n1037);
   U1065 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1038, Z => n1341);
   U1066 : MUXB2DL port map( A0 => b(27), A1 => b(26), SL => n8, Z => n1038);
   U1067 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1039, Z => n1342);
   U1068 : MUXB2DL port map( A0 => b(26), A1 => b(25), SL => n8, Z => n1039);
   U1069 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1040, Z => n1343);
   U1070 : MUXB2DL port map( A0 => b(25), A1 => b(24), SL => n8, Z => n1040);
   U1071 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1041, Z => n1344);
   U1072 : MUXB2DL port map( A0 => b(24), A1 => b(23), SL => n8, Z => n1041);
   U1073 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1042, Z => n1345);
   U1074 : MUXB2DL port map( A0 => b(23), A1 => b(22), SL => n8, Z => n1042);
   U1075 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1043, Z => n1346);
   U1076 : MUXB2DL port map( A0 => b(22), A1 => b(21), SL => n8, Z => n1043);
   U1077 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1044, Z => n1347);
   U1078 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n8, Z => n1044);
   U1079 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1045, Z => n1348);
   U1080 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n8, Z => n1045);
   U1081 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1046, Z => n1349);
   U1082 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n8, Z => n1046);
   U1083 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1047, Z => n1350);
   U1084 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n8, Z => n1047);
   U1085 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1048, Z => n1351);
   U1086 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n8, Z => n1048);
   U1087 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1049, Z => n1352);
   U1088 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n8, Z => n1049);
   U1089 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1050, Z => n1353);
   U1090 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n8, Z => n1050);
   U1091 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1051, Z => n1354);
   U1092 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n8, Z => n1051);
   U1093 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1052, Z => n1355);
   U1094 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n8, Z => n1052);
   U1095 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1053, Z => n1356);
   U1096 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n8, Z => n1053);
   U1097 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1054, Z => n1357);
   U1098 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n8, Z => n1054);
   U1099 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1055, Z => n1358);
   U1100 : MUXB2DL port map( A0 => n1543, A1 => b(9), SL => n8, Z => n1055);
   U1101 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1056, Z => n1359);
   U1102 : MUXB2DL port map( A0 => b(9), A1 => n1545, SL => n8, Z => n1056);
   U1103 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1057, Z => n1360);
   U1104 : MUXB2DL port map( A0 => n1545, A1 => b(7), SL => n8, Z => n1057);
   U1105 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1058, Z => n1361);
   U1106 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n8, Z => n1058);
   U1107 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1059, Z => n1362);
   U1108 : MUXB2DL port map( A0 => b(6), A1 => n1547, SL => n8, Z => n1059);
   U1109 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1060, Z => n1363);
   U1110 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n8, Z => n1060);
   U1111 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1061, Z => n1364);
   U1112 : MUXB2DL port map( A0 => n1549, A1 => n1551, SL => n8, Z => n1061);
   U1113 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1062, Z => n1365);
   U1114 : MUXB2DL port map( A0 => b(3), A1 => n1554, SL => n8, Z => n1062);
   U1115 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1063, Z => n1366);
   U1116 : MUXB2DL port map( A0 => n1553, A1 => b(1), SL => n8, Z => n1063);
   U1117 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1064, Z => n1367);
   U1118 : MUXB2DL port map( A0 => b(1), A1 => n1556, SL => n8, Z => n1064);
   U1119 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1065, Z => n1368);
   U1120 : NAN2M1D1 port map( A1 => n8, A2 => n1556, Z => n1065);
   U1121 : OAI21D1 port map( A1 => a(29), A2 => a(30), B => n1066, Z => n104);
   U1123 : EXNOR2D1 port map( A1 => a(29), A2 => a(30), Z => n106);
   U1125 : OAI21D1 port map( A1 => a(27), A2 => a(28), B => n1067, Z => n99);
   U1127 : EXNOR2D1 port map( A1 => a(27), A2 => a(28), Z => n103);
   U1129 : OAI21D1 port map( A1 => a(25), A2 => a(26), B => n1068, Z => n94);
   U1131 : EXNOR2D1 port map( A1 => a(25), A2 => a(26), Z => n98);
   U1135 : EXNOR2D1 port map( A1 => a(23), A2 => a(24), Z => n93);
   U1186 : ADHALFDL port map( A => n1278, B => n1093, CO => n780, S => n781);
   U1187 : OAI21D1 port map( A1 => a(1), A2 => a(2), B => n1080, Z => n1517);
   U1188 : OAI21D1 port map( A1 => a(3), A2 => a(4), B => n1079, Z => n1518);
   U1189 : OAI21D1 port map( A1 => a(7), A2 => a(8), B => n1077, Z => n1519);
   U1190 : AND2D1 port map( A1 => n1522, A2 => n305, Z => product(0));
   U1191 : AO21D1 port map( A1 => n215, A2 => n187, B => n188, Z => n1521);
   U1192 : OR2D1 port map( A1 => n1368, A2 => n1096, Z => n1522);
   U1193 : OA21M20D1 port map( A1 => n1523, A2 => n197, B => n194, Z => n190);
   U1194 : INVD1 port map( A => n215, Z => n214);
   U1195 : INVD1 port map( A => n233, Z => n232);
   U1196 : NAN2D1 port map( A1 => n313, A2 => n231, Z => n162);
   U1197 : INVD1 port map( A => n242, Z => n241);
   U1198 : INVD1 port map( A => n255, Z => n254);
   U1199 : INVD1 port map( A => n230, Z => n313);
   U1200 : INVD1 port map( A => n231, Z => n229);
   U1201 : INVD1 port map( A => n264, Z => n263);
   U1202 : NAN2D1 port map( A1 => n223, A2 => n1528, Z => n216);
   U1203 : INVD1 port map( A => n221, Z => n219);
   U1204 : NAN2D1 port map( A1 => n1530, A2 => n1529, Z => n243);
   U1205 : INVD1 port map( A => n248, Z => n246);
   U1206 : NAN2D1 port map( A1 => n1524, A2 => n1527, Z => n265);
   U1207 : INVD1 port map( A => n270, Z => n268);
   U1208 : NOR2D1 port map( A1 => n258, A2 => n261, Z => n256);
   U1209 : NOR2D1 port map( A1 => n236, A2 => n239, Z => n234);
   U1210 : NOR2D1 port map( A1 => n189, A2 => n201, Z => n187);
   U1211 : INVD1 port map( A => n209, Z => n211);
   U1212 : INVD1 port map( A => n206, Z => n204);
   U1213 : INVD1 port map( A => n275, Z => n273);
   U1214 : OR2D1 port map( A1 => n553, A2 => n574, Z => n1523);
   U1215 : NAN2D1 port map( A1 => n1523, A2 => n1526, Z => n189);
   U1216 : INVD1 port map( A => n199, Z => n197);
   U1217 : NAN2D1 port map( A1 => n667, A2 => n682, Z => n231);
   U1218 : INVD1 port map( A => n253, Z => n251);
   U1219 : NOR2D1 port map( A1 => n225, A2 => n230, Z => n223);
   U1220 : NAN2D1 port map( A1 => n1525, A2 => n310, Z => n201);
   U1221 : NOR2D1 port map( A1 => n683, A2 => n696, Z => n236);
   U1222 : NAN2D1 port map( A1 => n553, A2 => n574, Z => n194);
   U1223 : NOR2D1 port map( A1 => n667, A2 => n682, Z => n230);
   U1224 : INVD1 port map( A => n208, Z => n310);
   U1225 : NAN2D1 port map( A1 => n683, A2 => n696, Z => n237);
   U1226 : NAN2D1 port map( A1 => n1523, A2 => n194, Z => n156);
   U1227 : NAN2D1 port map( A1 => n1526, A2 => n199, Z => n157);
   U1228 : NAN2D1 port map( A1 => n1525, A2 => n206, Z => n158);
   U1229 : NAN2D1 port map( A1 => n310, A2 => n209, Z => n159);
   U1230 : NAN2D1 port map( A1 => n312, A2 => n226, Z => n161);
   U1231 : INVD1 port map( A => n225, Z => n312);
   U1232 : NAN2D1 port map( A1 => n1528, A2 => n221, Z => n160);
   U1233 : NAN2D1 port map( A1 => n314, A2 => n237, Z => n163);
   U1234 : INVD1 port map( A => n236, Z => n314);
   U1235 : NAN2D1 port map( A1 => n1530, A2 => n248, Z => n165);
   U1236 : NAN2D1 port map( A1 => n315, A2 => n240, Z => n164);
   U1237 : INVD1 port map( A => n239, Z => n315);
   U1238 : NAN2D1 port map( A1 => n1529, A2 => n253, Z => n166);
   U1239 : NAN2D1 port map( A1 => n318, A2 => n259, Z => n167);
   U1240 : INVD1 port map( A => n258, Z => n318);
   U1241 : NAN2D1 port map( A1 => n319, A2 => n262, Z => n168);
   U1242 : INVD1 port map( A => n261, Z => n319);
   U1243 : INVD1 port map( A => n277, Z => n276);
   U1244 : NAN2D1 port map( A1 => n1524, A2 => n270, Z => n169);
   U1245 : NAN2D1 port map( A1 => n1527, A2 => n275, Z => n170);
   U1246 : INVD1 port map( A => n286, Z => n285);
   U1247 : OR2D1 port map( A1 => n755, A2 => n762, Z => n1524);
   U1248 : NAN2D1 port map( A1 => n755, A2 => n762, Z => n270);
   U1249 : NOR2D1 port map( A1 => n280, A2 => n283, Z => n278);
   U1250 : OA21M20D1 port map( A1 => n1531, A2 => n294, B => n293, Z => n289);
   U1251 : NOR2D1 port map( A1 => n651, A2 => n666, Z => n225);
   U1252 : OA21M20D1 port map( A1 => n1532, A2 => n302, B => n301, Z => n297);
   U1253 : OR2D1 port map( A1 => n595, A2 => n614, Z => n1525);
   U1254 : NOR2D1 port map( A1 => n771, A2 => n776, Z => n280);
   U1255 : NOR2D1 port map( A1 => n745, A2 => n754, Z => n261);
   U1256 : NOR2D1 port map( A1 => n735, A2 => n744, Z => n258);
   U1257 : NAN2D1 port map( A1 => n763, A2 => n770, Z => n275);
   U1258 : OR2D1 port map( A1 => n575, A2 => n594, Z => n1526);
   U1259 : NAN2D1 port map( A1 => n575, A2 => n594, Z => n199);
   U1260 : NAN2D1 port map( A1 => n723, A2 => n734, Z => n253);
   U1261 : NAN2D1 port map( A1 => n651, A2 => n666, Z => n226);
   U1262 : OR2D1 port map( A1 => n763, A2 => n770, Z => n1527);
   U1263 : NAN2D1 port map( A1 => n595, A2 => n614, Z => n206);
   U1264 : OR2D1 port map( A1 => n633, A2 => n650, Z => n1528);
   U1265 : NAN2D1 port map( A1 => n745, A2 => n754, Z => n262);
   U1266 : OR2D1 port map( A1 => n723, A2 => n734, Z => n1529);
   U1267 : OR2D1 port map( A1 => n711, A2 => n722, Z => n1530);
   U1268 : NAN2D1 port map( A1 => n771, A2 => n776, Z => n281);
   U1269 : NAN2D1 port map( A1 => n615, A2 => n632, Z => n209);
   U1270 : NAN2D1 port map( A1 => n735, A2 => n744, Z => n259);
   U1271 : NOR2D1 port map( A1 => n697, A2 => n710, Z => n239);
   U1272 : NOR2D1 port map( A1 => n615, A2 => n632, Z => n208);
   U1273 : NAN2D1 port map( A1 => n633, A2 => n650, Z => n221);
   U1274 : NAN2D1 port map( A1 => n711, A2 => n722, Z => n248);
   U1275 : NAN2D1 port map( A1 => n697, A2 => n710, Z => n240);
   U1276 : NAN2D1 port map( A1 => n322, A2 => n281, Z => n171);
   U1277 : INVD1 port map( A => n280, Z => n322);
   U1278 : NAN2D1 port map( A1 => n323, A2 => n284, Z => n172);
   U1279 : INVD1 port map( A => n283, Z => n323);
   U1280 : NAN2D1 port map( A1 => n324, A2 => n288, Z => n173);
   U1281 : INVD1 port map( A => n287, Z => n324);
   U1282 : NAN2D1 port map( A1 => n1531, A2 => n293, Z => n174);
   U1283 : NAN2D1 port map( A1 => n326, A2 => n296, Z => n175);
   U1284 : INVD1 port map( A => n295, Z => n326);
   U1285 : NAN2D1 port map( A1 => n1532, A2 => n301, Z => n176);
   U1286 : EXOR2D1 port map( A1 => n178, A2 => n155, Z => product(31));
   U1287 : EXOR2D1 port map( A1 => n329, A2 => n344, Z => n155);
   U1288 : OR2D1 port map( A1 => n787, A2 => n789, Z => n1531);
   U1289 : OR2D1 port map( A1 => n793, A2 => n1366, Z => n1532);
   U1290 : NOR2D1 port map( A1 => n777, A2 => n782, Z => n283);
   U1291 : NAN2D1 port map( A1 => n787, A2 => n789, Z => n293);
   U1292 : NAN2D1 port map( A1 => n793, A2 => n1366, Z => n301);
   U1293 : NAN2D1 port map( A1 => n777, A2 => n782, Z => n284);
   U1294 : NOR2D1 port map( A1 => n783, A2 => n786, Z => n287);
   U1295 : NOR2D1 port map( A1 => n791, A2 => n792, Z => n295);
   U1296 : NAN2D1 port map( A1 => n783, A2 => n786, Z => n288);
   U1297 : NAN2D1 port map( A1 => n791, A2 => n792, Z => n296);
   U1298 : NAN2D1 port map( A1 => n1368, A2 => n1096, Z => n305);
   U1299 : NOR2D1 port map( A1 => n303, A2 => n305, Z => n302);
   U1300 : ADHALFDL port map( A => n1329, B => n1359, CO => n760, S => n761);
   U1301 : INVD1 port map( A => n1533, Z => n1542);
   U1302 : ADHALFDL port map( A => n1335, B => n1365, CO => n790, S => n791);
   U1303 : ADHALFDL port map( A => n1336, B => n1095, CO => n792, S => n793);
   U1304 : NOR2D1 port map( A1 => n1537, A2 => n30, Z => n1093);
   U1305 : INVD1 port map( A => n1535, Z => n1541);
   U1306 : ADHALFDL port map( A => n1331, B => n1361, CO => n774, S => n775);
   U1307 : INVD1 port map( A => n1534, Z => n1539);
   U1308 : ADHALFDL port map( A => n1252, B => n1092, CO => n768, S => n769);
   U1309 : ADHALFDL port map( A => n1333, B => n1363, CO => n784, S => n785);
   U1310 : INVD1 port map( A => n1536, Z => n1538);
   U1311 : ADHALFDL port map( A => n1306, B => n1094, CO => n788, S => n789);
   U1312 : INVD1 port map( A => n1537, Z => n1540);
   U1313 : INVD1 port map( A => n1548, Z => n1547);
   U1314 : INVD1 port map( A => n1555, Z => n1553);
   U1315 : INVD1 port map( A => n1546, Z => n1545);
   U1316 : INVD1 port map( A => n1544, Z => n1543);
   U1317 : INVD1 port map( A => n1555, Z => n1554);
   U1318 : INVD1 port map( A => n1552, Z => n1551);
   U1319 : INVD1 port map( A => n1557, Z => n1556);
   U1320 : INVD1 port map( A => n1550, Z => n1549);
   U1321 : ADHALFDL port map( A => n1206, B => n1090, CO => n732, S => n733);
   U1322 : ADHALFDL port map( A => n1168, B => n1088, CO => n680, S => n681);
   U1323 : ADHALFDL port map( A => n1152, B => n1087, CO => n648, S => n649);
   U1324 : ADHALFDL port map( A => n1228, B => n1091, CO => n752, S => n753);
   U1325 : ADHALFDL port map( A => n1186, B => n1089, CO => n708, S => n709);
   U1326 : ADHALFDL port map( A => n1138, B => n1086, CO => n612, S => n613);
   U1327 : INVD1 port map( A => n1367, Z => n303);
   U1328 : ADHALFDL port map( A => n1126, B => n1085, CO => n572, S => n573);
   U1329 : ADHALFDL port map( A => n1116, B => n1084, CO => n528, S => n529);
   U1330 : ADHALFDL port map( A => n1108, B => n1083, CO => n480, S => n481);
   U1331 : ADHALFDL port map( A => n1102, B => n1082, CO => n428, S => n429);
   U1332 : EXOR2D1 port map( A1 => n1307, A2 => n1337, Z => n343);
   U1333 : ADHALFDL port map( A => n1098, B => n1081, CO => n372, S => n373);
   U1334 : EXOR2D1 port map( A1 => a(1), A2 => a(2), Z => n1533);
   U1335 : ADHALFDL port map( A => n1323, B => n1353, CO => n694, S => n695);
   U1336 : EXOR2D1 port map( A1 => a(5), A2 => a(6), Z => n1534);
   U1337 : EXOR2D1 port map( A1 => a(3), A2 => a(4), Z => n1535);
   U1338 : EXOR2D1 port map( A1 => a(7), A2 => a(8), Z => n1536);
   U1339 : ADHALFDL port map( A => n1317, B => n1347, CO => n592, S => n593);
   U1340 : ADHALFDL port map( A => n1327, B => n1357, CO => n742, S => n743);
   U1341 : ADHALFDL port map( A => n1319, B => n1349, CO => n630, S => n631);
   U1342 : ADHALFDL port map( A => n1321, B => n1351, CO => n664, S => n665);
   U1343 : ADHALFDL port map( A => n1325, B => n1355, CO => n720, S => n721);
   U1344 : OA21D1 port map( A1 => a(5), A2 => a(6), B => n1078, Z => n1537);
   U1345 : INVD1 port map( A => a(3), Z => n1080);
   U1346 : EXNOR2D1 port map( A1 => a(11), A2 => a(12), Z => n56);
   U1347 : INVD1 port map( A => a(7), Z => n1078);
   U1348 : INVD1 port map( A => b(8), Z => n1546);
   U1349 : INVD1 port map( A => b(5), Z => n1548);
   U1350 : NAN2D1 port map( A1 => a(0), A2 => n6, Z => n3);
   U1351 : INVD1 port map( A => a(1), Z => n6);
   U1352 : INVD1 port map( A => b(2), Z => n1555);
   U1353 : INVD1 port map( A => b(10), Z => n1544);
   U1354 : INVD1 port map( A => a(9), Z => n1077);
   U1355 : INVD1 port map( A => b(3), Z => n1552);
   U1356 : EXNOR2D1 port map( A1 => a(13), A2 => a(14), Z => n63);
   U1357 : EXNOR2D1 port map( A1 => a(15), A2 => a(16), Z => n71);
   U1358 : INVD1 port map( A => b(4), Z => n1550);
   U1359 : INVD1 port map( A => a(5), Z => n1079);
   U1360 : INVD1 port map( A => b(0), Z => n1557);
   U1361 : EXNOR2D1 port map( A1 => a(9), A2 => a(10), Z => n48);
   U1362 : EXNOR2D1 port map( A1 => a(17), A2 => a(18), Z => n78);
   U1363 : AO21D1 port map( A1 => a(1), A2 => a(2), B => n1080, Z => n14);
   U1364 : AO21D1 port map( A1 => a(5), A2 => a(6), B => n1078, Z => n30);
   U1365 : EXNOR2D1 port map( A1 => a(19), A2 => a(20), Z => n83);
   U1366 : INVD1 port map( A => a(0), Z => n8);
   U1367 : AO21D1 port map( A1 => a(11), A2 => a(12), B => n1075, Z => n53);
   U1368 : INVD1 port map( A => a(13), Z => n1075);
   U1369 : ADHALFDL port map( A => n1315, B => n1345, CO => n550, S => n551);
   U1370 : AO21D1 port map( A1 => a(3), A2 => a(4), B => n1079, Z => n22);
   U1371 : AO21D1 port map( A1 => a(7), A2 => a(8), B => n1077, Z => n38);
   U1372 : OAI21D1 port map( A1 => a(11), A2 => a(12), B => n1075, Z => n50);
   U1373 : AO21D1 port map( A1 => a(13), A2 => a(14), B => n1074, Z => n61);
   U1374 : AO21D1 port map( A1 => a(15), A2 => a(16), B => n1073, Z => n69);
   U1375 : INVD1 port map( A => a(15), Z => n1074);
   U1376 : OAI21D1 port map( A1 => a(13), A2 => a(14), B => n1074, Z => n58);
   U1377 : INVD1 port map( A => a(17), Z => n1073);
   U1378 : OAI21D1 port map( A1 => a(15), A2 => a(16), B => n1073, Z => n66);
   U1379 : AO21D1 port map( A1 => a(9), A2 => a(10), B => n1076, Z => n45);
   U1380 : INVD1 port map( A => a(11), Z => n1076);
   U1381 : OAI21D1 port map( A1 => a(17), A2 => a(18), B => n1072, Z => n73);
   U1382 : INVD1 port map( A => a(19), Z => n1072);
   U1383 : OAI21D1 port map( A1 => a(9), A2 => a(10), B => n1076, Z => n42);
   U1384 : AO21D1 port map( A1 => a(17), A2 => a(18), B => n1072, Z => n76);
   U1385 : EXNOR2D1 port map( A1 => a(21), A2 => a(22), Z => n88);
   U1386 : OAI21D1 port map( A1 => a(19), A2 => a(20), B => n1071, Z => n79);
   U1387 : INVD1 port map( A => a(21), Z => n1071);
   U1388 : AO21D1 port map( A1 => a(19), A2 => a(20), B => n1071, Z => n81);
   U1389 : OAI21D1 port map( A1 => a(21), A2 => a(22), B => n1070, Z => n84);
   U1390 : INVD1 port map( A => a(23), Z => n1070);
   U1391 : AO21D1 port map( A1 => a(21), A2 => a(22), B => n1070, Z => n86);
   U1392 : ADHALFDL port map( A => n1313, B => n1343, CO => n504, S => n505);
   U1393 : OAI21D1 port map( A1 => a(23), A2 => a(24), B => n1069, Z => n89);
   U1394 : ADHALFDL port map( A => n1311, B => n1341, CO => n454, S => n455);
   U1395 : INVD1 port map( A => a(25), Z => n1069);
   U1396 : AO21D1 port map( A1 => a(23), A2 => a(24), B => n1069, Z => n91);
   U1397 : ADHALFDL port map( A => n1309, B => n1339, CO => n400, S => n401);
   U1398 : AO21D1 port map( A1 => a(25), A2 => a(26), B => n1068, Z => n96);
   U1399 : INVD1 port map( A => a(27), Z => n1068);
   U1400 : AO21D1 port map( A1 => a(27), A2 => a(28), B => n1067, Z => n101);
   U1401 : INVD1 port map( A => a(29), Z => n1067);
   U1402 : AO21D1 port map( A1 => a(29), A2 => a(30), B => n1066, Z => n105);
   U1403 : INVD1 port map( A => a(31), Z => n1066);

end hier_filter_none_5;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_gp_custom.all;

architecture hier_filter_none_5 of gp_custom_DW_mult_tc_7 is

   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AO21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component MUXB2DL
      port( A0, A1, SL : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component EXOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n6, n8, n14, n22, n30, n38, n42, n45, n48, n50, n53, n56, n58, 
      n61, n63, n66, n69, n71, n73, n76, n78, n79, n81, n83, n84, n86, n88, n89
      , n91, n93, n94, n96, n98, n99, n101, n103, n104, n105, n106, n155, n156,
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n178, n179, n180, n181, 
      n182, n183, n184, n185, n187, n188, n189, n190, n194, n195, n197, n199, 
      n200, n201, n202, n204, n206, n207, n208, n209, n211, n214, n215, n216, 
      n217, n219, n221, n222, n223, n224, n225, n226, n227, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n246, n248, n249, n251, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n268, n270, n271, n273, n275, 
      n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, 
      n288, n289, n293, n294, n295, n296, n297, n301, n302, n303, n305, n310, 
      n312, n313, n314, n315, n318, n319, n322, n323, n324, n326, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, 
      n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
      n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, 
      n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, 
      n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, 
      n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, 
      n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, 
      n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, 
      n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, 
      n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, 
      n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, 
      n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, 
      n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, 
      n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, 
      n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, 
      n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, 
      n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, 
      n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, 
      n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, 
      n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, 
      n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, 
      n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, 
      n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, 
      n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, 
      n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, 
      n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, 
      n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, 
      n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, 
      n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, 
      n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, 
      n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, 
      n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, 
      n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, 
      n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, 
      n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, 
      n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, 
      n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, 
      n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, 
      n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, 
      n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, 
      n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002
      , n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, 
      n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, 
      n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, 
      n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, 
      n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
      n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
      n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, 
      n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, 
      n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
      n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, 
      n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, 
      n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, 
      n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, 
      n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, 
      n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, 
      n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, 
      n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, 
      n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, 
      n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, 
      n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, 
      n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, 
      n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, 
      n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, 
      n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, 
      n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, 
      n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, 
      n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, 
      n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, 
      n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, 
      n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, 
      n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, 
      n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, 
      n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, 
      n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, 
      n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, 
      n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, 
      n1363, n1364, n1365, n1366, n1367, n1368, n1517, n1518, n1519, n1521, 
      n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, 
      n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, 
      n1542, n1543, n1544 : std_logic;

begin
   
   U125 : ADFULD1 port map( A => n345, B => n374, CI => n179, CO => n178, S => 
                           product(30));
   U126 : ADFULD1 port map( A => n375, B => n402, CI => n180, CO => n179, S => 
                           product(29));
   U127 : ADFULD1 port map( A => n403, B => n430, CI => n181, CO => n180, S => 
                           product(28));
   U128 : ADFULD1 port map( A => n431, B => n456, CI => n182, CO => n181, S => 
                           product(27));
   U129 : ADFULD1 port map( A => n457, B => n482, CI => n183, CO => n182, S => 
                           product(26));
   U130 : ADFULD1 port map( A => n483, B => n506, CI => n184, CO => n183, S => 
                           product(25));
   U131 : ADFULD1 port map( A => n507, B => n530, CI => n185, CO => n184, S => 
                           product(24));
   U132 : ADFULD1 port map( A => n531, B => n552, CI => n1521, CO => n185, S =>
                           product(23));
   U134 : EXOR2D1 port map( A1 => n195, A2 => n156, Z => product(22));
   U137 : OAI21D1 port map( A1 => n202, A2 => n189, B => n190, Z => n188);
   U146 : EXNOR2D1 port map( A1 => n200, A2 => n157, Z => product(21));
   U147 : AOI21D1 port map( A1 => n200, A2 => n1526, B => n197, Z => n195);
   U154 : EXNOR2D1 port map( A1 => n207, A2 => n158, Z => product(20));
   U155 : OAI21D1 port map( A1 => n214, A2 => n201, B => n202, Z => n200);
   U157 : AOI21D1 port map( A1 => n1525, A2 => n211, B => n204, Z => n202);
   U164 : EXOR2D1 port map( A1 => n214, A2 => n159, Z => product(19));
   U165 : OAI21D1 port map( A1 => n214, A2 => n208, B => n209, Z => n207);
   U174 : EXOR2D1 port map( A1 => n222, A2 => n160, Z => product(18));
   U176 : OAI21D1 port map( A1 => n233, A2 => n216, B => n217, Z => n215);
   U178 : AOI21D1 port map( A1 => n224, A2 => n1528, B => n219, Z => n217);
   U185 : EXOR2D1 port map( A1 => n227, A2 => n161, Z => product(17));
   U186 : AOI21D1 port map( A1 => n232, A2 => n223, B => n224, Z => n222);
   U188 : OAI21D1 port map( A1 => n225, A2 => n231, B => n226, Z => n224);
   U193 : EXNOR2D1 port map( A1 => n232, A2 => n162, Z => product(16));
   U194 : AOI21D1 port map( A1 => n232, A2 => n313, B => n229, Z => n227);
   U201 : EXNOR2D1 port map( A1 => n238, A2 => n163, Z => product(15));
   U203 : AOI21D1 port map( A1 => n242, A2 => n234, B => n235, Z => n233);
   U205 : OAI21D1 port map( A1 => n236, A2 => n240, B => n237, Z => n235);
   U210 : EXOR2D1 port map( A1 => n241, A2 => n164, Z => product(14));
   U211 : OAI21D1 port map( A1 => n241, A2 => n239, B => n240, Z => n238);
   U216 : EXOR2D1 port map( A1 => n249, A2 => n165, Z => product(13));
   U218 : OAI21D1 port map( A1 => n255, A2 => n243, B => n244, Z => n242);
   U220 : AOI21D1 port map( A1 => n1530, A2 => n251, B => n246, Z => n244);
   U227 : EXNOR2D1 port map( A1 => n254, A2 => n166, Z => product(12));
   U228 : AOI21D1 port map( A1 => n254, A2 => n1529, B => n251, Z => n249);
   U235 : EXNOR2D1 port map( A1 => n260, A2 => n167, Z => product(11));
   U237 : AOI21D1 port map( A1 => n256, A2 => n264, B => n257, Z => n255);
   U239 : OAI21D1 port map( A1 => n258, A2 => n262, B => n259, Z => n257);
   U244 : EXOR2D1 port map( A1 => n263, A2 => n168, Z => product(10));
   U245 : OAI21D1 port map( A1 => n263, A2 => n261, B => n262, Z => n260);
   U250 : EXOR2D1 port map( A1 => n271, A2 => n169, Z => product(9));
   U252 : OAI21D1 port map( A1 => n265, A2 => n277, B => n266, Z => n264);
   U254 : AOI21D1 port map( A1 => n1524, A2 => n273, B => n268, Z => n266);
   U261 : EXNOR2D1 port map( A1 => n276, A2 => n170, Z => product(8));
   U262 : AOI21D1 port map( A1 => n276, A2 => n1527, B => n273, Z => n271);
   U269 : EXNOR2D1 port map( A1 => n282, A2 => n171, Z => product(7));
   U271 : AOI21D1 port map( A1 => n278, A2 => n286, B => n279, Z => n277);
   U273 : OAI21D1 port map( A1 => n280, A2 => n284, B => n281, Z => n279);
   U278 : EXOR2D1 port map( A1 => n172, A2 => n285, Z => product(6));
   U279 : OAI21D1 port map( A1 => n285, A2 => n283, B => n284, Z => n282);
   U284 : EXOR2D1 port map( A1 => n173, A2 => n289, Z => product(5));
   U286 : OAI21D1 port map( A1 => n289, A2 => n287, B => n288, Z => n286);
   U291 : EXNOR2D1 port map( A1 => n174, A2 => n294, Z => product(4));
   U299 : EXOR2D1 port map( A1 => n297, A2 => n175, Z => product(3));
   U300 : OAI21D1 port map( A1 => n297, A2 => n295, B => n296, Z => n294);
   U305 : EXNOR2D1 port map( A1 => n176, A2 => n302, Z => product(2));
   U313 : EXOR2D1 port map( A1 => n303, A2 => n305, Z => product(1));
   U321 : EXOR3D1 port map( A1 => n346, A2 => n331, A3 => n330, Z => n329);
   U322 : EXOR3D1 port map( A1 => n332, A2 => n350, A3 => n348, Z => n330);
   U323 : EXOR3D1 port map( A1 => n352, A2 => n334, A3 => n333, Z => n331);
   U324 : EXOR3D1 port map( A1 => n354, A2 => n356, A3 => n335, Z => n332);
   U325 : EXOR3D1 port map( A1 => n337, A2 => n358, A3 => n336, Z => n333);
   U326 : EXOR3D1 port map( A1 => n339, A2 => n340, A3 => n360, Z => n334);
   U327 : EXOR3D1 port map( A1 => n342, A2 => n338, A3 => n341, Z => n335);
   U328 : EXOR3D1 port map( A1 => n366, A2 => n343, A3 => n362, Z => n336);
   U329 : EXOR3D1 port map( A1 => n368, A2 => n370, A3 => n364, Z => n337);
   U330 : EXOR3D1 port map( A1 => n1187, A2 => n1169, A3 => n372, Z => n338);
   U331 : EXOR3D1 port map( A1 => n1139, A2 => n1229, A3 => n1153, Z => n339);
   U332 : EXOR3D1 port map( A1 => n1103, A2 => n1117, A3 => n1109, Z => n340);
   U333 : EXOR3D1 port map( A1 => n1253, A2 => n1127, A3 => n1099, Z => n341);
   U334 : EXOR3D1 port map( A1 => n1097, A2 => n1279, A3 => n1207, Z => n342);
   U336 : ADFULD1 port map( A => n376, B => n349, CI => n347, CO => n344, S => 
                           n345);
   U337 : ADFULD1 port map( A => n351, B => n353, CI => n378, CO => n346, S => 
                           n347);
   U338 : ADFULD1 port map( A => n382, B => n355, CI => n380, CO => n348, S => 
                           n349);
   U339 : ADFULD1 port map( A => n359, B => n384, CI => n357, CO => n350, S => 
                           n351);
   U340 : ADFULD1 port map( A => n361, B => n388, CI => n386, CO => n352, S => 
                           n353);
   U341 : ADFULD1 port map( A => n365, B => n363, CI => n390, CO => n354, S => 
                           n355);
   U342 : ADFULD1 port map( A => n369, B => n371, CI => n367, CO => n356, S => 
                           n357);
   U343 : ADFULD1 port map( A => n398, B => n394, CI => n396, CO => n358, S => 
                           n359);
   U344 : ADFULD1 port map( A => n373, B => n400, CI => n392, CO => n360, S => 
                           n361);
   U345 : ADFULD1 port map( A => n1170, B => n1118, CI => n1140, CO => n362, S 
                           => n363);
   U346 : ADFULD1 port map( A => n1104, B => n1188, CI => n1110, CO => n364, S 
                           => n365);
   U347 : ADFULD1 port map( A => n1254, B => n1128, CI => n1230, CO => n366, S 
                           => n367);
   U348 : ADFULD1 port map( A => n1280, B => n1154, CI => n1208, CO => n368, S 
                           => n369);
   U349 : ADFULD1 port map( A => n1100, B => n1338, CI => n1308, CO => n370, S 
                           => n371);
   U351 : ADFULD1 port map( A => n404, B => n379, CI => n377, CO => n374, S => 
                           n375);
   U352 : ADFULD1 port map( A => n381, B => n408, CI => n406, CO => n376, S => 
                           n377);
   U353 : ADFULD1 port map( A => n410, B => n385, CI => n383, CO => n378, S => 
                           n379);
   U354 : ADFULD1 port map( A => n412, B => n389, CI => n387, CO => n380, S => 
                           n381);
   U355 : ADFULD1 port map( A => n391, B => n416, CI => n414, CO => n382, S => 
                           n383);
   U356 : ADFULD1 port map( A => n395, B => n397, CI => n399, CO => n384, S => 
                           n385);
   U357 : ADFULD1 port map( A => n418, B => n422, CI => n393, CO => n386, S => 
                           n387);
   U358 : ADFULD1 port map( A => n424, B => n426, CI => n420, CO => n388, S => 
                           n389);
   U359 : ADFULD1 port map( A => n428, B => n1171, CI => n401, CO => n390, S =>
                           n391);
   U360 : ADFULD1 port map( A => n1129, B => n1189, CI => n1141, CO => n392, S 
                           => n393);
   U361 : ADFULD1 port map( A => n1231, B => n1111, CI => n1105, CO => n394, S 
                           => n395);
   U362 : ADFULD1 port map( A => n1255, B => n1119, CI => n1101, CO => n396, S 
                           => n397);
   U363 : ADFULD1 port map( A => n1281, B => n1155, CI => n1209, CO => n398, S 
                           => n399);
   U365 : ADFULD1 port map( A => n432, B => n407, CI => n405, CO => n402, S => 
                           n403);
   U366 : ADFULD1 port map( A => n409, B => n436, CI => n434, CO => n404, S => 
                           n405);
   U367 : ADFULD1 port map( A => n438, B => n413, CI => n411, CO => n406, S => 
                           n407);
   U368 : ADFULD1 port map( A => n440, B => n417, CI => n415, CO => n408, S => 
                           n409);
   U369 : ADFULD1 port map( A => n444, B => n419, CI => n442, CO => n410, S => 
                           n411);
   U370 : ADFULD1 port map( A => n421, B => n423, CI => n425, CO => n412, S => 
                           n413);
   U371 : ADFULD1 port map( A => n448, B => n446, CI => n427, CO => n414, S => 
                           n415);
   U372 : ADFULD1 port map( A => n452, B => n429, CI => n450, CO => n416, S => 
                           n417);
   U373 : ADFULD1 port map( A => n1232, B => n1190, CI => n454, CO => n418, S 
                           => n419);
   U374 : ADFULD1 port map( A => n1142, B => n1256, CI => n1172, CO => n420, S 
                           => n421);
   U375 : ADFULD1 port map( A => n1112, B => n1130, CI => n1120, CO => n422, S 
                           => n423);
   U376 : ADFULD1 port map( A => n1282, B => n1156, CI => n1210, CO => n424, S 
                           => n425);
   U377 : ADFULD1 port map( A => n1106, B => n1340, CI => n1310, CO => n426, S 
                           => n427);
   U379 : ADFULD1 port map( A => n458, B => n435, CI => n433, CO => n430, S => 
                           n431);
   U380 : ADFULD1 port map( A => n437, B => n439, CI => n460, CO => n432, S => 
                           n433);
   U381 : ADFULD1 port map( A => n441, B => n464, CI => n462, CO => n434, S => 
                           n435);
   U382 : ADFULD1 port map( A => n466, B => n445, CI => n443, CO => n436, S => 
                           n437);
   U383 : ADFULD1 port map( A => n449, B => n451, CI => n468, CO => n438, S => 
                           n439);
   U384 : ADFULD1 port map( A => n453, B => n447, CI => n470, CO => n440, S => 
                           n441);
   U385 : ADFULD1 port map( A => n474, B => n472, CI => n476, CO => n442, S => 
                           n443);
   U386 : ADFULD1 port map( A => n455, B => n480, CI => n478, CO => n444, S => 
                           n445);
   U387 : ADFULD1 port map( A => n1131, B => n1191, CI => n1173, CO => n446, S 
                           => n447);
   U388 : ADFULD1 port map( A => n1113, B => n1233, CI => n1121, CO => n448, S 
                           => n449);
   U389 : ADFULD1 port map( A => n1283, B => n1143, CI => n1257, CO => n450, S 
                           => n451);
   U390 : ADFULD1 port map( A => n1107, B => n1157, CI => n1211, CO => n452, S 
                           => n453);
   U392 : ADFULD1 port map( A => n484, B => n461, CI => n459, CO => n456, S => 
                           n457);
   U393 : ADFULD1 port map( A => n486, B => n488, CI => n463, CO => n458, S => 
                           n459);
   U394 : ADFULD1 port map( A => n467, B => n469, CI => n465, CO => n460, S => 
                           n461);
   U395 : ADFULD1 port map( A => n492, B => n494, CI => n490, CO => n462, S => 
                           n463);
   U396 : ADFULD1 port map( A => n475, B => n477, CI => n471, CO => n464, S => 
                           n465);
   U397 : ADFULD1 port map( A => n479, B => n500, CI => n473, CO => n466, S => 
                           n467);
   U398 : ADFULD1 port map( A => n498, B => n502, CI => n496, CO => n468, S => 
                           n469);
   U399 : ADFULD1 port map( A => n504, B => n1192, CI => n481, CO => n470, S =>
                           n471);
   U400 : ADFULD1 port map( A => n1144, B => n1234, CI => n1158, CO => n472, S 
                           => n473);
   U401 : ADFULD1 port map( A => n1258, B => n1132, CI => n1122, CO => n474, S 
                           => n475);
   U402 : ADFULD1 port map( A => n1284, B => n1174, CI => n1212, CO => n476, S 
                           => n477);
   U403 : ADFULD1 port map( A => n1114, B => n1342, CI => n1312, CO => n478, S 
                           => n479);
   U405 : ADFULD1 port map( A => n508, B => n487, CI => n485, CO => n482, S => 
                           n483);
   U406 : ADFULD1 port map( A => n510, B => n512, CI => n489, CO => n484, S => 
                           n485);
   U407 : ADFULD1 port map( A => n493, B => n514, CI => n491, CO => n486, S => 
                           n487);
   U408 : ADFULD1 port map( A => n516, B => n518, CI => n495, CO => n488, S => 
                           n489);
   U409 : ADFULD1 port map( A => n501, B => n503, CI => n497, CO => n490, S => 
                           n491);
   U410 : ADFULD1 port map( A => n522, B => n524, CI => n499, CO => n492, S => 
                           n493);
   U411 : ADFULD1 port map( A => n526, B => n505, CI => n520, CO => n494, S => 
                           n495);
   U412 : ADFULD1 port map( A => n1235, B => n1259, CI => n528, CO => n496, S 
                           => n497);
   U413 : ADFULD1 port map( A => n1159, B => n1285, CI => n1193, CO => n498, S 
                           => n499);
   U414 : ADFULD1 port map( A => n1123, B => n1145, CI => n1133, CO => n500, S 
                           => n501);
   U415 : ADFULD1 port map( A => n1115, B => n1175, CI => n1213, CO => n502, S 
                           => n503);
   U417 : ADFULD1 port map( A => n532, B => n511, CI => n509, CO => n506, S => 
                           n507);
   U418 : ADFULD1 port map( A => n513, B => n536, CI => n534, CO => n508, S => 
                           n509);
   U419 : ADFULD1 port map( A => n517, B => n538, CI => n515, CO => n510, S => 
                           n511);
   U420 : ADFULD1 port map( A => n540, B => n542, CI => n519, CO => n512, S => 
                           n513);
   U421 : ADFULD1 port map( A => n525, B => n521, CI => n523, CO => n514, S => 
                           n515);
   U422 : ADFULD1 port map( A => n544, B => n546, CI => n527, CO => n516, S => 
                           n517);
   U423 : ADFULD1 port map( A => n529, B => n550, CI => n548, CO => n518, S => 
                           n519);
   U424 : ADFULD1 port map( A => n1194, B => n1260, CI => n1236, CO => n520, S 
                           => n521);
   U425 : ADFULD1 port map( A => n1134, B => n1286, CI => n1160, CO => n522, S 
                           => n523);
   U426 : ADFULD1 port map( A => n1124, B => n1176, CI => n1214, CO => n524, S 
                           => n525);
   U427 : ADFULD1 port map( A => n1146, B => n1344, CI => n1314, CO => n526, S 
                           => n527);
   U429 : ADFULD1 port map( A => n554, B => n535, CI => n533, CO => n530, S => 
                           n531);
   U430 : ADFULD1 port map( A => n556, B => n539, CI => n537, CO => n532, S => 
                           n533);
   U431 : ADFULD1 port map( A => n541, B => n560, CI => n558, CO => n534, S => 
                           n535);
   U432 : ADFULD1 port map( A => n562, B => n545, CI => n543, CO => n536, S => 
                           n537);
   U433 : ADFULD1 port map( A => n549, B => n564, CI => n547, CO => n538, S => 
                           n539);
   U434 : ADFULD1 port map( A => n566, B => n570, CI => n568, CO => n540, S => 
                           n541);
   U435 : ADFULD1 port map( A => n572, B => n1195, CI => n551, CO => n542, S =>
                           n543);
   U436 : ADFULD1 port map( A => n1135, B => n1237, CI => n1147, CO => n544, S 
                           => n545);
   U437 : ADFULD1 port map( A => n1287, B => n1161, CI => n1261, CO => n546, S 
                           => n547);
   U438 : ADFULD1 port map( A => n1125, B => n1177, CI => n1215, CO => n548, S 
                           => n549);
   U440 : ADFULD1 port map( A => n576, B => n557, CI => n555, CO => n552, S => 
                           n553);
   U441 : ADFULD1 port map( A => n559, B => n561, CI => n578, CO => n554, S => 
                           n555);
   U442 : ADFULD1 port map( A => n563, B => n582, CI => n580, CO => n556, S => 
                           n557);
   U443 : ADFULD1 port map( A => n565, B => n569, CI => n584, CO => n558, S => 
                           n559);
   U444 : ADFULD1 port map( A => n571, B => n586, CI => n567, CO => n560, S => 
                           n561);
   U445 : ADFULD1 port map( A => n590, B => n573, CI => n588, CO => n562, S => 
                           n563);
   U446 : ADFULD1 port map( A => n1196, B => n1238, CI => n592, CO => n564, S 
                           => n565);
   U447 : ADFULD1 port map( A => n1148, B => n1262, CI => n1162, CO => n566, S 
                           => n567);
   U448 : ADFULD1 port map( A => n1288, B => n1178, CI => n1216, CO => n568, S 
                           => n569);
   U449 : ADFULD1 port map( A => n1136, B => n1346, CI => n1316, CO => n570, S 
                           => n571);
   U451 : ADFULD1 port map( A => n596, B => n579, CI => n577, CO => n574, S => 
                           n575);
   U452 : ADFULD1 port map( A => n581, B => n583, CI => n598, CO => n576, S => 
                           n577);
   U453 : ADFULD1 port map( A => n585, B => n602, CI => n600, CO => n578, S => 
                           n579);
   U454 : ADFULD1 port map( A => n591, B => n589, CI => n604, CO => n580, S => 
                           n581);
   U455 : ADFULD1 port map( A => n606, B => n608, CI => n587, CO => n582, S => 
                           n583);
   U456 : ADFULD1 port map( A => n593, B => n612, CI => n610, CO => n584, S => 
                           n585);
   U457 : ADFULD1 port map( A => n1163, B => n1239, CI => n1197, CO => n586, S 
                           => n587);
   U458 : ADFULD1 port map( A => n1263, B => n1149, CI => n1137, CO => n588, S 
                           => n589);
   U459 : ADFULD1 port map( A => n1289, B => n1179, CI => n1217, CO => n590, S 
                           => n591);
   U461 : ADFULD1 port map( A => n616, B => n599, CI => n597, CO => n594, S => 
                           n595);
   U462 : ADFULD1 port map( A => n601, B => n603, CI => n618, CO => n596, S => 
                           n597);
   U463 : ADFULD1 port map( A => n622, B => n605, CI => n620, CO => n598, S => 
                           n599);
   U464 : ADFULD1 port map( A => n609, B => n611, CI => n607, CO => n600, S => 
                           n601);
   U465 : ADFULD1 port map( A => n626, B => n628, CI => n624, CO => n602, S => 
                           n603);
   U466 : ADFULD1 port map( A => n630, B => n1240, CI => n613, CO => n604, S =>
                           n605);
   U467 : ADFULD1 port map( A => n1150, B => n1264, CI => n1180, CO => n606, S 
                           => n607);
   U468 : ADFULD1 port map( A => n1290, B => n1198, CI => n1218, CO => n608, S 
                           => n609);
   U469 : ADFULD1 port map( A => n1164, B => n1348, CI => n1318, CO => n610, S 
                           => n611);
   U471 : ADFULD1 port map( A => n634, B => n619, CI => n617, CO => n614, S => 
                           n615);
   U472 : ADFULD1 port map( A => n621, B => n623, CI => n636, CO => n616, S => 
                           n617);
   U473 : ADFULD1 port map( A => n640, B => n625, CI => n638, CO => n618, S => 
                           n619);
   U474 : ADFULD1 port map( A => n627, B => n644, CI => n629, CO => n620, S => 
                           n621);
   U475 : ADFULD1 port map( A => n646, B => n631, CI => n642, CO => n622, S => 
                           n623);
   U476 : ADFULD1 port map( A => n1241, B => n1265, CI => n648, CO => n624, S 
                           => n625);
   U477 : ADFULD1 port map( A => n1291, B => n1181, CI => n1165, CO => n626, S 
                           => n627);
   U478 : ADFULD1 port map( A => n1151, B => n1199, CI => n1219, CO => n628, S 
                           => n629);
   U480 : ADFULD1 port map( A => n652, B => n637, CI => n635, CO => n632, S => 
                           n633);
   U481 : ADFULD1 port map( A => n639, B => n641, CI => n654, CO => n634, S => 
                           n635);
   U482 : ADFULD1 port map( A => n658, B => n645, CI => n656, CO => n636, S => 
                           n637);
   U483 : ADFULD1 port map( A => n647, B => n660, CI => n643, CO => n638, S => 
                           n639);
   U484 : ADFULD1 port map( A => n649, B => n664, CI => n662, CO => n640, S => 
                           n641);
   U485 : ADFULD1 port map( A => n1182, B => n1292, CI => n1242, CO => n642, S 
                           => n643);
   U486 : ADFULD1 port map( A => n1166, B => n1266, CI => n1220, CO => n644, S 
                           => n645);
   U487 : ADFULD1 port map( A => n1200, B => n1350, CI => n1320, CO => n646, S 
                           => n647);
   U489 : ADFULD1 port map( A => n668, B => n655, CI => n653, CO => n650, S => 
                           n651);
   U490 : ADFULD1 port map( A => n670, B => n659, CI => n657, CO => n652, S => 
                           n653);
   U491 : ADFULD1 port map( A => n663, B => n661, CI => n672, CO => n654, S => 
                           n655);
   U492 : ADFULD1 port map( A => n676, B => n678, CI => n674, CO => n656, S => 
                           n657);
   U493 : ADFULD1 port map( A => n680, B => n1267, CI => n665, CO => n658, S =>
                           n659);
   U494 : ADFULD1 port map( A => n1183, B => n1167, CI => n1243, CO => n660, S 
                           => n661);
   U495 : ADFULD1 port map( A => n1293, B => n1201, CI => n1221, CO => n662, S 
                           => n663);
   U497 : ADFULD1 port map( A => n684, B => n671, CI => n669, CO => n666, S => 
                           n667);
   U498 : ADFULD1 port map( A => n686, B => n688, CI => n673, CO => n668, S => 
                           n669);
   U499 : ADFULD1 port map( A => n677, B => n679, CI => n675, CO => n670, S => 
                           n671);
   U500 : ADFULD1 port map( A => n692, B => n681, CI => n690, CO => n672, S => 
                           n673);
   U501 : ADFULD1 port map( A => n1244, B => n1294, CI => n694, CO => n674, S 
                           => n675);
   U502 : ADFULD1 port map( A => n1184, B => n1268, CI => n1222, CO => n676, S 
                           => n677);
   U503 : ADFULD1 port map( A => n1202, B => n1352, CI => n1322, CO => n678, S 
                           => n679);
   U505 : ADFULD1 port map( A => n698, B => n687, CI => n685, CO => n682, S => 
                           n683);
   U506 : ADFULD1 port map( A => n700, B => n702, CI => n689, CO => n684, S => 
                           n685);
   U507 : ADFULD1 port map( A => n691, B => n704, CI => n693, CO => n686, S => 
                           n687);
   U508 : ADFULD1 port map( A => n695, B => n708, CI => n706, CO => n688, S => 
                           n689);
   U509 : ADFULD1 port map( A => n1185, B => n1245, CI => n1203, CO => n690, S 
                           => n691);
   U510 : ADFULD1 port map( A => n1295, B => n1269, CI => n1223, CO => n692, S 
                           => n693);
   U512 : ADFULD1 port map( A => n712, B => n701, CI => n699, CO => n696, S => 
                           n697);
   U513 : ADFULD1 port map( A => n703, B => n705, CI => n714, CO => n698, S => 
                           n699);
   U514 : ADFULD1 port map( A => n716, B => n718, CI => n707, CO => n700, S => 
                           n701);
   U515 : ADFULD1 port map( A => n720, B => n1270, CI => n709, CO => n702, S =>
                           n703);
   U516 : ADFULD1 port map( A => n1246, B => n1296, CI => n1224, CO => n704, S 
                           => n705);
   U517 : ADFULD1 port map( A => n1204, B => n1354, CI => n1324, CO => n706, S 
                           => n707);
   U519 : ADFULD1 port map( A => n724, B => n715, CI => n713, CO => n710, S => 
                           n711);
   U520 : ADFULD1 port map( A => n717, B => n719, CI => n726, CO => n712, S => 
                           n713);
   U521 : ADFULD1 port map( A => n730, B => n721, CI => n728, CO => n714, S => 
                           n715);
   U522 : ADFULD1 port map( A => n1205, B => n1247, CI => n732, CO => n716, S 
                           => n717);
   U523 : ADFULD1 port map( A => n1271, B => n1297, CI => n1225, CO => n718, S 
                           => n719);
   U525 : ADFULD1 port map( A => n736, B => n727, CI => n725, CO => n722, S => 
                           n723);
   U526 : ADFULD1 port map( A => n729, B => n731, CI => n738, CO => n724, S => 
                           n725);
   U527 : ADFULD1 port map( A => n733, B => n742, CI => n740, CO => n726, S => 
                           n727);
   U528 : ADFULD1 port map( A => n1272, B => n1298, CI => n1226, CO => n728, S 
                           => n729);
   U529 : ADFULD1 port map( A => n1248, B => n1356, CI => n1326, CO => n730, S 
                           => n731);
   U531 : ADFULD1 port map( A => n746, B => n739, CI => n737, CO => n734, S => 
                           n735);
   U532 : ADFULD1 port map( A => n748, B => n750, CI => n741, CO => n736, S => 
                           n737);
   U533 : ADFULD1 port map( A => n752, B => n1299, CI => n743, CO => n738, S =>
                           n739);
   U534 : ADFULD1 port map( A => n1273, B => n1249, CI => n1227, CO => n740, S 
                           => n741);
   U536 : ADFULD1 port map( A => n756, B => n749, CI => n747, CO => n744, S => 
                           n745);
   U537 : ADFULD1 port map( A => n758, B => n753, CI => n751, CO => n746, S => 
                           n747);
   U538 : ADFULD1 port map( A => n1274, B => n1300, CI => n760, CO => n748, S 
                           => n749);
   U539 : ADFULD1 port map( A => n1250, B => n1358, CI => n1328, CO => n750, S 
                           => n751);
   U541 : ADFULD1 port map( A => n764, B => n759, CI => n757, CO => n754, S => 
                           n755);
   U542 : ADFULD1 port map( A => n761, B => n768, CI => n766, CO => n756, S => 
                           n757);
   U543 : ADFULD1 port map( A => n1275, B => n1251, CI => n1301, CO => n758, S 
                           => n759);
   U545 : ADFULD1 port map( A => n767, B => n772, CI => n765, CO => n762, S => 
                           n763);
   U546 : ADFULD1 port map( A => n774, B => n1302, CI => n769, CO => n764, S =>
                           n765);
   U547 : ADFULD1 port map( A => n1276, B => n1360, CI => n1330, CO => n766, S 
                           => n767);
   U549 : ADFULD1 port map( A => n778, B => n775, CI => n773, CO => n770, S => 
                           n771);
   U550 : ADFULD1 port map( A => n1277, B => n1303, CI => n780, CO => n772, S 
                           => n773);
   U552 : ADFULD1 port map( A => n781, B => n784, CI => n779, CO => n776, S => 
                           n777);
   U553 : ADFULD1 port map( A => n1304, B => n1362, CI => n1332, CO => n778, S 
                           => n779);
   U555 : ADFULD1 port map( A => n788, B => n1305, CI => n785, CO => n782, S =>
                           n783);
   U557 : ADFULD1 port map( A => n1334, B => n1364, CI => n790, CO => n786, S 
                           => n787);
   U561 : NOR2M1D1 port map( A1 => n104, A2 => n105, Z => n1081);
   U562 : MUXB2DL port map( A0 => n104, A1 => n105, SL => n794, Z => n1097);
   U563 : MUXB2DL port map( A0 => b(1), A1 => n1543, SL => n106, Z => n794);
   U564 : MUXB2DL port map( A0 => n104, A1 => n105, SL => n795, Z => n1098);
   U565 : NAN2M1D1 port map( A1 => n106, A2 => b(0), Z => n795);
   U566 : NOR2M1D1 port map( A1 => n99, A2 => n101, Z => n1082);
   U567 : MUXB2DL port map( A0 => n99, A1 => n101, SL => n796, Z => n1099);
   U568 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n103, Z => n796);
   U569 : MUXB2DL port map( A0 => n99, A1 => n101, SL => n797, Z => n1100);
   U570 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n103, Z => n797);
   U571 : MUXB2DL port map( A0 => n99, A1 => n101, SL => n798, Z => n1101);
   U572 : MUXB2DL port map( A0 => b(1), A1 => n1543, SL => n103, Z => n798);
   U573 : MUXB2DL port map( A0 => n99, A1 => n101, SL => n799, Z => n1102);
   U574 : NAN2M1D1 port map( A1 => n103, A2 => b(0), Z => n799);
   U575 : NOR2M1D1 port map( A1 => n94, A2 => n96, Z => n1083);
   U576 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n800, Z => n1103);
   U577 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n98, Z => n800);
   U578 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n801, Z => n1104);
   U579 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n98, Z => n801);
   U580 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n802, Z => n1105);
   U581 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n98, Z => n802);
   U582 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n803, Z => n1106);
   U583 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n98, Z => n803);
   U584 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n804, Z => n1107);
   U585 : MUXB2DL port map( A0 => b(1), A1 => n1543, SL => n98, Z => n804);
   U586 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n805, Z => n1108);
   U587 : NAN2M1D1 port map( A1 => n98, A2 => b(0), Z => n805);
   U588 : NOR2M1D1 port map( A1 => n89, A2 => n91, Z => n1084);
   U589 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n806, Z => n1109);
   U590 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n93, Z => n806);
   U591 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n807, Z => n1110);
   U592 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n93, Z => n807);
   U593 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n808, Z => n1111);
   U594 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n93, Z => n808);
   U595 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n809, Z => n1112);
   U596 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n93, Z => n809);
   U597 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n810, Z => n1113);
   U598 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n93, Z => n810);
   U599 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n811, Z => n1114);
   U600 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n93, Z => n811);
   U601 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n812, Z => n1115);
   U602 : MUXB2DL port map( A0 => b(1), A1 => n1543, SL => n93, Z => n812);
   U603 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n813, Z => n1116);
   U604 : NAN2M1D1 port map( A1 => n93, A2 => n1543, Z => n813);
   U605 : NOR2M1D1 port map( A1 => n84, A2 => n86, Z => n1085);
   U606 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n814, Z => n1117);
   U607 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n88, Z => n814);
   U608 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n815, Z => n1118);
   U609 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n88, Z => n815);
   U610 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n816, Z => n1119);
   U611 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n88, Z => n816);
   U612 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n817, Z => n1120);
   U613 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n88, Z => n817);
   U614 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n818, Z => n1121);
   U615 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n88, Z => n818);
   U616 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n819, Z => n1122);
   U617 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n88, Z => n819);
   U618 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n820, Z => n1123);
   U619 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n88, Z => n820);
   U620 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n821, Z => n1124);
   U621 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n88, Z => n821);
   U622 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n822, Z => n1125);
   U623 : MUXB2DL port map( A0 => b(1), A1 => n1543, SL => n88, Z => n822);
   U624 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n823, Z => n1126);
   U625 : NAN2M1D1 port map( A1 => n88, A2 => n1543, Z => n823);
   U626 : NOR2M1D1 port map( A1 => n79, A2 => n81, Z => n1086);
   U627 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n824, Z => n1127);
   U628 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n83, Z => n824);
   U629 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n825, Z => n1128);
   U630 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n83, Z => n825);
   U631 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n826, Z => n1129);
   U632 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n83, Z => n826);
   U633 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n827, Z => n1130);
   U634 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n83, Z => n827);
   U635 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n828, Z => n1131);
   U636 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n83, Z => n828);
   U637 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n829, Z => n1132);
   U638 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n83, Z => n829);
   U639 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n830, Z => n1133);
   U640 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n83, Z => n830);
   U641 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n831, Z => n1134);
   U642 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n83, Z => n831);
   U643 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n832, Z => n1135);
   U644 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n83, Z => n832);
   U645 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n833, Z => n1136);
   U646 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n83, Z => n833);
   U647 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n834, Z => n1137);
   U648 : MUXB2DL port map( A0 => b(1), A1 => n1543, SL => n83, Z => n834);
   U649 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n835, Z => n1138);
   U650 : NAN2M1D1 port map( A1 => n83, A2 => b(0), Z => n835);
   U651 : NOR2M1D1 port map( A1 => n73, A2 => n76, Z => n1087);
   U652 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n836, Z => n1139);
   U653 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n78, Z => n836);
   U654 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n837, Z => n1140);
   U655 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n78, Z => n837);
   U656 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n838, Z => n1141);
   U657 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n78, Z => n838);
   U658 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n839, Z => n1142);
   U659 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n78, Z => n839);
   U660 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n840, Z => n1143);
   U661 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n78, Z => n840);
   U662 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n841, Z => n1144);
   U663 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n78, Z => n841);
   U664 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n842, Z => n1145);
   U665 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n78, Z => n842);
   U666 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n843, Z => n1146);
   U667 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n78, Z => n843);
   U668 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n844, Z => n1147);
   U669 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n78, Z => n844);
   U670 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n845, Z => n1148);
   U671 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n78, Z => n845);
   U672 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n846, Z => n1149);
   U673 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n78, Z => n846);
   U674 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n847, Z => n1150);
   U675 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n78, Z => n847);
   U676 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n848, Z => n1151);
   U677 : MUXB2DL port map( A0 => b(1), A1 => n1543, SL => n78, Z => n848);
   U678 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n849, Z => n1152);
   U679 : NAN2M1D1 port map( A1 => n78, A2 => n1543, Z => n849);
   U680 : NOR2M1D1 port map( A1 => n66, A2 => n69, Z => n1088);
   U681 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n850, Z => n1153);
   U682 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n71, Z => n850);
   U683 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n851, Z => n1154);
   U684 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n71, Z => n851);
   U685 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n852, Z => n1155);
   U686 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n71, Z => n852);
   U687 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n853, Z => n1156);
   U688 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n71, Z => n853);
   U689 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n854, Z => n1157);
   U690 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n71, Z => n854);
   U691 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n855, Z => n1158);
   U692 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n71, Z => n855);
   U693 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n856, Z => n1159);
   U694 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n71, Z => n856);
   U695 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n857, Z => n1160);
   U696 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n71, Z => n857);
   U697 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n858, Z => n1161);
   U698 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n71, Z => n858);
   U699 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n859, Z => n1162);
   U700 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n71, Z => n859);
   U701 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n860, Z => n1163);
   U702 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n71, Z => n860);
   U703 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n861, Z => n1164);
   U704 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n71, Z => n861);
   U705 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n862, Z => n1165);
   U706 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n71, Z => n862);
   U707 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n863, Z => n1166);
   U708 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n71, Z => n863);
   U709 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n864, Z => n1167);
   U710 : MUXB2DL port map( A0 => b(1), A1 => n1543, SL => n71, Z => n864);
   U711 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n865, Z => n1168);
   U712 : NAN2M1D1 port map( A1 => n71, A2 => b(0), Z => n865);
   U713 : NOR2M1D1 port map( A1 => n58, A2 => n61, Z => n1089);
   U714 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n866, Z => n1169);
   U715 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n63, Z => n866);
   U716 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n867, Z => n1170);
   U717 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n63, Z => n867);
   U718 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n868, Z => n1171);
   U719 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n63, Z => n868);
   U720 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n869, Z => n1172);
   U721 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n63, Z => n869);
   U722 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n870, Z => n1173);
   U723 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n63, Z => n870);
   U724 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n871, Z => n1174);
   U725 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n63, Z => n871);
   U726 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n872, Z => n1175);
   U727 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n63, Z => n872);
   U728 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n873, Z => n1176);
   U729 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n63, Z => n873);
   U730 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n874, Z => n1177);
   U731 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n63, Z => n874);
   U732 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n875, Z => n1178);
   U733 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n63, Z => n875);
   U734 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n876, Z => n1179);
   U735 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n63, Z => n876);
   U736 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n877, Z => n1180);
   U737 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n63, Z => n877);
   U738 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n878, Z => n1181);
   U739 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n63, Z => n878);
   U740 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n879, Z => n1182);
   U741 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n63, Z => n879);
   U742 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n880, Z => n1183);
   U743 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n63, Z => n880);
   U744 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n881, Z => n1184);
   U745 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n63, Z => n881);
   U746 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n882, Z => n1185);
   U747 : MUXB2DL port map( A0 => b(1), A1 => n1543, SL => n63, Z => n882);
   U748 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n883, Z => n1186);
   U749 : NAN2M1D1 port map( A1 => n63, A2 => b(0), Z => n883);
   U750 : NOR2M1D1 port map( A1 => n50, A2 => n53, Z => n1090);
   U751 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n884, Z => n1187);
   U752 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n56, Z => n884);
   U753 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n885, Z => n1188);
   U754 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n56, Z => n885);
   U755 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n886, Z => n1189);
   U756 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n56, Z => n886);
   U757 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n887, Z => n1190);
   U758 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n56, Z => n887);
   U759 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n888, Z => n1191);
   U760 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n56, Z => n888);
   U761 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n889, Z => n1192);
   U762 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n56, Z => n889);
   U763 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n890, Z => n1193);
   U764 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n56, Z => n890);
   U765 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n891, Z => n1194);
   U766 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n56, Z => n891);
   U767 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n892, Z => n1195);
   U768 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n56, Z => n892);
   U769 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n893, Z => n1196);
   U770 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n56, Z => n893);
   U771 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n894, Z => n1197);
   U772 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n56, Z => n894);
   U773 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n895, Z => n1198);
   U774 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n56, Z => n895);
   U775 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n896, Z => n1199);
   U776 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n56, Z => n896);
   U777 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n897, Z => n1200);
   U778 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n56, Z => n897);
   U779 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n898, Z => n1201);
   U780 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n56, Z => n898);
   U781 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n899, Z => n1202);
   U782 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n56, Z => n899);
   U783 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n900, Z => n1203);
   U784 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n56, Z => n900);
   U785 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n901, Z => n1204);
   U786 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n56, Z => n901);
   U787 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n902, Z => n1205);
   U788 : MUXB2DL port map( A0 => b(1), A1 => b(0), SL => n56, Z => n902);
   U789 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n903, Z => n1206);
   U790 : NAN2M1D1 port map( A1 => n56, A2 => n1543, Z => n903);
   U791 : NOR2M1D1 port map( A1 => n42, A2 => n45, Z => n1091);
   U792 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n904, Z => n1207);
   U793 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n48, Z => n904);
   U794 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n905, Z => n1208);
   U795 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n48, Z => n905);
   U796 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n906, Z => n1209);
   U797 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n48, Z => n906);
   U798 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n907, Z => n1210);
   U799 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n48, Z => n907);
   U800 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n908, Z => n1211);
   U801 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n48, Z => n908);
   U802 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n909, Z => n1212);
   U803 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n48, Z => n909);
   U804 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n910, Z => n1213);
   U805 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n48, Z => n910);
   U806 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n911, Z => n1214);
   U807 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n48, Z => n911);
   U808 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n912, Z => n1215);
   U809 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n48, Z => n912);
   U810 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n913, Z => n1216);
   U811 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n48, Z => n913);
   U812 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n914, Z => n1217);
   U813 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n48, Z => n914);
   U814 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n915, Z => n1218);
   U815 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n48, Z => n915);
   U816 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n916, Z => n1219);
   U817 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n48, Z => n916);
   U818 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n917, Z => n1220);
   U819 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n48, Z => n917);
   U820 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n918, Z => n1221);
   U821 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n48, Z => n918);
   U822 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n919, Z => n1222);
   U823 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n48, Z => n919);
   U824 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n920, Z => n1223);
   U825 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n48, Z => n920);
   U826 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n921, Z => n1224);
   U827 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n48, Z => n921);
   U828 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n922, Z => n1225);
   U829 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n48, Z => n922);
   U830 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n923, Z => n1226);
   U831 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n48, Z => n923);
   U832 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n924, Z => n1227);
   U833 : MUXB2DL port map( A0 => b(1), A1 => b(0), SL => n48, Z => n924);
   U834 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n925, Z => n1228);
   U835 : NAN2M1D1 port map( A1 => n48, A2 => b(0), Z => n925);
   U836 : NOR2M1D1 port map( A1 => n1519, A2 => n38, Z => n1092);
   U837 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n926, Z => n1229);
   U838 : MUXB2DL port map( A0 => b(23), A1 => b(22), SL => n1538, Z => n926);
   U839 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n927, Z => n1230);
   U840 : MUXB2DL port map( A0 => b(22), A1 => b(21), SL => n1538, Z => n927);
   U841 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n928, Z => n1231);
   U842 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n1538, Z => n928);
   U843 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n929, Z => n1232);
   U844 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n1538, Z => n929);
   U845 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n930, Z => n1233);
   U846 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n1538, Z => n930);
   U847 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n931, Z => n1234);
   U848 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n1538, Z => n931);
   U849 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n932, Z => n1235);
   U850 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n1538, Z => n932);
   U851 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n933, Z => n1236);
   U852 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n1538, Z => n933);
   U853 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n934, Z => n1237);
   U854 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n1538, Z => n934);
   U855 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n935, Z => n1238);
   U856 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n1538, Z => n935);
   U857 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n936, Z => n1239);
   U858 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n1538, Z => n936);
   U859 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n937, Z => n1240);
   U860 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n1538, Z => n937);
   U861 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n938, Z => n1241);
   U862 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n1538, Z => n938);
   U863 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n939, Z => n1242);
   U864 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n1538, Z => n939);
   U865 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n940, Z => n1243);
   U866 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n1538, Z => n940);
   U867 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n941, Z => n1244);
   U868 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n1538, Z => n941);
   U869 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n942, Z => n1245);
   U870 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n1538, Z => n942);
   U871 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n943, Z => n1246);
   U872 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n1538, Z => n943);
   U873 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n944, Z => n1247);
   U874 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n1538, Z => n944);
   U875 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n945, Z => n1248);
   U876 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n1538, Z => n945);
   U877 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n946, Z => n1249);
   U878 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n1538, Z => n946);
   U879 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n947, Z => n1250);
   U880 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n1538, Z => n947);
   U881 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n948, Z => n1251);
   U882 : MUXB2DL port map( A0 => b(1), A1 => b(0), SL => n1538, Z => n948);
   U883 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n949, Z => n1252);
   U884 : NAN2M1D1 port map( A1 => n1538, A2 => b(0), Z => n949);
   U886 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n950, Z => n1253);
   U887 : MUXB2DL port map( A0 => b(25), A1 => b(24), SL => n1539, Z => n950);
   U888 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n951, Z => n1254);
   U889 : MUXB2DL port map( A0 => b(24), A1 => b(23), SL => n1539, Z => n951);
   U890 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n952, Z => n1255);
   U891 : MUXB2DL port map( A0 => b(23), A1 => b(22), SL => n1539, Z => n952);
   U892 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n953, Z => n1256);
   U893 : MUXB2DL port map( A0 => b(22), A1 => b(21), SL => n1539, Z => n953);
   U894 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n954, Z => n1257);
   U895 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n1539, Z => n954);
   U896 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n955, Z => n1258);
   U897 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n1539, Z => n955);
   U898 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n956, Z => n1259);
   U899 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n1539, Z => n956);
   U900 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n957, Z => n1260);
   U901 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n1539, Z => n957);
   U902 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n958, Z => n1261);
   U903 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n1539, Z => n958);
   U904 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n959, Z => n1262);
   U905 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n1539, Z => n959);
   U906 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n960, Z => n1263);
   U907 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n1539, Z => n960);
   U908 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n961, Z => n1264);
   U909 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n1539, Z => n961);
   U910 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n962, Z => n1265);
   U911 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n1539, Z => n962);
   U912 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n963, Z => n1266);
   U913 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n1539, Z => n963);
   U914 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n964, Z => n1267);
   U915 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n1539, Z => n964);
   U916 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n965, Z => n1268);
   U917 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n1539, Z => n965);
   U918 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n966, Z => n1269);
   U919 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n1539, Z => n966);
   U920 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n967, Z => n1270);
   U921 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n1539, Z => n967);
   U922 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n968, Z => n1271);
   U923 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n1539, Z => n968);
   U924 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n969, Z => n1272);
   U925 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n1539, Z => n969);
   U926 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n970, Z => n1273);
   U927 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n1539, Z => n970);
   U928 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n971, Z => n1274);
   U929 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n1539, Z => n971);
   U930 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n972, Z => n1275);
   U931 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n1539, Z => n972);
   U932 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n973, Z => n1276);
   U933 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n1539, Z => n973);
   U934 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n974, Z => n1277);
   U935 : MUXB2DL port map( A0 => b(1), A1 => b(0), SL => n1539, Z => n974);
   U936 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n975, Z => n1278);
   U937 : NAN2M1D1 port map( A1 => n1539, A2 => b(0), Z => n975);
   U938 : NOR2M1D1 port map( A1 => n1518, A2 => n22, Z => n1094);
   U939 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n976, Z => n1279);
   U940 : MUXB2DL port map( A0 => b(27), A1 => b(26), SL => n1541, Z => n976);
   U941 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n977, Z => n1280);
   U942 : MUXB2DL port map( A0 => b(26), A1 => b(25), SL => n1541, Z => n977);
   U943 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n978, Z => n1281);
   U944 : MUXB2DL port map( A0 => b(25), A1 => b(24), SL => n1541, Z => n978);
   U945 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n979, Z => n1282);
   U946 : MUXB2DL port map( A0 => b(24), A1 => b(23), SL => n1541, Z => n979);
   U947 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n980, Z => n1283);
   U948 : MUXB2DL port map( A0 => b(23), A1 => b(22), SL => n1541, Z => n980);
   U949 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n981, Z => n1284);
   U950 : MUXB2DL port map( A0 => b(22), A1 => b(21), SL => n1541, Z => n981);
   U951 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n982, Z => n1285);
   U952 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n1541, Z => n982);
   U953 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n983, Z => n1286);
   U954 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n1541, Z => n983);
   U955 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n984, Z => n1287);
   U956 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n1541, Z => n984);
   U957 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n985, Z => n1288);
   U958 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n1541, Z => n985);
   U959 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n986, Z => n1289);
   U960 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n1541, Z => n986);
   U961 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n987, Z => n1290);
   U962 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n1541, Z => n987);
   U963 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n988, Z => n1291);
   U964 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n1541, Z => n988);
   U965 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n989, Z => n1292);
   U966 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n1541, Z => n989);
   U967 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n990, Z => n1293);
   U968 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n1541, Z => n990);
   U969 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n991, Z => n1294);
   U970 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n1541, Z => n991);
   U971 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n992, Z => n1295);
   U972 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n1541, Z => n992);
   U973 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n993, Z => n1296);
   U974 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n1541, Z => n993);
   U975 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n994, Z => n1297);
   U976 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n1541, Z => n994);
   U977 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n995, Z => n1298);
   U978 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n1541, Z => n995);
   U979 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n996, Z => n1299);
   U980 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n1541, Z => n996);
   U981 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n997, Z => n1300);
   U982 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n1541, Z => n997);
   U983 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n998, Z => n1301);
   U984 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n1541, Z => n998);
   U985 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n999, Z => n1302);
   U986 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n1541, Z => n999);
   U987 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n1000, Z => n1303);
   U988 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n1541, Z => n1000);
   U989 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n1001, Z => n1304);
   U990 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n1541, Z => n1001);
   U991 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n1002, Z => n1305);
   U992 : MUXB2DL port map( A0 => b(1), A1 => n1543, SL => n1541, Z => n1002);
   U993 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n1003, Z => n1306);
   U994 : NAN2M1D1 port map( A1 => n1541, A2 => b(0), Z => n1003);
   U995 : NOR2M1D1 port map( A1 => n1517, A2 => n14, Z => n1095);
   U996 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1004, Z => n1307);
   U997 : MUXB2DL port map( A0 => b(29), A1 => b(28), SL => n1542, Z => n1004);
   U998 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1005, Z => n1308);
   U999 : MUXB2DL port map( A0 => b(28), A1 => b(27), SL => n1542, Z => n1005);
   U1000 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1006, Z => n1309);
   U1001 : MUXB2DL port map( A0 => b(27), A1 => b(26), SL => n1542, Z => n1006)
                           ;
   U1002 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1007, Z => n1310);
   U1003 : MUXB2DL port map( A0 => b(26), A1 => b(25), SL => n1542, Z => n1007)
                           ;
   U1004 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1008, Z => n1311);
   U1005 : MUXB2DL port map( A0 => b(25), A1 => b(24), SL => n1542, Z => n1008)
                           ;
   U1006 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1009, Z => n1312);
   U1007 : MUXB2DL port map( A0 => b(24), A1 => b(23), SL => n1542, Z => n1009)
                           ;
   U1008 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1010, Z => n1313);
   U1009 : MUXB2DL port map( A0 => b(23), A1 => b(22), SL => n1542, Z => n1010)
                           ;
   U1010 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1011, Z => n1314);
   U1011 : MUXB2DL port map( A0 => b(22), A1 => b(21), SL => n1542, Z => n1011)
                           ;
   U1012 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1012, Z => n1315);
   U1013 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n1542, Z => n1012)
                           ;
   U1014 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1013, Z => n1316);
   U1015 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n1542, Z => n1013)
                           ;
   U1016 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1014, Z => n1317);
   U1017 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n1542, Z => n1014)
                           ;
   U1018 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1015, Z => n1318);
   U1019 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n1542, Z => n1015)
                           ;
   U1020 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1016, Z => n1319);
   U1021 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n1542, Z => n1016)
                           ;
   U1022 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1017, Z => n1320);
   U1023 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n1542, Z => n1017)
                           ;
   U1024 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1018, Z => n1321);
   U1025 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n1542, Z => n1018)
                           ;
   U1026 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1019, Z => n1322);
   U1027 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n1542, Z => n1019)
                           ;
   U1028 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1020, Z => n1323);
   U1029 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n1542, Z => n1020)
                           ;
   U1030 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1021, Z => n1324);
   U1031 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n1542, Z => n1021)
                           ;
   U1032 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1022, Z => n1325);
   U1033 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n1542, Z => n1022)
                           ;
   U1034 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1023, Z => n1326);
   U1035 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n1542, Z => n1023);
   U1036 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1024, Z => n1327);
   U1037 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n1542, Z => n1024);
   U1038 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1025, Z => n1328);
   U1039 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n1542, Z => n1025);
   U1040 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1026, Z => n1329);
   U1041 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n1542, Z => n1026);
   U1042 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1027, Z => n1330);
   U1043 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n1542, Z => n1027);
   U1044 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1028, Z => n1331);
   U1045 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n1542, Z => n1028);
   U1046 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1029, Z => n1332);
   U1047 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n1542, Z => n1029);
   U1048 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1030, Z => n1333);
   U1049 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n1542, Z => n1030);
   U1050 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1031, Z => n1334);
   U1051 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n1542, Z => n1031);
   U1052 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1032, Z => n1335);
   U1053 : MUXB2DL port map( A0 => b(1), A1 => n1543, SL => n1542, Z => n1032);
   U1054 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1033, Z => n1336);
   U1055 : NAN2M1D1 port map( A1 => n1542, A2 => b(0), Z => n1033);
   U1056 : NOR2M1D1 port map( A1 => n3, A2 => n6, Z => n1096);
   U1057 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1034, Z => n1337);
   U1058 : MUXB2DL port map( A0 => b(31), A1 => b(30), SL => n8, Z => n1034);
   U1059 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1035, Z => n1338);
   U1060 : MUXB2DL port map( A0 => b(30), A1 => b(29), SL => n8, Z => n1035);
   U1061 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1036, Z => n1339);
   U1062 : MUXB2DL port map( A0 => b(29), A1 => b(28), SL => n8, Z => n1036);
   U1063 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1037, Z => n1340);
   U1064 : MUXB2DL port map( A0 => b(28), A1 => b(27), SL => n8, Z => n1037);
   U1065 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1038, Z => n1341);
   U1066 : MUXB2DL port map( A0 => b(27), A1 => b(26), SL => n8, Z => n1038);
   U1067 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1039, Z => n1342);
   U1068 : MUXB2DL port map( A0 => b(26), A1 => b(25), SL => n8, Z => n1039);
   U1069 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1040, Z => n1343);
   U1070 : MUXB2DL port map( A0 => b(25), A1 => b(24), SL => n8, Z => n1040);
   U1071 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1041, Z => n1344);
   U1072 : MUXB2DL port map( A0 => b(24), A1 => b(23), SL => n8, Z => n1041);
   U1073 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1042, Z => n1345);
   U1074 : MUXB2DL port map( A0 => b(23), A1 => b(22), SL => n8, Z => n1042);
   U1075 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1043, Z => n1346);
   U1076 : MUXB2DL port map( A0 => b(22), A1 => b(21), SL => n8, Z => n1043);
   U1077 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1044, Z => n1347);
   U1078 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n8, Z => n1044);
   U1079 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1045, Z => n1348);
   U1080 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n8, Z => n1045);
   U1081 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1046, Z => n1349);
   U1082 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n8, Z => n1046);
   U1083 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1047, Z => n1350);
   U1084 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n8, Z => n1047);
   U1085 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1048, Z => n1351);
   U1086 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n8, Z => n1048);
   U1087 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1049, Z => n1352);
   U1088 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n8, Z => n1049);
   U1089 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1050, Z => n1353);
   U1090 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n8, Z => n1050);
   U1091 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1051, Z => n1354);
   U1092 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n8, Z => n1051);
   U1093 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1052, Z => n1355);
   U1094 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n8, Z => n1052);
   U1095 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1053, Z => n1356);
   U1096 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n8, Z => n1053);
   U1097 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1054, Z => n1357);
   U1098 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n8, Z => n1054);
   U1099 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1055, Z => n1358);
   U1100 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n8, Z => n1055);
   U1101 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1056, Z => n1359);
   U1102 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n8, Z => n1056);
   U1103 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1057, Z => n1360);
   U1104 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n8, Z => n1057);
   U1105 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1058, Z => n1361);
   U1106 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n8, Z => n1058);
   U1107 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1059, Z => n1362);
   U1108 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n8, Z => n1059);
   U1109 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1060, Z => n1363);
   U1110 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n8, Z => n1060);
   U1111 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1061, Z => n1364);
   U1112 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n8, Z => n1061);
   U1113 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1062, Z => n1365);
   U1114 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n8, Z => n1062);
   U1115 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1063, Z => n1366);
   U1116 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n8, Z => n1063);
   U1117 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1064, Z => n1367);
   U1118 : MUXB2DL port map( A0 => b(1), A1 => n1543, SL => n8, Z => n1064);
   U1119 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1065, Z => n1368);
   U1120 : NAN2M1D1 port map( A1 => n8, A2 => n1543, Z => n1065);
   U1121 : OAI21D1 port map( A1 => a(29), A2 => a(30), B => n1066, Z => n104);
   U1123 : EXNOR2D1 port map( A1 => a(29), A2 => a(30), Z => n106);
   U1125 : OAI21D1 port map( A1 => a(27), A2 => a(28), B => n1067, Z => n99);
   U1127 : EXNOR2D1 port map( A1 => a(27), A2 => a(28), Z => n103);
   U1129 : OAI21D1 port map( A1 => a(25), A2 => a(26), B => n1068, Z => n94);
   U1131 : EXNOR2D1 port map( A1 => a(25), A2 => a(26), Z => n98);
   U1135 : EXNOR2D1 port map( A1 => a(23), A2 => a(24), Z => n93);
   U1186 : ADHALFDL port map( A => n1278, B => n1093, CO => n780, S => n781);
   U1187 : OAI21D1 port map( A1 => a(1), A2 => a(2), B => n1080, Z => n1517);
   U1188 : OAI21D1 port map( A1 => a(3), A2 => a(4), B => n1079, Z => n1518);
   U1189 : OAI21D1 port map( A1 => a(7), A2 => a(8), B => n1077, Z => n1519);
   U1190 : AND2D1 port map( A1 => n1522, A2 => n305, Z => product(0));
   U1191 : AO21D1 port map( A1 => n215, A2 => n187, B => n188, Z => n1521);
   U1192 : OR2D1 port map( A1 => n1368, A2 => n1096, Z => n1522);
   U1193 : OA21M20D1 port map( A1 => n1523, A2 => n197, B => n194, Z => n190);
   U1194 : INVD1 port map( A => n215, Z => n214);
   U1195 : INVD1 port map( A => n233, Z => n232);
   U1196 : NAN2D1 port map( A1 => n313, A2 => n231, Z => n162);
   U1197 : INVD1 port map( A => n242, Z => n241);
   U1198 : INVD1 port map( A => n255, Z => n254);
   U1199 : INVD1 port map( A => n230, Z => n313);
   U1200 : INVD1 port map( A => n231, Z => n229);
   U1201 : INVD1 port map( A => n264, Z => n263);
   U1202 : NAN2D1 port map( A1 => n223, A2 => n1528, Z => n216);
   U1203 : INVD1 port map( A => n221, Z => n219);
   U1204 : NAN2D1 port map( A1 => n1530, A2 => n1529, Z => n243);
   U1205 : INVD1 port map( A => n248, Z => n246);
   U1206 : NAN2D1 port map( A1 => n1524, A2 => n1527, Z => n265);
   U1207 : INVD1 port map( A => n270, Z => n268);
   U1208 : NOR2D1 port map( A1 => n258, A2 => n261, Z => n256);
   U1209 : NOR2D1 port map( A1 => n236, A2 => n239, Z => n234);
   U1210 : NOR2D1 port map( A1 => n189, A2 => n201, Z => n187);
   U1211 : INVD1 port map( A => n209, Z => n211);
   U1212 : INVD1 port map( A => n206, Z => n204);
   U1213 : INVD1 port map( A => n275, Z => n273);
   U1214 : OR2D1 port map( A1 => n553, A2 => n574, Z => n1523);
   U1215 : NAN2D1 port map( A1 => n1523, A2 => n1526, Z => n189);
   U1216 : INVD1 port map( A => n199, Z => n197);
   U1217 : INVD1 port map( A => n253, Z => n251);
   U1218 : NAN2D1 port map( A1 => n667, A2 => n682, Z => n231);
   U1219 : NOR2D1 port map( A1 => n225, A2 => n230, Z => n223);
   U1220 : NAN2D1 port map( A1 => n1525, A2 => n310, Z => n201);
   U1221 : NOR2D1 port map( A1 => n683, A2 => n696, Z => n236);
   U1222 : NAN2D1 port map( A1 => n553, A2 => n574, Z => n194);
   U1223 : INVD1 port map( A => n208, Z => n310);
   U1224 : NOR2D1 port map( A1 => n667, A2 => n682, Z => n230);
   U1225 : NAN2D1 port map( A1 => n683, A2 => n696, Z => n237);
   U1226 : NAN2D1 port map( A1 => n1523, A2 => n194, Z => n156);
   U1227 : NAN2D1 port map( A1 => n1526, A2 => n199, Z => n157);
   U1228 : NAN2D1 port map( A1 => n1525, A2 => n206, Z => n158);
   U1229 : NAN2D1 port map( A1 => n310, A2 => n209, Z => n159);
   U1230 : NAN2D1 port map( A1 => n312, A2 => n226, Z => n161);
   U1231 : INVD1 port map( A => n225, Z => n312);
   U1232 : NAN2D1 port map( A1 => n1528, A2 => n221, Z => n160);
   U1233 : NAN2D1 port map( A1 => n314, A2 => n237, Z => n163);
   U1234 : INVD1 port map( A => n236, Z => n314);
   U1235 : NAN2D1 port map( A1 => n1530, A2 => n248, Z => n165);
   U1236 : NAN2D1 port map( A1 => n315, A2 => n240, Z => n164);
   U1237 : INVD1 port map( A => n239, Z => n315);
   U1238 : NAN2D1 port map( A1 => n1529, A2 => n253, Z => n166);
   U1239 : NAN2D1 port map( A1 => n318, A2 => n259, Z => n167);
   U1240 : INVD1 port map( A => n258, Z => n318);
   U1241 : NAN2D1 port map( A1 => n319, A2 => n262, Z => n168);
   U1242 : INVD1 port map( A => n261, Z => n319);
   U1243 : INVD1 port map( A => n277, Z => n276);
   U1244 : NAN2D1 port map( A1 => n1524, A2 => n270, Z => n169);
   U1245 : NAN2D1 port map( A1 => n1527, A2 => n275, Z => n170);
   U1246 : INVD1 port map( A => n286, Z => n285);
   U1247 : OR2D1 port map( A1 => n755, A2 => n762, Z => n1524);
   U1248 : NAN2D1 port map( A1 => n755, A2 => n762, Z => n270);
   U1249 : NOR2D1 port map( A1 => n280, A2 => n283, Z => n278);
   U1250 : OA21M20D1 port map( A1 => n1531, A2 => n294, B => n293, Z => n289);
   U1251 : NOR2D1 port map( A1 => n651, A2 => n666, Z => n225);
   U1252 : OA21M20D1 port map( A1 => n1532, A2 => n302, B => n301, Z => n297);
   U1253 : OR2D1 port map( A1 => n595, A2 => n614, Z => n1525);
   U1254 : NOR2D1 port map( A1 => n771, A2 => n776, Z => n280);
   U1255 : NOR2D1 port map( A1 => n745, A2 => n754, Z => n261);
   U1256 : NOR2D1 port map( A1 => n735, A2 => n744, Z => n258);
   U1257 : NAN2D1 port map( A1 => n763, A2 => n770, Z => n275);
   U1258 : OR2D1 port map( A1 => n575, A2 => n594, Z => n1526);
   U1259 : NAN2D1 port map( A1 => n575, A2 => n594, Z => n199);
   U1260 : NAN2D1 port map( A1 => n723, A2 => n734, Z => n253);
   U1261 : NAN2D1 port map( A1 => n651, A2 => n666, Z => n226);
   U1262 : OR2D1 port map( A1 => n763, A2 => n770, Z => n1527);
   U1263 : NAN2D1 port map( A1 => n595, A2 => n614, Z => n206);
   U1264 : OR2D1 port map( A1 => n633, A2 => n650, Z => n1528);
   U1265 : OR2D1 port map( A1 => n723, A2 => n734, Z => n1529);
   U1266 : NAN2D1 port map( A1 => n745, A2 => n754, Z => n262);
   U1267 : OR2D1 port map( A1 => n711, A2 => n722, Z => n1530);
   U1268 : NAN2D1 port map( A1 => n615, A2 => n632, Z => n209);
   U1269 : NAN2D1 port map( A1 => n771, A2 => n776, Z => n281);
   U1270 : NAN2D1 port map( A1 => n735, A2 => n744, Z => n259);
   U1271 : NOR2D1 port map( A1 => n615, A2 => n632, Z => n208);
   U1272 : NOR2D1 port map( A1 => n697, A2 => n710, Z => n239);
   U1273 : NAN2D1 port map( A1 => n711, A2 => n722, Z => n248);
   U1274 : NAN2D1 port map( A1 => n633, A2 => n650, Z => n221);
   U1275 : NAN2D1 port map( A1 => n697, A2 => n710, Z => n240);
   U1276 : NAN2D1 port map( A1 => n322, A2 => n281, Z => n171);
   U1277 : INVD1 port map( A => n280, Z => n322);
   U1278 : NAN2D1 port map( A1 => n323, A2 => n284, Z => n172);
   U1279 : INVD1 port map( A => n283, Z => n323);
   U1280 : NAN2D1 port map( A1 => n324, A2 => n288, Z => n173);
   U1281 : INVD1 port map( A => n287, Z => n324);
   U1282 : NAN2D1 port map( A1 => n1531, A2 => n293, Z => n174);
   U1283 : NAN2D1 port map( A1 => n326, A2 => n296, Z => n175);
   U1284 : INVD1 port map( A => n295, Z => n326);
   U1285 : NAN2D1 port map( A1 => n1532, A2 => n301, Z => n176);
   U1286 : OR2D1 port map( A1 => n787, A2 => n789, Z => n1531);
   U1287 : OR2D1 port map( A1 => n793, A2 => n1366, Z => n1532);
   U1288 : NOR2D1 port map( A1 => n777, A2 => n782, Z => n283);
   U1289 : NAN2D1 port map( A1 => n787, A2 => n789, Z => n293);
   U1290 : NAN2D1 port map( A1 => n793, A2 => n1366, Z => n301);
   U1291 : NAN2D1 port map( A1 => n777, A2 => n782, Z => n284);
   U1292 : NOR2D1 port map( A1 => n783, A2 => n786, Z => n287);
   U1293 : NOR2D1 port map( A1 => n791, A2 => n792, Z => n295);
   U1294 : NAN2D1 port map( A1 => n783, A2 => n786, Z => n288);
   U1295 : NAN2D1 port map( A1 => n791, A2 => n792, Z => n296);
   U1296 : NAN2D1 port map( A1 => n1368, A2 => n1096, Z => n305);
   U1297 : NOR2D1 port map( A1 => n303, A2 => n305, Z => n302);
   U1298 : INVD1 port map( A => n1533, Z => n1542);
   U1299 : EXOR2D1 port map( A1 => n178, A2 => n155, Z => product(31));
   U1300 : EXOR2D1 port map( A1 => n329, A2 => n344, Z => n155);
   U1301 : ADHALFDL port map( A => n1335, B => n1365, CO => n790, S => n791);
   U1302 : ADHALFDL port map( A => n1336, B => n1095, CO => n792, S => n793);
   U1303 : NOR2D1 port map( A1 => n1537, A2 => n30, Z => n1093);
   U1304 : INVD1 port map( A => n1535, Z => n1541);
   U1305 : ADHALFDL port map( A => n1331, B => n1361, CO => n774, S => n775);
   U1306 : INVD1 port map( A => n1534, Z => n1539);
   U1307 : ADHALFDL port map( A => n1252, B => n1092, CO => n768, S => n769);
   U1308 : INVD1 port map( A => n1536, Z => n1538);
   U1309 : ADHALFDL port map( A => n1333, B => n1363, CO => n784, S => n785);
   U1310 : ADHALFDL port map( A => n1306, B => n1094, CO => n788, S => n789);
   U1311 : INVD1 port map( A => n1537, Z => n1540);
   U1312 : ADHALFDL port map( A => n1206, B => n1090, CO => n732, S => n733);
   U1313 : ADHALFDL port map( A => n1168, B => n1088, CO => n680, S => n681);
   U1314 : ADHALFDL port map( A => n1152, B => n1087, CO => n648, S => n649);
   U1315 : ADHALFDL port map( A => n1228, B => n1091, CO => n752, S => n753);
   U1316 : ADHALFDL port map( A => n1186, B => n1089, CO => n708, S => n709);
   U1317 : ADHALFDL port map( A => n1138, B => n1086, CO => n612, S => n613);
   U1318 : INVD1 port map( A => n1367, Z => n303);
   U1319 : ADHALFDL port map( A => n1126, B => n1085, CO => n572, S => n573);
   U1320 : ADHALFDL port map( A => n1116, B => n1084, CO => n528, S => n529);
   U1321 : ADHALFDL port map( A => n1108, B => n1083, CO => n480, S => n481);
   U1322 : ADHALFDL port map( A => n1102, B => n1082, CO => n428, S => n429);
   U1323 : ADHALFDL port map( A => n1098, B => n1081, CO => n372, S => n373);
   U1324 : ADHALFDL port map( A => n1329, B => n1359, CO => n760, S => n761);
   U1325 : EXOR2D1 port map( A1 => a(1), A2 => a(2), Z => n1533);
   U1326 : ADHALFDL port map( A => n1323, B => n1353, CO => n694, S => n695);
   U1327 : EXOR2D1 port map( A1 => a(5), A2 => a(6), Z => n1534);
   U1328 : EXOR2D1 port map( A1 => a(3), A2 => a(4), Z => n1535);
   U1329 : EXOR2D1 port map( A1 => a(7), A2 => a(8), Z => n1536);
   U1330 : ADHALFDL port map( A => n1317, B => n1347, CO => n592, S => n593);
   U1331 : ADHALFDL port map( A => n1327, B => n1357, CO => n742, S => n743);
   U1332 : ADHALFDL port map( A => n1319, B => n1349, CO => n630, S => n631);
   U1333 : ADHALFDL port map( A => n1321, B => n1351, CO => n664, S => n665);
   U1334 : ADHALFDL port map( A => n1325, B => n1355, CO => n720, S => n721);
   U1335 : OA21D1 port map( A1 => a(5), A2 => a(6), B => n1078, Z => n1537);
   U1336 : INVD1 port map( A => a(3), Z => n1080);
   U1337 : EXNOR2D1 port map( A1 => a(11), A2 => a(12), Z => n56);
   U1338 : INVD1 port map( A => a(7), Z => n1078);
   U1339 : NAN2D1 port map( A1 => a(0), A2 => n6, Z => n3);
   U1340 : INVD1 port map( A => a(1), Z => n6);
   U1341 : INVD1 port map( A => a(9), Z => n1077);
   U1342 : EXNOR2D1 port map( A1 => a(13), A2 => a(14), Z => n63);
   U1343 : EXNOR2D1 port map( A1 => a(15), A2 => a(16), Z => n71);
   U1344 : INVD1 port map( A => a(5), Z => n1079);
   U1345 : EXNOR2D1 port map( A1 => a(9), A2 => a(10), Z => n48);
   U1346 : AO21D1 port map( A1 => a(1), A2 => a(2), B => n1080, Z => n14);
   U1347 : EXNOR2D1 port map( A1 => a(17), A2 => a(18), Z => n78);
   U1348 : INVD1 port map( A => n1544, Z => n1543);
   U1349 : AO21D1 port map( A1 => a(5), A2 => a(6), B => n1078, Z => n30);
   U1350 : INVD1 port map( A => a(0), Z => n8);
   U1351 : EXNOR2D1 port map( A1 => a(19), A2 => a(20), Z => n83);
   U1352 : AO21D1 port map( A1 => a(11), A2 => a(12), B => n1075, Z => n53);
   U1353 : INVD1 port map( A => a(13), Z => n1075);
   U1354 : ADHALFDL port map( A => n1315, B => n1345, CO => n550, S => n551);
   U1355 : AO21D1 port map( A1 => a(3), A2 => a(4), B => n1079, Z => n22);
   U1356 : AO21D1 port map( A1 => a(7), A2 => a(8), B => n1077, Z => n38);
   U1357 : OAI21D1 port map( A1 => a(11), A2 => a(12), B => n1075, Z => n50);
   U1358 : AO21D1 port map( A1 => a(13), A2 => a(14), B => n1074, Z => n61);
   U1359 : AO21D1 port map( A1 => a(15), A2 => a(16), B => n1073, Z => n69);
   U1360 : INVD1 port map( A => a(15), Z => n1074);
   U1361 : OAI21D1 port map( A1 => a(13), A2 => a(14), B => n1074, Z => n58);
   U1362 : INVD1 port map( A => a(17), Z => n1073);
   U1363 : OAI21D1 port map( A1 => a(15), A2 => a(16), B => n1073, Z => n66);
   U1364 : AO21D1 port map( A1 => a(9), A2 => a(10), B => n1076, Z => n45);
   U1365 : INVD1 port map( A => a(11), Z => n1076);
   U1366 : OAI21D1 port map( A1 => a(17), A2 => a(18), B => n1072, Z => n73);
   U1367 : INVD1 port map( A => a(19), Z => n1072);
   U1368 : OAI21D1 port map( A1 => a(9), A2 => a(10), B => n1076, Z => n42);
   U1369 : AO21D1 port map( A1 => a(17), A2 => a(18), B => n1072, Z => n76);
   U1370 : EXNOR2D1 port map( A1 => a(21), A2 => a(22), Z => n88);
   U1371 : OAI21D1 port map( A1 => a(19), A2 => a(20), B => n1071, Z => n79);
   U1372 : INVD1 port map( A => a(21), Z => n1071);
   U1373 : AO21D1 port map( A1 => a(19), A2 => a(20), B => n1071, Z => n81);
   U1374 : OAI21D1 port map( A1 => a(21), A2 => a(22), B => n1070, Z => n84);
   U1375 : INVD1 port map( A => a(23), Z => n1070);
   U1376 : AO21D1 port map( A1 => a(21), A2 => a(22), B => n1070, Z => n86);
   U1377 : ADHALFDL port map( A => n1313, B => n1343, CO => n504, S => n505);
   U1378 : ADHALFDL port map( A => n1311, B => n1341, CO => n454, S => n455);
   U1379 : OAI21D1 port map( A1 => a(23), A2 => a(24), B => n1069, Z => n89);
   U1380 : INVD1 port map( A => a(25), Z => n1069);
   U1381 : AO21D1 port map( A1 => a(23), A2 => a(24), B => n1069, Z => n91);
   U1382 : ADHALFDL port map( A => n1309, B => n1339, CO => n400, S => n401);
   U1383 : AO21D1 port map( A1 => a(25), A2 => a(26), B => n1068, Z => n96);
   U1384 : INVD1 port map( A => a(27), Z => n1068);
   U1385 : EXOR2D1 port map( A1 => n1307, A2 => n1337, Z => n343);
   U1386 : AO21D1 port map( A1 => a(27), A2 => a(28), B => n1067, Z => n101);
   U1387 : INVD1 port map( A => a(29), Z => n1067);
   U1388 : AO21D1 port map( A1 => a(29), A2 => a(30), B => n1066, Z => n105);
   U1389 : INVD1 port map( A => b(0), Z => n1544);
   U1390 : INVD1 port map( A => a(31), Z => n1066);

end hier_filter_none_5;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_gp_custom.all;

architecture hier_filter_none_5 of gp_custom_DW_mult_tc_6 is

   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AO21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component MUXB2DL
      port( A0, A1, SL : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component EXOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n6, n8, n14, n22, n30, n38, n42, n45, n48, n50, n53, n56, n58, 
      n61, n63, n66, n69, n71, n73, n76, n78, n79, n81, n83, n84, n86, n88, n89
      , n91, n93, n94, n96, n98, n99, n101, n103, n104, n105, n106, n155, n156,
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n178, n179, n180, n181, 
      n182, n183, n184, n185, n187, n188, n189, n190, n194, n195, n197, n199, 
      n200, n201, n202, n204, n206, n207, n208, n209, n211, n214, n215, n216, 
      n217, n219, n221, n222, n223, n224, n225, n226, n227, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n246, n248, n249, n251, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n268, n270, n271, n273, n275, 
      n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, 
      n288, n289, n293, n294, n295, n296, n297, n301, n302, n303, n305, n310, 
      n312, n313, n314, n315, n318, n319, n322, n323, n324, n326, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, 
      n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
      n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, 
      n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, 
      n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, 
      n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, 
      n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, 
      n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, 
      n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, 
      n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, 
      n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, 
      n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, 
      n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, 
      n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, 
      n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, 
      n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, 
      n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, 
      n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, 
      n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, 
      n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, 
      n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, 
      n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, 
      n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, 
      n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, 
      n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, 
      n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, 
      n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, 
      n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, 
      n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, 
      n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, 
      n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, 
      n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, 
      n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, 
      n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, 
      n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, 
      n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, 
      n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, 
      n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, 
      n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, 
      n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, 
      n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002
      , n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, 
      n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, 
      n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, 
      n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, 
      n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
      n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
      n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, 
      n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, 
      n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
      n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, 
      n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, 
      n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, 
      n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, 
      n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, 
      n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, 
      n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, 
      n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, 
      n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, 
      n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, 
      n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, 
      n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, 
      n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, 
      n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, 
      n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, 
      n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, 
      n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, 
      n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, 
      n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, 
      n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, 
      n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, 
      n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, 
      n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, 
      n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, 
      n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, 
      n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, 
      n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, 
      n1363, n1364, n1365, n1366, n1367, n1368, n1517, n1518, n1519, n1521, 
      n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, 
      n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, 
      n1542, n1543, n1544, n1545, n1546 : std_logic;

begin
   
   U125 : ADFULD1 port map( A => n345, B => n374, CI => n179, CO => n178, S => 
                           product(30));
   U126 : ADFULD1 port map( A => n375, B => n402, CI => n180, CO => n179, S => 
                           product(29));
   U127 : ADFULD1 port map( A => n403, B => n430, CI => n181, CO => n180, S => 
                           product(28));
   U128 : ADFULD1 port map( A => n431, B => n456, CI => n182, CO => n181, S => 
                           product(27));
   U129 : ADFULD1 port map( A => n457, B => n482, CI => n183, CO => n182, S => 
                           product(26));
   U130 : ADFULD1 port map( A => n483, B => n506, CI => n184, CO => n183, S => 
                           product(25));
   U131 : ADFULD1 port map( A => n507, B => n530, CI => n185, CO => n184, S => 
                           product(24));
   U132 : ADFULD1 port map( A => n531, B => n552, CI => n1521, CO => n185, S =>
                           product(23));
   U134 : EXOR2D1 port map( A1 => n195, A2 => n156, Z => product(22));
   U137 : OAI21D1 port map( A1 => n202, A2 => n189, B => n190, Z => n188);
   U146 : EXNOR2D1 port map( A1 => n200, A2 => n157, Z => product(21));
   U147 : AOI21D1 port map( A1 => n200, A2 => n1526, B => n197, Z => n195);
   U154 : EXNOR2D1 port map( A1 => n207, A2 => n158, Z => product(20));
   U155 : OAI21D1 port map( A1 => n214, A2 => n201, B => n202, Z => n200);
   U157 : AOI21D1 port map( A1 => n1525, A2 => n211, B => n204, Z => n202);
   U164 : EXOR2D1 port map( A1 => n214, A2 => n159, Z => product(19));
   U165 : OAI21D1 port map( A1 => n214, A2 => n208, B => n209, Z => n207);
   U174 : EXOR2D1 port map( A1 => n222, A2 => n160, Z => product(18));
   U176 : OAI21D1 port map( A1 => n233, A2 => n216, B => n217, Z => n215);
   U178 : AOI21D1 port map( A1 => n224, A2 => n1528, B => n219, Z => n217);
   U185 : EXOR2D1 port map( A1 => n227, A2 => n161, Z => product(17));
   U186 : AOI21D1 port map( A1 => n232, A2 => n223, B => n224, Z => n222);
   U188 : OAI21D1 port map( A1 => n225, A2 => n231, B => n226, Z => n224);
   U193 : EXNOR2D1 port map( A1 => n232, A2 => n162, Z => product(16));
   U194 : AOI21D1 port map( A1 => n232, A2 => n313, B => n229, Z => n227);
   U201 : EXNOR2D1 port map( A1 => n238, A2 => n163, Z => product(15));
   U203 : AOI21D1 port map( A1 => n242, A2 => n234, B => n235, Z => n233);
   U205 : OAI21D1 port map( A1 => n236, A2 => n240, B => n237, Z => n235);
   U210 : EXOR2D1 port map( A1 => n241, A2 => n164, Z => product(14));
   U211 : OAI21D1 port map( A1 => n241, A2 => n239, B => n240, Z => n238);
   U216 : EXOR2D1 port map( A1 => n249, A2 => n165, Z => product(13));
   U218 : OAI21D1 port map( A1 => n255, A2 => n243, B => n244, Z => n242);
   U220 : AOI21D1 port map( A1 => n1530, A2 => n251, B => n246, Z => n244);
   U227 : EXNOR2D1 port map( A1 => n254, A2 => n166, Z => product(12));
   U228 : AOI21D1 port map( A1 => n254, A2 => n1529, B => n251, Z => n249);
   U235 : EXNOR2D1 port map( A1 => n260, A2 => n167, Z => product(11));
   U237 : AOI21D1 port map( A1 => n256, A2 => n264, B => n257, Z => n255);
   U239 : OAI21D1 port map( A1 => n258, A2 => n262, B => n259, Z => n257);
   U244 : EXOR2D1 port map( A1 => n263, A2 => n168, Z => product(10));
   U245 : OAI21D1 port map( A1 => n263, A2 => n261, B => n262, Z => n260);
   U250 : EXOR2D1 port map( A1 => n271, A2 => n169, Z => product(9));
   U252 : OAI21D1 port map( A1 => n265, A2 => n277, B => n266, Z => n264);
   U254 : AOI21D1 port map( A1 => n1524, A2 => n273, B => n268, Z => n266);
   U261 : EXNOR2D1 port map( A1 => n276, A2 => n170, Z => product(8));
   U262 : AOI21D1 port map( A1 => n276, A2 => n1527, B => n273, Z => n271);
   U269 : EXNOR2D1 port map( A1 => n282, A2 => n171, Z => product(7));
   U271 : AOI21D1 port map( A1 => n278, A2 => n286, B => n279, Z => n277);
   U273 : OAI21D1 port map( A1 => n280, A2 => n284, B => n281, Z => n279);
   U278 : EXOR2D1 port map( A1 => n172, A2 => n285, Z => product(6));
   U279 : OAI21D1 port map( A1 => n285, A2 => n283, B => n284, Z => n282);
   U284 : EXOR2D1 port map( A1 => n173, A2 => n289, Z => product(5));
   U286 : OAI21D1 port map( A1 => n289, A2 => n287, B => n288, Z => n286);
   U291 : EXNOR2D1 port map( A1 => n174, A2 => n294, Z => product(4));
   U299 : EXOR2D1 port map( A1 => n297, A2 => n175, Z => product(3));
   U300 : OAI21D1 port map( A1 => n297, A2 => n295, B => n296, Z => n294);
   U305 : EXNOR2D1 port map( A1 => n176, A2 => n302, Z => product(2));
   U313 : EXOR2D1 port map( A1 => n303, A2 => n305, Z => product(1));
   U321 : EXOR3D1 port map( A1 => n346, A2 => n331, A3 => n330, Z => n329);
   U322 : EXOR3D1 port map( A1 => n332, A2 => n350, A3 => n348, Z => n330);
   U323 : EXOR3D1 port map( A1 => n352, A2 => n334, A3 => n333, Z => n331);
   U324 : EXOR3D1 port map( A1 => n354, A2 => n356, A3 => n335, Z => n332);
   U325 : EXOR3D1 port map( A1 => n337, A2 => n358, A3 => n336, Z => n333);
   U326 : EXOR3D1 port map( A1 => n339, A2 => n340, A3 => n360, Z => n334);
   U327 : EXOR3D1 port map( A1 => n342, A2 => n338, A3 => n341, Z => n335);
   U328 : EXOR3D1 port map( A1 => n366, A2 => n343, A3 => n362, Z => n336);
   U329 : EXOR3D1 port map( A1 => n368, A2 => n370, A3 => n364, Z => n337);
   U330 : EXOR3D1 port map( A1 => n1187, A2 => n1169, A3 => n372, Z => n338);
   U331 : EXOR3D1 port map( A1 => n1139, A2 => n1229, A3 => n1153, Z => n339);
   U332 : EXOR3D1 port map( A1 => n1103, A2 => n1117, A3 => n1109, Z => n340);
   U333 : EXOR3D1 port map( A1 => n1253, A2 => n1127, A3 => n1099, Z => n341);
   U334 : EXOR3D1 port map( A1 => n1097, A2 => n1279, A3 => n1207, Z => n342);
   U336 : ADFULD1 port map( A => n376, B => n349, CI => n347, CO => n344, S => 
                           n345);
   U337 : ADFULD1 port map( A => n351, B => n353, CI => n378, CO => n346, S => 
                           n347);
   U338 : ADFULD1 port map( A => n382, B => n355, CI => n380, CO => n348, S => 
                           n349);
   U339 : ADFULD1 port map( A => n359, B => n384, CI => n357, CO => n350, S => 
                           n351);
   U340 : ADFULD1 port map( A => n361, B => n388, CI => n386, CO => n352, S => 
                           n353);
   U341 : ADFULD1 port map( A => n365, B => n363, CI => n390, CO => n354, S => 
                           n355);
   U342 : ADFULD1 port map( A => n369, B => n371, CI => n367, CO => n356, S => 
                           n357);
   U343 : ADFULD1 port map( A => n398, B => n394, CI => n396, CO => n358, S => 
                           n359);
   U344 : ADFULD1 port map( A => n373, B => n400, CI => n392, CO => n360, S => 
                           n361);
   U345 : ADFULD1 port map( A => n1170, B => n1118, CI => n1140, CO => n362, S 
                           => n363);
   U346 : ADFULD1 port map( A => n1104, B => n1188, CI => n1110, CO => n364, S 
                           => n365);
   U347 : ADFULD1 port map( A => n1254, B => n1128, CI => n1230, CO => n366, S 
                           => n367);
   U348 : ADFULD1 port map( A => n1280, B => n1154, CI => n1208, CO => n368, S 
                           => n369);
   U349 : ADFULD1 port map( A => n1100, B => n1338, CI => n1308, CO => n370, S 
                           => n371);
   U351 : ADFULD1 port map( A => n404, B => n379, CI => n377, CO => n374, S => 
                           n375);
   U352 : ADFULD1 port map( A => n381, B => n408, CI => n406, CO => n376, S => 
                           n377);
   U353 : ADFULD1 port map( A => n410, B => n385, CI => n383, CO => n378, S => 
                           n379);
   U354 : ADFULD1 port map( A => n412, B => n389, CI => n387, CO => n380, S => 
                           n381);
   U355 : ADFULD1 port map( A => n391, B => n416, CI => n414, CO => n382, S => 
                           n383);
   U356 : ADFULD1 port map( A => n395, B => n397, CI => n399, CO => n384, S => 
                           n385);
   U357 : ADFULD1 port map( A => n418, B => n422, CI => n393, CO => n386, S => 
                           n387);
   U358 : ADFULD1 port map( A => n424, B => n426, CI => n420, CO => n388, S => 
                           n389);
   U359 : ADFULD1 port map( A => n428, B => n1171, CI => n401, CO => n390, S =>
                           n391);
   U360 : ADFULD1 port map( A => n1129, B => n1189, CI => n1141, CO => n392, S 
                           => n393);
   U361 : ADFULD1 port map( A => n1231, B => n1111, CI => n1105, CO => n394, S 
                           => n395);
   U362 : ADFULD1 port map( A => n1255, B => n1119, CI => n1101, CO => n396, S 
                           => n397);
   U363 : ADFULD1 port map( A => n1281, B => n1155, CI => n1209, CO => n398, S 
                           => n399);
   U365 : ADFULD1 port map( A => n432, B => n407, CI => n405, CO => n402, S => 
                           n403);
   U366 : ADFULD1 port map( A => n409, B => n436, CI => n434, CO => n404, S => 
                           n405);
   U367 : ADFULD1 port map( A => n438, B => n413, CI => n411, CO => n406, S => 
                           n407);
   U368 : ADFULD1 port map( A => n440, B => n417, CI => n415, CO => n408, S => 
                           n409);
   U369 : ADFULD1 port map( A => n444, B => n419, CI => n442, CO => n410, S => 
                           n411);
   U370 : ADFULD1 port map( A => n421, B => n423, CI => n425, CO => n412, S => 
                           n413);
   U371 : ADFULD1 port map( A => n448, B => n446, CI => n427, CO => n414, S => 
                           n415);
   U372 : ADFULD1 port map( A => n452, B => n429, CI => n450, CO => n416, S => 
                           n417);
   U373 : ADFULD1 port map( A => n1232, B => n1190, CI => n454, CO => n418, S 
                           => n419);
   U374 : ADFULD1 port map( A => n1142, B => n1256, CI => n1172, CO => n420, S 
                           => n421);
   U375 : ADFULD1 port map( A => n1112, B => n1130, CI => n1120, CO => n422, S 
                           => n423);
   U376 : ADFULD1 port map( A => n1282, B => n1156, CI => n1210, CO => n424, S 
                           => n425);
   U377 : ADFULD1 port map( A => n1106, B => n1340, CI => n1310, CO => n426, S 
                           => n427);
   U379 : ADFULD1 port map( A => n458, B => n435, CI => n433, CO => n430, S => 
                           n431);
   U380 : ADFULD1 port map( A => n437, B => n439, CI => n460, CO => n432, S => 
                           n433);
   U381 : ADFULD1 port map( A => n441, B => n464, CI => n462, CO => n434, S => 
                           n435);
   U382 : ADFULD1 port map( A => n466, B => n445, CI => n443, CO => n436, S => 
                           n437);
   U383 : ADFULD1 port map( A => n449, B => n451, CI => n468, CO => n438, S => 
                           n439);
   U384 : ADFULD1 port map( A => n453, B => n447, CI => n470, CO => n440, S => 
                           n441);
   U385 : ADFULD1 port map( A => n474, B => n472, CI => n476, CO => n442, S => 
                           n443);
   U386 : ADFULD1 port map( A => n455, B => n480, CI => n478, CO => n444, S => 
                           n445);
   U387 : ADFULD1 port map( A => n1131, B => n1191, CI => n1173, CO => n446, S 
                           => n447);
   U388 : ADFULD1 port map( A => n1113, B => n1233, CI => n1121, CO => n448, S 
                           => n449);
   U389 : ADFULD1 port map( A => n1283, B => n1143, CI => n1257, CO => n450, S 
                           => n451);
   U390 : ADFULD1 port map( A => n1107, B => n1157, CI => n1211, CO => n452, S 
                           => n453);
   U392 : ADFULD1 port map( A => n484, B => n461, CI => n459, CO => n456, S => 
                           n457);
   U393 : ADFULD1 port map( A => n486, B => n488, CI => n463, CO => n458, S => 
                           n459);
   U394 : ADFULD1 port map( A => n467, B => n469, CI => n465, CO => n460, S => 
                           n461);
   U395 : ADFULD1 port map( A => n492, B => n494, CI => n490, CO => n462, S => 
                           n463);
   U396 : ADFULD1 port map( A => n475, B => n477, CI => n471, CO => n464, S => 
                           n465);
   U397 : ADFULD1 port map( A => n479, B => n500, CI => n473, CO => n466, S => 
                           n467);
   U398 : ADFULD1 port map( A => n498, B => n502, CI => n496, CO => n468, S => 
                           n469);
   U399 : ADFULD1 port map( A => n504, B => n1192, CI => n481, CO => n470, S =>
                           n471);
   U400 : ADFULD1 port map( A => n1144, B => n1234, CI => n1158, CO => n472, S 
                           => n473);
   U401 : ADFULD1 port map( A => n1258, B => n1132, CI => n1122, CO => n474, S 
                           => n475);
   U402 : ADFULD1 port map( A => n1284, B => n1174, CI => n1212, CO => n476, S 
                           => n477);
   U403 : ADFULD1 port map( A => n1114, B => n1342, CI => n1312, CO => n478, S 
                           => n479);
   U405 : ADFULD1 port map( A => n508, B => n487, CI => n485, CO => n482, S => 
                           n483);
   U406 : ADFULD1 port map( A => n510, B => n512, CI => n489, CO => n484, S => 
                           n485);
   U407 : ADFULD1 port map( A => n493, B => n514, CI => n491, CO => n486, S => 
                           n487);
   U408 : ADFULD1 port map( A => n516, B => n518, CI => n495, CO => n488, S => 
                           n489);
   U409 : ADFULD1 port map( A => n501, B => n503, CI => n497, CO => n490, S => 
                           n491);
   U410 : ADFULD1 port map( A => n522, B => n524, CI => n499, CO => n492, S => 
                           n493);
   U411 : ADFULD1 port map( A => n526, B => n505, CI => n520, CO => n494, S => 
                           n495);
   U412 : ADFULD1 port map( A => n1235, B => n1259, CI => n528, CO => n496, S 
                           => n497);
   U413 : ADFULD1 port map( A => n1159, B => n1285, CI => n1193, CO => n498, S 
                           => n499);
   U414 : ADFULD1 port map( A => n1123, B => n1145, CI => n1133, CO => n500, S 
                           => n501);
   U415 : ADFULD1 port map( A => n1115, B => n1175, CI => n1213, CO => n502, S 
                           => n503);
   U417 : ADFULD1 port map( A => n532, B => n511, CI => n509, CO => n506, S => 
                           n507);
   U418 : ADFULD1 port map( A => n513, B => n536, CI => n534, CO => n508, S => 
                           n509);
   U419 : ADFULD1 port map( A => n517, B => n538, CI => n515, CO => n510, S => 
                           n511);
   U420 : ADFULD1 port map( A => n540, B => n542, CI => n519, CO => n512, S => 
                           n513);
   U421 : ADFULD1 port map( A => n525, B => n521, CI => n523, CO => n514, S => 
                           n515);
   U422 : ADFULD1 port map( A => n544, B => n546, CI => n527, CO => n516, S => 
                           n517);
   U423 : ADFULD1 port map( A => n529, B => n550, CI => n548, CO => n518, S => 
                           n519);
   U424 : ADFULD1 port map( A => n1194, B => n1260, CI => n1236, CO => n520, S 
                           => n521);
   U425 : ADFULD1 port map( A => n1134, B => n1286, CI => n1160, CO => n522, S 
                           => n523);
   U426 : ADFULD1 port map( A => n1124, B => n1176, CI => n1214, CO => n524, S 
                           => n525);
   U427 : ADFULD1 port map( A => n1146, B => n1344, CI => n1314, CO => n526, S 
                           => n527);
   U429 : ADFULD1 port map( A => n554, B => n535, CI => n533, CO => n530, S => 
                           n531);
   U430 : ADFULD1 port map( A => n556, B => n539, CI => n537, CO => n532, S => 
                           n533);
   U431 : ADFULD1 port map( A => n541, B => n560, CI => n558, CO => n534, S => 
                           n535);
   U432 : ADFULD1 port map( A => n562, B => n545, CI => n543, CO => n536, S => 
                           n537);
   U433 : ADFULD1 port map( A => n549, B => n564, CI => n547, CO => n538, S => 
                           n539);
   U434 : ADFULD1 port map( A => n566, B => n570, CI => n568, CO => n540, S => 
                           n541);
   U435 : ADFULD1 port map( A => n572, B => n1195, CI => n551, CO => n542, S =>
                           n543);
   U436 : ADFULD1 port map( A => n1135, B => n1237, CI => n1147, CO => n544, S 
                           => n545);
   U437 : ADFULD1 port map( A => n1287, B => n1161, CI => n1261, CO => n546, S 
                           => n547);
   U438 : ADFULD1 port map( A => n1125, B => n1177, CI => n1215, CO => n548, S 
                           => n549);
   U440 : ADFULD1 port map( A => n576, B => n557, CI => n555, CO => n552, S => 
                           n553);
   U441 : ADFULD1 port map( A => n559, B => n561, CI => n578, CO => n554, S => 
                           n555);
   U442 : ADFULD1 port map( A => n563, B => n582, CI => n580, CO => n556, S => 
                           n557);
   U443 : ADFULD1 port map( A => n565, B => n569, CI => n584, CO => n558, S => 
                           n559);
   U444 : ADFULD1 port map( A => n571, B => n586, CI => n567, CO => n560, S => 
                           n561);
   U445 : ADFULD1 port map( A => n590, B => n573, CI => n588, CO => n562, S => 
                           n563);
   U446 : ADFULD1 port map( A => n1196, B => n1238, CI => n592, CO => n564, S 
                           => n565);
   U447 : ADFULD1 port map( A => n1148, B => n1262, CI => n1162, CO => n566, S 
                           => n567);
   U448 : ADFULD1 port map( A => n1288, B => n1178, CI => n1216, CO => n568, S 
                           => n569);
   U449 : ADFULD1 port map( A => n1136, B => n1346, CI => n1316, CO => n570, S 
                           => n571);
   U451 : ADFULD1 port map( A => n596, B => n579, CI => n577, CO => n574, S => 
                           n575);
   U452 : ADFULD1 port map( A => n581, B => n583, CI => n598, CO => n576, S => 
                           n577);
   U453 : ADFULD1 port map( A => n585, B => n602, CI => n600, CO => n578, S => 
                           n579);
   U454 : ADFULD1 port map( A => n591, B => n589, CI => n604, CO => n580, S => 
                           n581);
   U455 : ADFULD1 port map( A => n606, B => n608, CI => n587, CO => n582, S => 
                           n583);
   U456 : ADFULD1 port map( A => n593, B => n612, CI => n610, CO => n584, S => 
                           n585);
   U457 : ADFULD1 port map( A => n1163, B => n1239, CI => n1197, CO => n586, S 
                           => n587);
   U458 : ADFULD1 port map( A => n1263, B => n1149, CI => n1137, CO => n588, S 
                           => n589);
   U459 : ADFULD1 port map( A => n1289, B => n1179, CI => n1217, CO => n590, S 
                           => n591);
   U461 : ADFULD1 port map( A => n616, B => n599, CI => n597, CO => n594, S => 
                           n595);
   U462 : ADFULD1 port map( A => n601, B => n603, CI => n618, CO => n596, S => 
                           n597);
   U463 : ADFULD1 port map( A => n622, B => n605, CI => n620, CO => n598, S => 
                           n599);
   U464 : ADFULD1 port map( A => n609, B => n611, CI => n607, CO => n600, S => 
                           n601);
   U465 : ADFULD1 port map( A => n626, B => n628, CI => n624, CO => n602, S => 
                           n603);
   U466 : ADFULD1 port map( A => n630, B => n1240, CI => n613, CO => n604, S =>
                           n605);
   U467 : ADFULD1 port map( A => n1150, B => n1264, CI => n1180, CO => n606, S 
                           => n607);
   U468 : ADFULD1 port map( A => n1290, B => n1198, CI => n1218, CO => n608, S 
                           => n609);
   U469 : ADFULD1 port map( A => n1164, B => n1348, CI => n1318, CO => n610, S 
                           => n611);
   U471 : ADFULD1 port map( A => n634, B => n619, CI => n617, CO => n614, S => 
                           n615);
   U472 : ADFULD1 port map( A => n621, B => n623, CI => n636, CO => n616, S => 
                           n617);
   U473 : ADFULD1 port map( A => n640, B => n625, CI => n638, CO => n618, S => 
                           n619);
   U474 : ADFULD1 port map( A => n627, B => n644, CI => n629, CO => n620, S => 
                           n621);
   U475 : ADFULD1 port map( A => n646, B => n631, CI => n642, CO => n622, S => 
                           n623);
   U476 : ADFULD1 port map( A => n1241, B => n1265, CI => n648, CO => n624, S 
                           => n625);
   U477 : ADFULD1 port map( A => n1291, B => n1181, CI => n1165, CO => n626, S 
                           => n627);
   U478 : ADFULD1 port map( A => n1151, B => n1199, CI => n1219, CO => n628, S 
                           => n629);
   U480 : ADFULD1 port map( A => n652, B => n637, CI => n635, CO => n632, S => 
                           n633);
   U481 : ADFULD1 port map( A => n639, B => n641, CI => n654, CO => n634, S => 
                           n635);
   U482 : ADFULD1 port map( A => n658, B => n645, CI => n656, CO => n636, S => 
                           n637);
   U483 : ADFULD1 port map( A => n647, B => n660, CI => n643, CO => n638, S => 
                           n639);
   U484 : ADFULD1 port map( A => n649, B => n664, CI => n662, CO => n640, S => 
                           n641);
   U485 : ADFULD1 port map( A => n1182, B => n1292, CI => n1242, CO => n642, S 
                           => n643);
   U486 : ADFULD1 port map( A => n1166, B => n1266, CI => n1220, CO => n644, S 
                           => n645);
   U487 : ADFULD1 port map( A => n1200, B => n1350, CI => n1320, CO => n646, S 
                           => n647);
   U489 : ADFULD1 port map( A => n668, B => n655, CI => n653, CO => n650, S => 
                           n651);
   U490 : ADFULD1 port map( A => n670, B => n659, CI => n657, CO => n652, S => 
                           n653);
   U491 : ADFULD1 port map( A => n663, B => n661, CI => n672, CO => n654, S => 
                           n655);
   U492 : ADFULD1 port map( A => n676, B => n678, CI => n674, CO => n656, S => 
                           n657);
   U493 : ADFULD1 port map( A => n680, B => n1267, CI => n665, CO => n658, S =>
                           n659);
   U494 : ADFULD1 port map( A => n1183, B => n1167, CI => n1243, CO => n660, S 
                           => n661);
   U495 : ADFULD1 port map( A => n1293, B => n1201, CI => n1221, CO => n662, S 
                           => n663);
   U497 : ADFULD1 port map( A => n684, B => n671, CI => n669, CO => n666, S => 
                           n667);
   U498 : ADFULD1 port map( A => n686, B => n688, CI => n673, CO => n668, S => 
                           n669);
   U499 : ADFULD1 port map( A => n677, B => n679, CI => n675, CO => n670, S => 
                           n671);
   U500 : ADFULD1 port map( A => n692, B => n681, CI => n690, CO => n672, S => 
                           n673);
   U501 : ADFULD1 port map( A => n1244, B => n1294, CI => n694, CO => n674, S 
                           => n675);
   U502 : ADFULD1 port map( A => n1184, B => n1268, CI => n1222, CO => n676, S 
                           => n677);
   U503 : ADFULD1 port map( A => n1202, B => n1352, CI => n1322, CO => n678, S 
                           => n679);
   U505 : ADFULD1 port map( A => n698, B => n687, CI => n685, CO => n682, S => 
                           n683);
   U506 : ADFULD1 port map( A => n700, B => n702, CI => n689, CO => n684, S => 
                           n685);
   U507 : ADFULD1 port map( A => n691, B => n704, CI => n693, CO => n686, S => 
                           n687);
   U508 : ADFULD1 port map( A => n695, B => n708, CI => n706, CO => n688, S => 
                           n689);
   U509 : ADFULD1 port map( A => n1185, B => n1245, CI => n1203, CO => n690, S 
                           => n691);
   U510 : ADFULD1 port map( A => n1295, B => n1269, CI => n1223, CO => n692, S 
                           => n693);
   U512 : ADFULD1 port map( A => n712, B => n701, CI => n699, CO => n696, S => 
                           n697);
   U513 : ADFULD1 port map( A => n703, B => n705, CI => n714, CO => n698, S => 
                           n699);
   U514 : ADFULD1 port map( A => n716, B => n718, CI => n707, CO => n700, S => 
                           n701);
   U515 : ADFULD1 port map( A => n720, B => n1270, CI => n709, CO => n702, S =>
                           n703);
   U516 : ADFULD1 port map( A => n1246, B => n1296, CI => n1224, CO => n704, S 
                           => n705);
   U517 : ADFULD1 port map( A => n1204, B => n1354, CI => n1324, CO => n706, S 
                           => n707);
   U519 : ADFULD1 port map( A => n724, B => n715, CI => n713, CO => n710, S => 
                           n711);
   U520 : ADFULD1 port map( A => n717, B => n719, CI => n726, CO => n712, S => 
                           n713);
   U521 : ADFULD1 port map( A => n730, B => n721, CI => n728, CO => n714, S => 
                           n715);
   U522 : ADFULD1 port map( A => n1205, B => n1247, CI => n732, CO => n716, S 
                           => n717);
   U523 : ADFULD1 port map( A => n1271, B => n1297, CI => n1225, CO => n718, S 
                           => n719);
   U525 : ADFULD1 port map( A => n736, B => n727, CI => n725, CO => n722, S => 
                           n723);
   U526 : ADFULD1 port map( A => n729, B => n731, CI => n738, CO => n724, S => 
                           n725);
   U527 : ADFULD1 port map( A => n733, B => n742, CI => n740, CO => n726, S => 
                           n727);
   U528 : ADFULD1 port map( A => n1272, B => n1298, CI => n1226, CO => n728, S 
                           => n729);
   U529 : ADFULD1 port map( A => n1248, B => n1356, CI => n1326, CO => n730, S 
                           => n731);
   U531 : ADFULD1 port map( A => n746, B => n739, CI => n737, CO => n734, S => 
                           n735);
   U532 : ADFULD1 port map( A => n748, B => n750, CI => n741, CO => n736, S => 
                           n737);
   U533 : ADFULD1 port map( A => n752, B => n1299, CI => n743, CO => n738, S =>
                           n739);
   U534 : ADFULD1 port map( A => n1273, B => n1249, CI => n1227, CO => n740, S 
                           => n741);
   U536 : ADFULD1 port map( A => n756, B => n749, CI => n747, CO => n744, S => 
                           n745);
   U537 : ADFULD1 port map( A => n758, B => n753, CI => n751, CO => n746, S => 
                           n747);
   U538 : ADFULD1 port map( A => n1274, B => n1300, CI => n760, CO => n748, S 
                           => n749);
   U539 : ADFULD1 port map( A => n1250, B => n1358, CI => n1328, CO => n750, S 
                           => n751);
   U541 : ADFULD1 port map( A => n764, B => n759, CI => n757, CO => n754, S => 
                           n755);
   U542 : ADFULD1 port map( A => n761, B => n768, CI => n766, CO => n756, S => 
                           n757);
   U543 : ADFULD1 port map( A => n1275, B => n1251, CI => n1301, CO => n758, S 
                           => n759);
   U545 : ADFULD1 port map( A => n767, B => n772, CI => n765, CO => n762, S => 
                           n763);
   U546 : ADFULD1 port map( A => n774, B => n1302, CI => n769, CO => n764, S =>
                           n765);
   U547 : ADFULD1 port map( A => n1276, B => n1360, CI => n1330, CO => n766, S 
                           => n767);
   U549 : ADFULD1 port map( A => n778, B => n775, CI => n773, CO => n770, S => 
                           n771);
   U550 : ADFULD1 port map( A => n1277, B => n1303, CI => n780, CO => n772, S 
                           => n773);
   U552 : ADFULD1 port map( A => n781, B => n784, CI => n779, CO => n776, S => 
                           n777);
   U553 : ADFULD1 port map( A => n1304, B => n1362, CI => n1332, CO => n778, S 
                           => n779);
   U555 : ADFULD1 port map( A => n788, B => n1305, CI => n785, CO => n782, S =>
                           n783);
   U557 : ADFULD1 port map( A => n1334, B => n1364, CI => n790, CO => n786, S 
                           => n787);
   U561 : NOR2M1D1 port map( A1 => n104, A2 => n105, Z => n1081);
   U562 : MUXB2DL port map( A0 => n104, A1 => n105, SL => n794, Z => n1097);
   U563 : MUXB2DL port map( A0 => b(1), A1 => b(0), SL => n106, Z => n794);
   U564 : MUXB2DL port map( A0 => n104, A1 => n105, SL => n795, Z => n1098);
   U565 : NAN2M1D1 port map( A1 => n106, A2 => b(0), Z => n795);
   U566 : NOR2M1D1 port map( A1 => n99, A2 => n101, Z => n1082);
   U567 : MUXB2DL port map( A0 => n99, A1 => n101, SL => n796, Z => n1099);
   U568 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n103, Z => n796);
   U569 : MUXB2DL port map( A0 => n99, A1 => n101, SL => n797, Z => n1100);
   U570 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n103, Z => n797);
   U571 : MUXB2DL port map( A0 => n99, A1 => n101, SL => n798, Z => n1101);
   U572 : MUXB2DL port map( A0 => b(1), A1 => b(0), SL => n103, Z => n798);
   U573 : MUXB2DL port map( A0 => n99, A1 => n101, SL => n799, Z => n1102);
   U574 : NAN2M1D1 port map( A1 => n103, A2 => b(0), Z => n799);
   U575 : NOR2M1D1 port map( A1 => n94, A2 => n96, Z => n1083);
   U576 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n800, Z => n1103);
   U577 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n98, Z => n800);
   U578 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n801, Z => n1104);
   U579 : MUXB2DL port map( A0 => b(4), A1 => n1543, SL => n98, Z => n801);
   U580 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n802, Z => n1105);
   U581 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n98, Z => n802);
   U582 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n803, Z => n1106);
   U583 : MUXB2DL port map( A0 => b(2), A1 => n1545, SL => n98, Z => n803);
   U584 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n804, Z => n1107);
   U585 : MUXB2DL port map( A0 => b(1), A1 => b(0), SL => n98, Z => n804);
   U586 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n805, Z => n1108);
   U587 : NAN2M1D1 port map( A1 => n98, A2 => b(0), Z => n805);
   U588 : NOR2M1D1 port map( A1 => n89, A2 => n91, Z => n1084);
   U589 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n806, Z => n1109);
   U590 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n93, Z => n806);
   U591 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n807, Z => n1110);
   U592 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n93, Z => n807);
   U593 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n808, Z => n1111);
   U594 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n93, Z => n808);
   U595 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n809, Z => n1112);
   U596 : MUXB2DL port map( A0 => b(4), A1 => n1543, SL => n93, Z => n809);
   U597 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n810, Z => n1113);
   U598 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n93, Z => n810);
   U599 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n811, Z => n1114);
   U600 : MUXB2DL port map( A0 => b(2), A1 => n1545, SL => n93, Z => n811);
   U601 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n812, Z => n1115);
   U602 : MUXB2DL port map( A0 => b(1), A1 => b(0), SL => n93, Z => n812);
   U603 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n813, Z => n1116);
   U604 : NAN2M1D1 port map( A1 => n93, A2 => b(0), Z => n813);
   U605 : NOR2M1D1 port map( A1 => n84, A2 => n86, Z => n1085);
   U606 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n814, Z => n1117);
   U607 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n88, Z => n814);
   U608 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n815, Z => n1118);
   U609 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n88, Z => n815);
   U610 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n816, Z => n1119);
   U611 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n88, Z => n816);
   U612 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n817, Z => n1120);
   U613 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n88, Z => n817);
   U614 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n818, Z => n1121);
   U615 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n88, Z => n818);
   U616 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n819, Z => n1122);
   U617 : MUXB2DL port map( A0 => b(4), A1 => n1543, SL => n88, Z => n819);
   U618 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n820, Z => n1123);
   U619 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n88, Z => n820);
   U620 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n821, Z => n1124);
   U621 : MUXB2DL port map( A0 => b(2), A1 => n1545, SL => n88, Z => n821);
   U622 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n822, Z => n1125);
   U623 : MUXB2DL port map( A0 => b(1), A1 => b(0), SL => n88, Z => n822);
   U624 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n823, Z => n1126);
   U625 : NAN2M1D1 port map( A1 => n88, A2 => b(0), Z => n823);
   U626 : NOR2M1D1 port map( A1 => n79, A2 => n81, Z => n1086);
   U627 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n824, Z => n1127);
   U628 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n83, Z => n824);
   U629 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n825, Z => n1128);
   U630 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n83, Z => n825);
   U631 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n826, Z => n1129);
   U632 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n83, Z => n826);
   U633 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n827, Z => n1130);
   U634 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n83, Z => n827);
   U635 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n828, Z => n1131);
   U636 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n83, Z => n828);
   U637 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n829, Z => n1132);
   U638 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n83, Z => n829);
   U639 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n830, Z => n1133);
   U640 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n83, Z => n830);
   U641 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n831, Z => n1134);
   U642 : MUXB2DL port map( A0 => b(4), A1 => n1543, SL => n83, Z => n831);
   U643 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n832, Z => n1135);
   U644 : MUXB2DL port map( A0 => n1543, A1 => b(2), SL => n83, Z => n832);
   U645 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n833, Z => n1136);
   U646 : MUXB2DL port map( A0 => b(2), A1 => n1545, SL => n83, Z => n833);
   U647 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n834, Z => n1137);
   U648 : MUXB2DL port map( A0 => b(1), A1 => b(0), SL => n83, Z => n834);
   U649 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n835, Z => n1138);
   U650 : NAN2M1D1 port map( A1 => n83, A2 => b(0), Z => n835);
   U651 : NOR2M1D1 port map( A1 => n73, A2 => n76, Z => n1087);
   U652 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n836, Z => n1139);
   U653 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n78, Z => n836);
   U654 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n837, Z => n1140);
   U655 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n78, Z => n837);
   U656 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n838, Z => n1141);
   U657 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n78, Z => n838);
   U658 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n839, Z => n1142);
   U659 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n78, Z => n839);
   U660 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n840, Z => n1143);
   U661 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n78, Z => n840);
   U662 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n841, Z => n1144);
   U663 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n78, Z => n841);
   U664 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n842, Z => n1145);
   U665 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n78, Z => n842);
   U666 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n843, Z => n1146);
   U667 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n78, Z => n843);
   U668 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n844, Z => n1147);
   U669 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n78, Z => n844);
   U670 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n845, Z => n1148);
   U671 : MUXB2DL port map( A0 => b(4), A1 => n1543, SL => n78, Z => n845);
   U672 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n846, Z => n1149);
   U673 : MUXB2DL port map( A0 => n1543, A1 => b(2), SL => n78, Z => n846);
   U674 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n847, Z => n1150);
   U675 : MUXB2DL port map( A0 => b(2), A1 => n1545, SL => n78, Z => n847);
   U676 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n848, Z => n1151);
   U677 : MUXB2DL port map( A0 => b(1), A1 => b(0), SL => n78, Z => n848);
   U678 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n849, Z => n1152);
   U679 : NAN2M1D1 port map( A1 => n78, A2 => b(0), Z => n849);
   U680 : NOR2M1D1 port map( A1 => n66, A2 => n69, Z => n1088);
   U681 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n850, Z => n1153);
   U682 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n71, Z => n850);
   U683 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n851, Z => n1154);
   U684 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n71, Z => n851);
   U685 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n852, Z => n1155);
   U686 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n71, Z => n852);
   U687 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n853, Z => n1156);
   U688 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n71, Z => n853);
   U689 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n854, Z => n1157);
   U690 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n71, Z => n854);
   U691 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n855, Z => n1158);
   U692 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n71, Z => n855);
   U693 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n856, Z => n1159);
   U694 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n71, Z => n856);
   U695 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n857, Z => n1160);
   U696 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n71, Z => n857);
   U697 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n858, Z => n1161);
   U698 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n71, Z => n858);
   U699 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n859, Z => n1162);
   U700 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n71, Z => n859);
   U701 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n860, Z => n1163);
   U702 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n71, Z => n860);
   U703 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n861, Z => n1164);
   U704 : MUXB2DL port map( A0 => b(4), A1 => n1543, SL => n71, Z => n861);
   U705 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n862, Z => n1165);
   U706 : MUXB2DL port map( A0 => n1543, A1 => b(2), SL => n71, Z => n862);
   U707 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n863, Z => n1166);
   U708 : MUXB2DL port map( A0 => b(2), A1 => n1545, SL => n71, Z => n863);
   U709 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n864, Z => n1167);
   U710 : MUXB2DL port map( A0 => b(1), A1 => b(0), SL => n71, Z => n864);
   U711 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n865, Z => n1168);
   U712 : NAN2M1D1 port map( A1 => n71, A2 => b(0), Z => n865);
   U713 : NOR2M1D1 port map( A1 => n58, A2 => n61, Z => n1089);
   U714 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n866, Z => n1169);
   U715 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n63, Z => n866);
   U716 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n867, Z => n1170);
   U717 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n63, Z => n867);
   U718 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n868, Z => n1171);
   U719 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n63, Z => n868);
   U720 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n869, Z => n1172);
   U721 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n63, Z => n869);
   U722 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n870, Z => n1173);
   U723 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n63, Z => n870);
   U724 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n871, Z => n1174);
   U725 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n63, Z => n871);
   U726 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n872, Z => n1175);
   U727 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n63, Z => n872);
   U728 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n873, Z => n1176);
   U729 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n63, Z => n873);
   U730 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n874, Z => n1177);
   U731 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n63, Z => n874);
   U732 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n875, Z => n1178);
   U733 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n63, Z => n875);
   U734 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n876, Z => n1179);
   U735 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n63, Z => n876);
   U736 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n877, Z => n1180);
   U737 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n63, Z => n877);
   U738 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n878, Z => n1181);
   U739 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n63, Z => n878);
   U740 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n879, Z => n1182);
   U741 : MUXB2DL port map( A0 => b(4), A1 => n1543, SL => n63, Z => n879);
   U742 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n880, Z => n1183);
   U743 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n63, Z => n880);
   U744 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n881, Z => n1184);
   U745 : MUXB2DL port map( A0 => b(2), A1 => n1545, SL => n63, Z => n881);
   U746 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n882, Z => n1185);
   U747 : MUXB2DL port map( A0 => n1545, A1 => b(0), SL => n63, Z => n882);
   U748 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n883, Z => n1186);
   U749 : NAN2M1D1 port map( A1 => n63, A2 => b(0), Z => n883);
   U750 : NOR2M1D1 port map( A1 => n50, A2 => n53, Z => n1090);
   U751 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n884, Z => n1187);
   U752 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n56, Z => n884);
   U753 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n885, Z => n1188);
   U754 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n56, Z => n885);
   U755 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n886, Z => n1189);
   U756 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n56, Z => n886);
   U757 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n887, Z => n1190);
   U758 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n56, Z => n887);
   U759 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n888, Z => n1191);
   U760 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n56, Z => n888);
   U761 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n889, Z => n1192);
   U762 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n56, Z => n889);
   U763 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n890, Z => n1193);
   U764 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n56, Z => n890);
   U765 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n891, Z => n1194);
   U766 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n56, Z => n891);
   U767 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n892, Z => n1195);
   U768 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n56, Z => n892);
   U769 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n893, Z => n1196);
   U770 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n56, Z => n893);
   U771 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n894, Z => n1197);
   U772 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n56, Z => n894);
   U773 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n895, Z => n1198);
   U774 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n56, Z => n895);
   U775 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n896, Z => n1199);
   U776 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n56, Z => n896);
   U777 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n897, Z => n1200);
   U778 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n56, Z => n897);
   U779 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n898, Z => n1201);
   U780 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n56, Z => n898);
   U781 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n899, Z => n1202);
   U782 : MUXB2DL port map( A0 => b(4), A1 => n1543, SL => n56, Z => n899);
   U783 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n900, Z => n1203);
   U784 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n56, Z => n900);
   U785 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n901, Z => n1204);
   U786 : MUXB2DL port map( A0 => b(2), A1 => n1545, SL => n56, Z => n901);
   U787 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n902, Z => n1205);
   U788 : MUXB2DL port map( A0 => n1545, A1 => b(0), SL => n56, Z => n902);
   U789 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n903, Z => n1206);
   U790 : NAN2M1D1 port map( A1 => n56, A2 => b(0), Z => n903);
   U791 : NOR2M1D1 port map( A1 => n42, A2 => n45, Z => n1091);
   U792 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n904, Z => n1207);
   U793 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n48, Z => n904);
   U794 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n905, Z => n1208);
   U795 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n48, Z => n905);
   U796 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n906, Z => n1209);
   U797 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n48, Z => n906);
   U798 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n907, Z => n1210);
   U799 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n48, Z => n907);
   U800 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n908, Z => n1211);
   U801 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n48, Z => n908);
   U802 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n909, Z => n1212);
   U803 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n48, Z => n909);
   U804 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n910, Z => n1213);
   U805 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n48, Z => n910);
   U806 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n911, Z => n1214);
   U807 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n48, Z => n911);
   U808 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n912, Z => n1215);
   U809 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n48, Z => n912);
   U810 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n913, Z => n1216);
   U811 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n48, Z => n913);
   U812 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n914, Z => n1217);
   U813 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n48, Z => n914);
   U814 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n915, Z => n1218);
   U815 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n48, Z => n915);
   U816 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n916, Z => n1219);
   U817 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n48, Z => n916);
   U818 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n917, Z => n1220);
   U819 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n48, Z => n917);
   U820 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n918, Z => n1221);
   U821 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n48, Z => n918);
   U822 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n919, Z => n1222);
   U823 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n48, Z => n919);
   U824 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n920, Z => n1223);
   U825 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n48, Z => n920);
   U826 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n921, Z => n1224);
   U827 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n48, Z => n921);
   U828 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n922, Z => n1225);
   U829 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n48, Z => n922);
   U830 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n923, Z => n1226);
   U831 : MUXB2DL port map( A0 => b(2), A1 => n1545, SL => n48, Z => n923);
   U832 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n924, Z => n1227);
   U833 : MUXB2DL port map( A0 => n1545, A1 => b(0), SL => n48, Z => n924);
   U834 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n925, Z => n1228);
   U835 : NAN2M1D1 port map( A1 => n48, A2 => b(0), Z => n925);
   U836 : NOR2M1D1 port map( A1 => n1519, A2 => n38, Z => n1092);
   U837 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n926, Z => n1229);
   U838 : MUXB2DL port map( A0 => b(23), A1 => b(22), SL => n1538, Z => n926);
   U839 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n927, Z => n1230);
   U840 : MUXB2DL port map( A0 => b(22), A1 => b(21), SL => n1538, Z => n927);
   U841 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n928, Z => n1231);
   U842 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n1538, Z => n928);
   U843 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n929, Z => n1232);
   U844 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n1538, Z => n929);
   U845 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n930, Z => n1233);
   U846 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n1538, Z => n930);
   U847 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n931, Z => n1234);
   U848 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n1538, Z => n931);
   U849 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n932, Z => n1235);
   U850 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n1538, Z => n932);
   U851 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n933, Z => n1236);
   U852 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n1538, Z => n933);
   U853 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n934, Z => n1237);
   U854 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n1538, Z => n934);
   U855 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n935, Z => n1238);
   U856 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n1538, Z => n935);
   U857 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n936, Z => n1239);
   U858 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n1538, Z => n936);
   U859 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n937, Z => n1240);
   U860 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n1538, Z => n937);
   U861 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n938, Z => n1241);
   U862 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n1538, Z => n938);
   U863 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n939, Z => n1242);
   U864 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n1538, Z => n939);
   U865 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n940, Z => n1243);
   U866 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n1538, Z => n940);
   U867 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n941, Z => n1244);
   U868 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n1538, Z => n941);
   U869 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n942, Z => n1245);
   U870 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n1538, Z => n942);
   U871 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n943, Z => n1246);
   U872 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n1538, Z => n943);
   U873 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n944, Z => n1247);
   U874 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n1538, Z => n944);
   U875 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n945, Z => n1248);
   U876 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n1538, Z => n945);
   U877 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n946, Z => n1249);
   U878 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n1538, Z => n946);
   U879 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n947, Z => n1250);
   U880 : MUXB2DL port map( A0 => b(2), A1 => n1545, SL => n1538, Z => n947);
   U881 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n948, Z => n1251);
   U882 : MUXB2DL port map( A0 => b(1), A1 => b(0), SL => n1538, Z => n948);
   U883 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n949, Z => n1252);
   U884 : NAN2M1D1 port map( A1 => n1538, A2 => b(0), Z => n949);
   U886 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n950, Z => n1253);
   U887 : MUXB2DL port map( A0 => b(25), A1 => b(24), SL => n1539, Z => n950);
   U888 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n951, Z => n1254);
   U889 : MUXB2DL port map( A0 => b(24), A1 => b(23), SL => n1539, Z => n951);
   U890 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n952, Z => n1255);
   U891 : MUXB2DL port map( A0 => b(23), A1 => b(22), SL => n1539, Z => n952);
   U892 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n953, Z => n1256);
   U893 : MUXB2DL port map( A0 => b(22), A1 => b(21), SL => n1539, Z => n953);
   U894 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n954, Z => n1257);
   U895 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n1539, Z => n954);
   U896 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n955, Z => n1258);
   U897 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n1539, Z => n955);
   U898 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n956, Z => n1259);
   U899 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n1539, Z => n956);
   U900 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n957, Z => n1260);
   U901 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n1539, Z => n957);
   U902 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n958, Z => n1261);
   U903 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n1539, Z => n958);
   U904 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n959, Z => n1262);
   U905 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n1539, Z => n959);
   U906 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n960, Z => n1263);
   U907 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n1539, Z => n960);
   U908 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n961, Z => n1264);
   U909 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n1539, Z => n961);
   U910 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n962, Z => n1265);
   U911 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n1539, Z => n962);
   U912 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n963, Z => n1266);
   U913 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n1539, Z => n963);
   U914 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n964, Z => n1267);
   U915 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n1539, Z => n964);
   U916 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n965, Z => n1268);
   U917 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n1539, Z => n965);
   U918 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n966, Z => n1269);
   U919 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n1539, Z => n966);
   U920 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n967, Z => n1270);
   U921 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n1539, Z => n967);
   U922 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n968, Z => n1271);
   U923 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n1539, Z => n968);
   U924 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n969, Z => n1272);
   U925 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n1539, Z => n969);
   U926 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n970, Z => n1273);
   U927 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n1539, Z => n970);
   U928 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n971, Z => n1274);
   U929 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n1539, Z => n971);
   U930 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n972, Z => n1275);
   U931 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n1539, Z => n972);
   U932 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n973, Z => n1276);
   U933 : MUXB2DL port map( A0 => b(2), A1 => n1545, SL => n1539, Z => n973);
   U934 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n974, Z => n1277);
   U935 : MUXB2DL port map( A0 => b(1), A1 => b(0), SL => n1539, Z => n974);
   U936 : MUXB2DL port map( A0 => n1540, A1 => n30, SL => n975, Z => n1278);
   U937 : NAN2M1D1 port map( A1 => n1539, A2 => b(0), Z => n975);
   U938 : NOR2M1D1 port map( A1 => n1518, A2 => n22, Z => n1094);
   U939 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n976, Z => n1279);
   U940 : MUXB2DL port map( A0 => b(27), A1 => b(26), SL => n1541, Z => n976);
   U941 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n977, Z => n1280);
   U942 : MUXB2DL port map( A0 => b(26), A1 => b(25), SL => n1541, Z => n977);
   U943 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n978, Z => n1281);
   U944 : MUXB2DL port map( A0 => b(25), A1 => b(24), SL => n1541, Z => n978);
   U945 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n979, Z => n1282);
   U946 : MUXB2DL port map( A0 => b(24), A1 => b(23), SL => n1541, Z => n979);
   U947 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n980, Z => n1283);
   U948 : MUXB2DL port map( A0 => b(23), A1 => b(22), SL => n1541, Z => n980);
   U949 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n981, Z => n1284);
   U950 : MUXB2DL port map( A0 => b(22), A1 => b(21), SL => n1541, Z => n981);
   U951 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n982, Z => n1285);
   U952 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n1541, Z => n982);
   U953 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n983, Z => n1286);
   U954 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n1541, Z => n983);
   U955 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n984, Z => n1287);
   U956 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n1541, Z => n984);
   U957 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n985, Z => n1288);
   U958 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n1541, Z => n985);
   U959 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n986, Z => n1289);
   U960 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n1541, Z => n986);
   U961 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n987, Z => n1290);
   U962 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n1541, Z => n987);
   U963 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n988, Z => n1291);
   U964 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n1541, Z => n988);
   U965 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n989, Z => n1292);
   U966 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n1541, Z => n989);
   U967 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n990, Z => n1293);
   U968 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n1541, Z => n990);
   U969 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n991, Z => n1294);
   U970 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n1541, Z => n991);
   U971 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n992, Z => n1295);
   U972 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n1541, Z => n992);
   U973 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n993, Z => n1296);
   U974 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n1541, Z => n993);
   U975 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n994, Z => n1297);
   U976 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n1541, Z => n994);
   U977 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n995, Z => n1298);
   U978 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n1541, Z => n995);
   U979 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n996, Z => n1299);
   U980 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n1541, Z => n996);
   U981 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n997, Z => n1300);
   U982 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n1541, Z => n997);
   U983 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n998, Z => n1301);
   U984 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n1541, Z => n998);
   U985 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n999, Z => n1302);
   U986 : MUXB2DL port map( A0 => b(4), A1 => n1543, SL => n1541, Z => n999);
   U987 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n1000, Z => n1303);
   U988 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n1541, Z => n1000);
   U989 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n1001, Z => n1304);
   U990 : MUXB2DL port map( A0 => b(2), A1 => n1545, SL => n1541, Z => n1001);
   U991 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n1002, Z => n1305);
   U992 : MUXB2DL port map( A0 => b(1), A1 => b(0), SL => n1541, Z => n1002);
   U993 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n1003, Z => n1306);
   U994 : NAN2M1D1 port map( A1 => n1541, A2 => b(0), Z => n1003);
   U995 : NOR2M1D1 port map( A1 => n1517, A2 => n14, Z => n1095);
   U996 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1004, Z => n1307);
   U997 : MUXB2DL port map( A0 => b(29), A1 => b(28), SL => n1542, Z => n1004);
   U998 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1005, Z => n1308);
   U999 : MUXB2DL port map( A0 => b(28), A1 => b(27), SL => n1542, Z => n1005);
   U1000 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1006, Z => n1309);
   U1001 : MUXB2DL port map( A0 => b(27), A1 => b(26), SL => n1542, Z => n1006)
                           ;
   U1002 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1007, Z => n1310);
   U1003 : MUXB2DL port map( A0 => b(26), A1 => b(25), SL => n1542, Z => n1007)
                           ;
   U1004 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1008, Z => n1311);
   U1005 : MUXB2DL port map( A0 => b(25), A1 => b(24), SL => n1542, Z => n1008)
                           ;
   U1006 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1009, Z => n1312);
   U1007 : MUXB2DL port map( A0 => b(24), A1 => b(23), SL => n1542, Z => n1009)
                           ;
   U1008 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1010, Z => n1313);
   U1009 : MUXB2DL port map( A0 => b(23), A1 => b(22), SL => n1542, Z => n1010)
                           ;
   U1010 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1011, Z => n1314);
   U1011 : MUXB2DL port map( A0 => b(22), A1 => b(21), SL => n1542, Z => n1011)
                           ;
   U1012 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1012, Z => n1315);
   U1013 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n1542, Z => n1012)
                           ;
   U1014 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1013, Z => n1316);
   U1015 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n1542, Z => n1013)
                           ;
   U1016 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1014, Z => n1317);
   U1017 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n1542, Z => n1014)
                           ;
   U1018 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1015, Z => n1318);
   U1019 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n1542, Z => n1015)
                           ;
   U1020 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1016, Z => n1319);
   U1021 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n1542, Z => n1016)
                           ;
   U1022 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1017, Z => n1320);
   U1023 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n1542, Z => n1017)
                           ;
   U1024 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1018, Z => n1321);
   U1025 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n1542, Z => n1018)
                           ;
   U1026 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1019, Z => n1322);
   U1027 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n1542, Z => n1019)
                           ;
   U1028 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1020, Z => n1323);
   U1029 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n1542, Z => n1020)
                           ;
   U1030 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1021, Z => n1324);
   U1031 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n1542, Z => n1021)
                           ;
   U1032 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1022, Z => n1325);
   U1033 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n1542, Z => n1022)
                           ;
   U1034 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1023, Z => n1326);
   U1035 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n1542, Z => n1023);
   U1036 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1024, Z => n1327);
   U1037 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n1542, Z => n1024);
   U1038 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1025, Z => n1328);
   U1039 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n1542, Z => n1025);
   U1040 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1026, Z => n1329);
   U1041 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n1542, Z => n1026);
   U1042 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1027, Z => n1330);
   U1043 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n1542, Z => n1027);
   U1044 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1028, Z => n1331);
   U1045 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n1542, Z => n1028);
   U1046 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1029, Z => n1332);
   U1047 : MUXB2DL port map( A0 => b(4), A1 => n1543, SL => n1542, Z => n1029);
   U1048 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1030, Z => n1333);
   U1049 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n1542, Z => n1030);
   U1050 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1031, Z => n1334);
   U1051 : MUXB2DL port map( A0 => b(2), A1 => n1545, SL => n1542, Z => n1031);
   U1052 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1032, Z => n1335);
   U1053 : MUXB2DL port map( A0 => b(1), A1 => b(0), SL => n1542, Z => n1032);
   U1054 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1033, Z => n1336);
   U1055 : NAN2M1D1 port map( A1 => n1542, A2 => b(0), Z => n1033);
   U1056 : NOR2M1D1 port map( A1 => n3, A2 => n6, Z => n1096);
   U1057 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1034, Z => n1337);
   U1058 : MUXB2DL port map( A0 => b(31), A1 => b(30), SL => n8, Z => n1034);
   U1059 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1035, Z => n1338);
   U1060 : MUXB2DL port map( A0 => b(30), A1 => b(29), SL => n8, Z => n1035);
   U1061 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1036, Z => n1339);
   U1062 : MUXB2DL port map( A0 => b(29), A1 => b(28), SL => n8, Z => n1036);
   U1063 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1037, Z => n1340);
   U1064 : MUXB2DL port map( A0 => b(28), A1 => b(27), SL => n8, Z => n1037);
   U1065 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1038, Z => n1341);
   U1066 : MUXB2DL port map( A0 => b(27), A1 => b(26), SL => n8, Z => n1038);
   U1067 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1039, Z => n1342);
   U1068 : MUXB2DL port map( A0 => b(26), A1 => b(25), SL => n8, Z => n1039);
   U1069 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1040, Z => n1343);
   U1070 : MUXB2DL port map( A0 => b(25), A1 => b(24), SL => n8, Z => n1040);
   U1071 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1041, Z => n1344);
   U1072 : MUXB2DL port map( A0 => b(24), A1 => b(23), SL => n8, Z => n1041);
   U1073 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1042, Z => n1345);
   U1074 : MUXB2DL port map( A0 => b(23), A1 => b(22), SL => n8, Z => n1042);
   U1075 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1043, Z => n1346);
   U1076 : MUXB2DL port map( A0 => b(22), A1 => b(21), SL => n8, Z => n1043);
   U1077 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1044, Z => n1347);
   U1078 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n8, Z => n1044);
   U1079 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1045, Z => n1348);
   U1080 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n8, Z => n1045);
   U1081 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1046, Z => n1349);
   U1082 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n8, Z => n1046);
   U1083 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1047, Z => n1350);
   U1084 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n8, Z => n1047);
   U1085 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1048, Z => n1351);
   U1086 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n8, Z => n1048);
   U1087 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1049, Z => n1352);
   U1088 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n8, Z => n1049);
   U1089 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1050, Z => n1353);
   U1090 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n8, Z => n1050);
   U1091 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1051, Z => n1354);
   U1092 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n8, Z => n1051);
   U1093 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1052, Z => n1355);
   U1094 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n8, Z => n1052);
   U1095 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1053, Z => n1356);
   U1096 : MUXB2DL port map( A0 => b(12), A1 => b(11), SL => n8, Z => n1053);
   U1097 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1054, Z => n1357);
   U1098 : MUXB2DL port map( A0 => b(11), A1 => b(10), SL => n8, Z => n1054);
   U1099 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1055, Z => n1358);
   U1100 : MUXB2DL port map( A0 => b(10), A1 => b(9), SL => n8, Z => n1055);
   U1101 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1056, Z => n1359);
   U1102 : MUXB2DL port map( A0 => b(9), A1 => b(8), SL => n8, Z => n1056);
   U1103 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1057, Z => n1360);
   U1104 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n8, Z => n1057);
   U1105 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1058, Z => n1361);
   U1106 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n8, Z => n1058);
   U1107 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1059, Z => n1362);
   U1108 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n8, Z => n1059);
   U1109 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1060, Z => n1363);
   U1110 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n8, Z => n1060);
   U1111 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1061, Z => n1364);
   U1112 : MUXB2DL port map( A0 => b(4), A1 => n1543, SL => n8, Z => n1061);
   U1113 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1062, Z => n1365);
   U1114 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n8, Z => n1062);
   U1115 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1063, Z => n1366);
   U1116 : MUXB2DL port map( A0 => b(2), A1 => n1545, SL => n8, Z => n1063);
   U1117 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1064, Z => n1367);
   U1118 : MUXB2DL port map( A0 => b(1), A1 => b(0), SL => n8, Z => n1064);
   U1119 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1065, Z => n1368);
   U1120 : NAN2M1D1 port map( A1 => n8, A2 => b(0), Z => n1065);
   U1121 : OAI21D1 port map( A1 => a(29), A2 => a(30), B => n1066, Z => n104);
   U1123 : EXNOR2D1 port map( A1 => a(29), A2 => a(30), Z => n106);
   U1125 : OAI21D1 port map( A1 => a(27), A2 => a(28), B => n1067, Z => n99);
   U1127 : EXNOR2D1 port map( A1 => a(27), A2 => a(28), Z => n103);
   U1129 : OAI21D1 port map( A1 => a(25), A2 => a(26), B => n1068, Z => n94);
   U1131 : EXNOR2D1 port map( A1 => a(25), A2 => a(26), Z => n98);
   U1135 : EXNOR2D1 port map( A1 => a(23), A2 => a(24), Z => n93);
   U1186 : ADHALFDL port map( A => n1278, B => n1093, CO => n780, S => n781);
   U1187 : OAI21D1 port map( A1 => a(1), A2 => a(2), B => n1080, Z => n1517);
   U1188 : OAI21D1 port map( A1 => a(3), A2 => a(4), B => n1079, Z => n1518);
   U1189 : OAI21D1 port map( A1 => a(7), A2 => a(8), B => n1077, Z => n1519);
   U1190 : AND2D1 port map( A1 => n1522, A2 => n305, Z => product(0));
   U1191 : AO21D1 port map( A1 => n215, A2 => n187, B => n188, Z => n1521);
   U1192 : OR2D1 port map( A1 => n1368, A2 => n1096, Z => n1522);
   U1193 : OA21M20D1 port map( A1 => n1523, A2 => n197, B => n194, Z => n190);
   U1194 : INVD1 port map( A => n215, Z => n214);
   U1195 : INVD1 port map( A => n233, Z => n232);
   U1196 : NAN2D1 port map( A1 => n313, A2 => n231, Z => n162);
   U1197 : INVD1 port map( A => n242, Z => n241);
   U1198 : INVD1 port map( A => n255, Z => n254);
   U1199 : INVD1 port map( A => n230, Z => n313);
   U1200 : INVD1 port map( A => n231, Z => n229);
   U1201 : INVD1 port map( A => n264, Z => n263);
   U1202 : NAN2D1 port map( A1 => n223, A2 => n1528, Z => n216);
   U1203 : INVD1 port map( A => n221, Z => n219);
   U1204 : NAN2D1 port map( A1 => n1530, A2 => n1529, Z => n243);
   U1205 : INVD1 port map( A => n248, Z => n246);
   U1206 : NAN2D1 port map( A1 => n1524, A2 => n1527, Z => n265);
   U1207 : INVD1 port map( A => n270, Z => n268);
   U1208 : NOR2D1 port map( A1 => n258, A2 => n261, Z => n256);
   U1209 : NOR2D1 port map( A1 => n236, A2 => n239, Z => n234);
   U1210 : NOR2D1 port map( A1 => n189, A2 => n201, Z => n187);
   U1211 : INVD1 port map( A => n209, Z => n211);
   U1212 : INVD1 port map( A => n206, Z => n204);
   U1213 : INVD1 port map( A => n275, Z => n273);
   U1214 : OR2D1 port map( A1 => n553, A2 => n574, Z => n1523);
   U1215 : NAN2D1 port map( A1 => n1523, A2 => n1526, Z => n189);
   U1216 : INVD1 port map( A => n199, Z => n197);
   U1217 : INVD1 port map( A => n253, Z => n251);
   U1218 : NAN2D1 port map( A1 => n667, A2 => n682, Z => n231);
   U1219 : NOR2D1 port map( A1 => n225, A2 => n230, Z => n223);
   U1220 : NAN2D1 port map( A1 => n1525, A2 => n310, Z => n201);
   U1221 : NOR2D1 port map( A1 => n683, A2 => n696, Z => n236);
   U1222 : NAN2D1 port map( A1 => n553, A2 => n574, Z => n194);
   U1223 : INVD1 port map( A => n208, Z => n310);
   U1224 : NOR2D1 port map( A1 => n667, A2 => n682, Z => n230);
   U1225 : NAN2D1 port map( A1 => n683, A2 => n696, Z => n237);
   U1226 : NAN2D1 port map( A1 => n1523, A2 => n194, Z => n156);
   U1227 : NAN2D1 port map( A1 => n1526, A2 => n199, Z => n157);
   U1228 : NAN2D1 port map( A1 => n1525, A2 => n206, Z => n158);
   U1229 : NAN2D1 port map( A1 => n310, A2 => n209, Z => n159);
   U1230 : NAN2D1 port map( A1 => n312, A2 => n226, Z => n161);
   U1231 : INVD1 port map( A => n225, Z => n312);
   U1232 : NAN2D1 port map( A1 => n1528, A2 => n221, Z => n160);
   U1233 : NAN2D1 port map( A1 => n314, A2 => n237, Z => n163);
   U1234 : INVD1 port map( A => n236, Z => n314);
   U1235 : NAN2D1 port map( A1 => n1530, A2 => n248, Z => n165);
   U1236 : NAN2D1 port map( A1 => n315, A2 => n240, Z => n164);
   U1237 : INVD1 port map( A => n239, Z => n315);
   U1238 : NAN2D1 port map( A1 => n1529, A2 => n253, Z => n166);
   U1239 : NAN2D1 port map( A1 => n318, A2 => n259, Z => n167);
   U1240 : INVD1 port map( A => n258, Z => n318);
   U1241 : NAN2D1 port map( A1 => n319, A2 => n262, Z => n168);
   U1242 : INVD1 port map( A => n261, Z => n319);
   U1243 : INVD1 port map( A => n277, Z => n276);
   U1244 : NAN2D1 port map( A1 => n1524, A2 => n270, Z => n169);
   U1245 : NAN2D1 port map( A1 => n1527, A2 => n275, Z => n170);
   U1246 : INVD1 port map( A => n286, Z => n285);
   U1247 : OR2D1 port map( A1 => n755, A2 => n762, Z => n1524);
   U1248 : NAN2D1 port map( A1 => n755, A2 => n762, Z => n270);
   U1249 : NOR2D1 port map( A1 => n280, A2 => n283, Z => n278);
   U1250 : OA21M20D1 port map( A1 => n1531, A2 => n294, B => n293, Z => n289);
   U1251 : NOR2D1 port map( A1 => n651, A2 => n666, Z => n225);
   U1252 : OA21M20D1 port map( A1 => n1532, A2 => n302, B => n301, Z => n297);
   U1253 : OR2D1 port map( A1 => n595, A2 => n614, Z => n1525);
   U1254 : NOR2D1 port map( A1 => n771, A2 => n776, Z => n280);
   U1255 : NOR2D1 port map( A1 => n745, A2 => n754, Z => n261);
   U1256 : NOR2D1 port map( A1 => n735, A2 => n744, Z => n258);
   U1257 : NAN2D1 port map( A1 => n763, A2 => n770, Z => n275);
   U1258 : OR2D1 port map( A1 => n575, A2 => n594, Z => n1526);
   U1259 : NAN2D1 port map( A1 => n575, A2 => n594, Z => n199);
   U1260 : NAN2D1 port map( A1 => n723, A2 => n734, Z => n253);
   U1261 : NAN2D1 port map( A1 => n651, A2 => n666, Z => n226);
   U1262 : OR2D1 port map( A1 => n763, A2 => n770, Z => n1527);
   U1263 : NAN2D1 port map( A1 => n595, A2 => n614, Z => n206);
   U1264 : OR2D1 port map( A1 => n633, A2 => n650, Z => n1528);
   U1265 : OR2D1 port map( A1 => n723, A2 => n734, Z => n1529);
   U1266 : NAN2D1 port map( A1 => n745, A2 => n754, Z => n262);
   U1267 : OR2D1 port map( A1 => n711, A2 => n722, Z => n1530);
   U1268 : NAN2D1 port map( A1 => n615, A2 => n632, Z => n209);
   U1269 : NAN2D1 port map( A1 => n771, A2 => n776, Z => n281);
   U1270 : NAN2D1 port map( A1 => n735, A2 => n744, Z => n259);
   U1271 : NOR2D1 port map( A1 => n615, A2 => n632, Z => n208);
   U1272 : NOR2D1 port map( A1 => n697, A2 => n710, Z => n239);
   U1273 : NAN2D1 port map( A1 => n711, A2 => n722, Z => n248);
   U1274 : NAN2D1 port map( A1 => n633, A2 => n650, Z => n221);
   U1275 : NAN2D1 port map( A1 => n697, A2 => n710, Z => n240);
   U1276 : NAN2D1 port map( A1 => n322, A2 => n281, Z => n171);
   U1277 : INVD1 port map( A => n280, Z => n322);
   U1278 : NAN2D1 port map( A1 => n323, A2 => n284, Z => n172);
   U1279 : INVD1 port map( A => n283, Z => n323);
   U1280 : NAN2D1 port map( A1 => n324, A2 => n288, Z => n173);
   U1281 : INVD1 port map( A => n287, Z => n324);
   U1282 : NAN2D1 port map( A1 => n1531, A2 => n293, Z => n174);
   U1283 : NAN2D1 port map( A1 => n326, A2 => n296, Z => n175);
   U1284 : INVD1 port map( A => n295, Z => n326);
   U1285 : NAN2D1 port map( A1 => n1532, A2 => n301, Z => n176);
   U1286 : OR2D1 port map( A1 => n787, A2 => n789, Z => n1531);
   U1287 : OR2D1 port map( A1 => n793, A2 => n1366, Z => n1532);
   U1288 : NOR2D1 port map( A1 => n777, A2 => n782, Z => n283);
   U1289 : NAN2D1 port map( A1 => n787, A2 => n789, Z => n293);
   U1290 : NAN2D1 port map( A1 => n793, A2 => n1366, Z => n301);
   U1291 : NAN2D1 port map( A1 => n777, A2 => n782, Z => n284);
   U1292 : NOR2D1 port map( A1 => n783, A2 => n786, Z => n287);
   U1293 : NOR2D1 port map( A1 => n791, A2 => n792, Z => n295);
   U1294 : NAN2D1 port map( A1 => n783, A2 => n786, Z => n288);
   U1295 : NAN2D1 port map( A1 => n791, A2 => n792, Z => n296);
   U1296 : NAN2D1 port map( A1 => n1368, A2 => n1096, Z => n305);
   U1297 : NOR2D1 port map( A1 => n303, A2 => n305, Z => n302);
   U1298 : INVD1 port map( A => n1533, Z => n1542);
   U1299 : EXOR2D1 port map( A1 => n178, A2 => n155, Z => product(31));
   U1300 : EXOR2D1 port map( A1 => n329, A2 => n344, Z => n155);
   U1301 : ADHALFDL port map( A => n1335, B => n1365, CO => n790, S => n791);
   U1302 : ADHALFDL port map( A => n1336, B => n1095, CO => n792, S => n793);
   U1303 : INVD1 port map( A => n1534, Z => n1539);
   U1304 : NOR2D1 port map( A1 => n1537, A2 => n30, Z => n1093);
   U1305 : INVD1 port map( A => n1535, Z => n1541);
   U1306 : INVD1 port map( A => n1536, Z => n1538);
   U1307 : ADHALFDL port map( A => n1331, B => n1361, CO => n774, S => n775);
   U1308 : ADHALFDL port map( A => n1252, B => n1092, CO => n768, S => n769);
   U1309 : ADHALFDL port map( A => n1333, B => n1363, CO => n784, S => n785);
   U1310 : ADHALFDL port map( A => n1306, B => n1094, CO => n788, S => n789);
   U1311 : INVD1 port map( A => n1537, Z => n1540);
   U1312 : ADHALFDL port map( A => n1206, B => n1090, CO => n732, S => n733);
   U1313 : ADHALFDL port map( A => n1168, B => n1088, CO => n680, S => n681);
   U1314 : ADHALFDL port map( A => n1152, B => n1087, CO => n648, S => n649);
   U1315 : ADHALFDL port map( A => n1228, B => n1091, CO => n752, S => n753);
   U1316 : ADHALFDL port map( A => n1186, B => n1089, CO => n708, S => n709);
   U1317 : ADHALFDL port map( A => n1138, B => n1086, CO => n612, S => n613);
   U1318 : INVD1 port map( A => n1367, Z => n303);
   U1319 : ADHALFDL port map( A => n1126, B => n1085, CO => n572, S => n573);
   U1320 : ADHALFDL port map( A => n1116, B => n1084, CO => n528, S => n529);
   U1321 : ADHALFDL port map( A => n1108, B => n1083, CO => n480, S => n481);
   U1322 : ADHALFDL port map( A => n1102, B => n1082, CO => n428, S => n429);
   U1323 : ADHALFDL port map( A => n1098, B => n1081, CO => n372, S => n373);
   U1324 : ADHALFDL port map( A => n1329, B => n1359, CO => n760, S => n761);
   U1325 : EXOR2D1 port map( A1 => a(1), A2 => a(2), Z => n1533);
   U1326 : ADHALFDL port map( A => n1323, B => n1353, CO => n694, S => n695);
   U1327 : EXOR2D1 port map( A1 => a(5), A2 => a(6), Z => n1534);
   U1328 : EXOR2D1 port map( A1 => a(3), A2 => a(4), Z => n1535);
   U1329 : EXOR2D1 port map( A1 => a(7), A2 => a(8), Z => n1536);
   U1330 : ADHALFDL port map( A => n1317, B => n1347, CO => n592, S => n593);
   U1331 : ADHALFDL port map( A => n1327, B => n1357, CO => n742, S => n743);
   U1332 : ADHALFDL port map( A => n1319, B => n1349, CO => n630, S => n631);
   U1333 : ADHALFDL port map( A => n1321, B => n1351, CO => n664, S => n665);
   U1334 : ADHALFDL port map( A => n1325, B => n1355, CO => n720, S => n721);
   U1335 : OA21D1 port map( A1 => a(5), A2 => a(6), B => n1078, Z => n1537);
   U1336 : INVD1 port map( A => a(3), Z => n1080);
   U1337 : EXNOR2D1 port map( A1 => a(11), A2 => a(12), Z => n56);
   U1338 : INVD1 port map( A => a(7), Z => n1078);
   U1339 : NAN2D1 port map( A1 => a(0), A2 => n6, Z => n3);
   U1340 : INVD1 port map( A => a(1), Z => n6);
   U1341 : INVD1 port map( A => a(9), Z => n1077);
   U1342 : EXNOR2D1 port map( A1 => a(13), A2 => a(14), Z => n63);
   U1343 : EXNOR2D1 port map( A1 => a(15), A2 => a(16), Z => n71);
   U1344 : INVD1 port map( A => a(5), Z => n1079);
   U1345 : EXNOR2D1 port map( A1 => a(9), A2 => a(10), Z => n48);
   U1346 : INVD1 port map( A => n1546, Z => n1545);
   U1347 : EXNOR2D1 port map( A1 => a(17), A2 => a(18), Z => n78);
   U1348 : AO21D1 port map( A1 => a(1), A2 => a(2), B => n1080, Z => n14);
   U1349 : INVD1 port map( A => n1544, Z => n1543);
   U1350 : AO21D1 port map( A1 => a(5), A2 => a(6), B => n1078, Z => n30);
   U1351 : INVD1 port map( A => a(0), Z => n8);
   U1352 : EXNOR2D1 port map( A1 => a(19), A2 => a(20), Z => n83);
   U1353 : AO21D1 port map( A1 => a(11), A2 => a(12), B => n1075, Z => n53);
   U1354 : INVD1 port map( A => a(13), Z => n1075);
   U1355 : ADHALFDL port map( A => n1315, B => n1345, CO => n550, S => n551);
   U1356 : AO21D1 port map( A1 => a(3), A2 => a(4), B => n1079, Z => n22);
   U1357 : AO21D1 port map( A1 => a(7), A2 => a(8), B => n1077, Z => n38);
   U1358 : OAI21D1 port map( A1 => a(11), A2 => a(12), B => n1075, Z => n50);
   U1359 : AO21D1 port map( A1 => a(13), A2 => a(14), B => n1074, Z => n61);
   U1360 : AO21D1 port map( A1 => a(15), A2 => a(16), B => n1073, Z => n69);
   U1361 : INVD1 port map( A => a(15), Z => n1074);
   U1362 : OAI21D1 port map( A1 => a(13), A2 => a(14), B => n1074, Z => n58);
   U1363 : INVD1 port map( A => a(17), Z => n1073);
   U1364 : OAI21D1 port map( A1 => a(15), A2 => a(16), B => n1073, Z => n66);
   U1365 : AO21D1 port map( A1 => a(9), A2 => a(10), B => n1076, Z => n45);
   U1366 : INVD1 port map( A => a(11), Z => n1076);
   U1367 : OAI21D1 port map( A1 => a(17), A2 => a(18), B => n1072, Z => n73);
   U1368 : INVD1 port map( A => a(19), Z => n1072);
   U1369 : OAI21D1 port map( A1 => a(9), A2 => a(10), B => n1076, Z => n42);
   U1370 : AO21D1 port map( A1 => a(17), A2 => a(18), B => n1072, Z => n76);
   U1371 : EXNOR2D1 port map( A1 => a(21), A2 => a(22), Z => n88);
   U1372 : OAI21D1 port map( A1 => a(19), A2 => a(20), B => n1071, Z => n79);
   U1373 : INVD1 port map( A => a(21), Z => n1071);
   U1374 : AO21D1 port map( A1 => a(19), A2 => a(20), B => n1071, Z => n81);
   U1375 : OAI21D1 port map( A1 => a(21), A2 => a(22), B => n1070, Z => n84);
   U1376 : INVD1 port map( A => a(23), Z => n1070);
   U1377 : AO21D1 port map( A1 => a(21), A2 => a(22), B => n1070, Z => n86);
   U1378 : ADHALFDL port map( A => n1313, B => n1343, CO => n504, S => n505);
   U1379 : OAI21D1 port map( A1 => a(23), A2 => a(24), B => n1069, Z => n89);
   U1380 : ADHALFDL port map( A => n1311, B => n1341, CO => n454, S => n455);
   U1381 : INVD1 port map( A => a(25), Z => n1069);
   U1382 : AO21D1 port map( A1 => a(23), A2 => a(24), B => n1069, Z => n91);
   U1383 : ADHALFDL port map( A => n1309, B => n1339, CO => n400, S => n401);
   U1384 : AO21D1 port map( A1 => a(25), A2 => a(26), B => n1068, Z => n96);
   U1385 : INVD1 port map( A => a(27), Z => n1068);
   U1386 : EXOR2D1 port map( A1 => n1307, A2 => n1337, Z => n343);
   U1387 : AO21D1 port map( A1 => a(27), A2 => a(28), B => n1067, Z => n101);
   U1388 : INVD1 port map( A => a(29), Z => n1067);
   U1389 : AO21D1 port map( A1 => a(29), A2 => a(30), B => n1066, Z => n105);
   U1390 : INVD1 port map( A => b(1), Z => n1546);
   U1391 : INVD1 port map( A => b(3), Z => n1544);
   U1392 : INVD1 port map( A => a(31), Z => n1066);

end hier_filter_none_5;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_gp_custom.all;

architecture hier_filter_none_5 of gp_custom_DW_mult_tc_5 is

   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AO21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OA21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component MUXB2DL
      port( A0, A1, SL : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component EXOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n6, n8, n14, n22, n30, n38, n42, n45, n48, n50, n53, n56, n58, 
      n61, n63, n66, n69, n71, n73, n76, n78, n79, n81, n83, n84, n86, n88, n89
      , n91, n93, n94, n96, n98, n99, n101, n103, n104, n105, n106, n155, n156,
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n178, n179, n180, n181, 
      n182, n183, n184, n185, n187, n188, n189, n190, n194, n195, n197, n199, 
      n200, n201, n202, n204, n206, n207, n208, n209, n211, n214, n215, n216, 
      n217, n219, n221, n222, n223, n224, n225, n226, n227, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n246, n248, n249, n251, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n268, n270, n271, n273, n275, 
      n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, 
      n288, n289, n293, n294, n295, n296, n297, n301, n302, n303, n305, n310, 
      n312, n313, n314, n315, n318, n319, n322, n323, n324, n326, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, 
      n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
      n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, 
      n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, 
      n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, 
      n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, 
      n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, 
      n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, 
      n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, 
      n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, 
      n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, 
      n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, 
      n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, 
      n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, 
      n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, 
      n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, 
      n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, 
      n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, 
      n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, 
      n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, 
      n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, 
      n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, 
      n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, 
      n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, 
      n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, 
      n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, 
      n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, 
      n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, 
      n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, 
      n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, 
      n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, 
      n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, 
      n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, 
      n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, 
      n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, 
      n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, 
      n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, 
      n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, 
      n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, 
      n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, 
      n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002
      , n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, 
      n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, 
      n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, 
      n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, 
      n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
      n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
      n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, 
      n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, 
      n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
      n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, 
      n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, 
      n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, 
      n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, 
      n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, 
      n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, 
      n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, 
      n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, 
      n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, 
      n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, 
      n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, 
      n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, 
      n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, 
      n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, 
      n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, 
      n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, 
      n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, 
      n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, 
      n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, 
      n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, 
      n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, 
      n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, 
      n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, 
      n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, 
      n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, 
      n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, 
      n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, 
      n1363, n1364, n1365, n1366, n1367, n1368, n1517, n1518, n1519, n1521, 
      n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, 
      n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, 
      n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549 : std_logic;

begin
   
   U125 : ADFULD1 port map( A => n345, B => n374, CI => n179, CO => n178, S => 
                           product(30));
   U126 : ADFULD1 port map( A => n375, B => n402, CI => n180, CO => n179, S => 
                           product(29));
   U127 : ADFULD1 port map( A => n403, B => n430, CI => n181, CO => n180, S => 
                           product(28));
   U128 : ADFULD1 port map( A => n431, B => n456, CI => n182, CO => n181, S => 
                           product(27));
   U129 : ADFULD1 port map( A => n457, B => n482, CI => n183, CO => n182, S => 
                           product(26));
   U130 : ADFULD1 port map( A => n483, B => n506, CI => n184, CO => n183, S => 
                           product(25));
   U131 : ADFULD1 port map( A => n507, B => n530, CI => n185, CO => n184, S => 
                           product(24));
   U132 : ADFULD1 port map( A => n531, B => n552, CI => n1521, CO => n185, S =>
                           product(23));
   U134 : EXOR2D1 port map( A1 => n195, A2 => n156, Z => product(22));
   U137 : OAI21D1 port map( A1 => n202, A2 => n189, B => n190, Z => n188);
   U146 : EXNOR2D1 port map( A1 => n200, A2 => n157, Z => product(21));
   U147 : AOI21D1 port map( A1 => n200, A2 => n1526, B => n197, Z => n195);
   U154 : EXNOR2D1 port map( A1 => n207, A2 => n158, Z => product(20));
   U155 : OAI21D1 port map( A1 => n214, A2 => n201, B => n202, Z => n200);
   U157 : AOI21D1 port map( A1 => n1525, A2 => n211, B => n204, Z => n202);
   U164 : EXOR2D1 port map( A1 => n214, A2 => n159, Z => product(19));
   U165 : OAI21D1 port map( A1 => n214, A2 => n208, B => n209, Z => n207);
   U174 : EXOR2D1 port map( A1 => n222, A2 => n160, Z => product(18));
   U176 : OAI21D1 port map( A1 => n233, A2 => n216, B => n217, Z => n215);
   U178 : AOI21D1 port map( A1 => n224, A2 => n1528, B => n219, Z => n217);
   U185 : EXOR2D1 port map( A1 => n227, A2 => n161, Z => product(17));
   U186 : AOI21D1 port map( A1 => n232, A2 => n223, B => n224, Z => n222);
   U188 : OAI21D1 port map( A1 => n225, A2 => n231, B => n226, Z => n224);
   U193 : EXNOR2D1 port map( A1 => n232, A2 => n162, Z => product(16));
   U194 : AOI21D1 port map( A1 => n232, A2 => n313, B => n229, Z => n227);
   U201 : EXNOR2D1 port map( A1 => n238, A2 => n163, Z => product(15));
   U203 : AOI21D1 port map( A1 => n242, A2 => n234, B => n235, Z => n233);
   U205 : OAI21D1 port map( A1 => n236, A2 => n240, B => n237, Z => n235);
   U210 : EXOR2D1 port map( A1 => n241, A2 => n164, Z => product(14));
   U211 : OAI21D1 port map( A1 => n241, A2 => n239, B => n240, Z => n238);
   U216 : EXOR2D1 port map( A1 => n249, A2 => n165, Z => product(13));
   U218 : OAI21D1 port map( A1 => n255, A2 => n243, B => n244, Z => n242);
   U220 : AOI21D1 port map( A1 => n1530, A2 => n251, B => n246, Z => n244);
   U227 : EXNOR2D1 port map( A1 => n254, A2 => n166, Z => product(12));
   U228 : AOI21D1 port map( A1 => n254, A2 => n1529, B => n251, Z => n249);
   U235 : EXNOR2D1 port map( A1 => n260, A2 => n167, Z => product(11));
   U237 : AOI21D1 port map( A1 => n256, A2 => n264, B => n257, Z => n255);
   U239 : OAI21D1 port map( A1 => n258, A2 => n262, B => n259, Z => n257);
   U244 : EXOR2D1 port map( A1 => n263, A2 => n168, Z => product(10));
   U245 : OAI21D1 port map( A1 => n263, A2 => n261, B => n262, Z => n260);
   U250 : EXOR2D1 port map( A1 => n271, A2 => n169, Z => product(9));
   U252 : OAI21D1 port map( A1 => n265, A2 => n277, B => n266, Z => n264);
   U254 : AOI21D1 port map( A1 => n1524, A2 => n273, B => n268, Z => n266);
   U261 : EXNOR2D1 port map( A1 => n276, A2 => n170, Z => product(8));
   U262 : AOI21D1 port map( A1 => n276, A2 => n1527, B => n273, Z => n271);
   U269 : EXNOR2D1 port map( A1 => n282, A2 => n171, Z => product(7));
   U271 : AOI21D1 port map( A1 => n278, A2 => n286, B => n279, Z => n277);
   U273 : OAI21D1 port map( A1 => n280, A2 => n284, B => n281, Z => n279);
   U278 : EXOR2D1 port map( A1 => n172, A2 => n285, Z => product(6));
   U279 : OAI21D1 port map( A1 => n285, A2 => n283, B => n284, Z => n282);
   U284 : EXOR2D1 port map( A1 => n173, A2 => n289, Z => product(5));
   U286 : OAI21D1 port map( A1 => n289, A2 => n287, B => n288, Z => n286);
   U291 : EXNOR2D1 port map( A1 => n174, A2 => n294, Z => product(4));
   U299 : EXOR2D1 port map( A1 => n297, A2 => n175, Z => product(3));
   U300 : OAI21D1 port map( A1 => n297, A2 => n295, B => n296, Z => n294);
   U305 : EXNOR2D1 port map( A1 => n176, A2 => n302, Z => product(2));
   U313 : EXOR2D1 port map( A1 => n303, A2 => n305, Z => product(1));
   U321 : EXOR3D1 port map( A1 => n346, A2 => n331, A3 => n330, Z => n329);
   U322 : EXOR3D1 port map( A1 => n332, A2 => n350, A3 => n348, Z => n330);
   U323 : EXOR3D1 port map( A1 => n352, A2 => n334, A3 => n333, Z => n331);
   U324 : EXOR3D1 port map( A1 => n354, A2 => n356, A3 => n335, Z => n332);
   U325 : EXOR3D1 port map( A1 => n337, A2 => n358, A3 => n336, Z => n333);
   U326 : EXOR3D1 port map( A1 => n339, A2 => n340, A3 => n360, Z => n334);
   U327 : EXOR3D1 port map( A1 => n342, A2 => n338, A3 => n341, Z => n335);
   U328 : EXOR3D1 port map( A1 => n366, A2 => n343, A3 => n362, Z => n336);
   U329 : EXOR3D1 port map( A1 => n368, A2 => n370, A3 => n364, Z => n337);
   U330 : EXOR3D1 port map( A1 => n1187, A2 => n1169, A3 => n372, Z => n338);
   U331 : EXOR3D1 port map( A1 => n1139, A2 => n1229, A3 => n1153, Z => n339);
   U332 : EXOR3D1 port map( A1 => n1103, A2 => n1117, A3 => n1109, Z => n340);
   U333 : EXOR3D1 port map( A1 => n1253, A2 => n1127, A3 => n1099, Z => n341);
   U334 : EXOR3D1 port map( A1 => n1097, A2 => n1279, A3 => n1207, Z => n342);
   U336 : ADFULD1 port map( A => n376, B => n349, CI => n347, CO => n344, S => 
                           n345);
   U337 : ADFULD1 port map( A => n351, B => n353, CI => n378, CO => n346, S => 
                           n347);
   U338 : ADFULD1 port map( A => n382, B => n355, CI => n380, CO => n348, S => 
                           n349);
   U339 : ADFULD1 port map( A => n359, B => n384, CI => n357, CO => n350, S => 
                           n351);
   U340 : ADFULD1 port map( A => n361, B => n388, CI => n386, CO => n352, S => 
                           n353);
   U341 : ADFULD1 port map( A => n365, B => n363, CI => n390, CO => n354, S => 
                           n355);
   U342 : ADFULD1 port map( A => n369, B => n371, CI => n367, CO => n356, S => 
                           n357);
   U343 : ADFULD1 port map( A => n398, B => n394, CI => n396, CO => n358, S => 
                           n359);
   U344 : ADFULD1 port map( A => n373, B => n400, CI => n392, CO => n360, S => 
                           n361);
   U345 : ADFULD1 port map( A => n1170, B => n1118, CI => n1140, CO => n362, S 
                           => n363);
   U346 : ADFULD1 port map( A => n1104, B => n1188, CI => n1110, CO => n364, S 
                           => n365);
   U347 : ADFULD1 port map( A => n1254, B => n1128, CI => n1230, CO => n366, S 
                           => n367);
   U348 : ADFULD1 port map( A => n1280, B => n1154, CI => n1208, CO => n368, S 
                           => n369);
   U349 : ADFULD1 port map( A => n1100, B => n1338, CI => n1308, CO => n370, S 
                           => n371);
   U351 : ADFULD1 port map( A => n404, B => n379, CI => n377, CO => n374, S => 
                           n375);
   U352 : ADFULD1 port map( A => n381, B => n408, CI => n406, CO => n376, S => 
                           n377);
   U353 : ADFULD1 port map( A => n410, B => n385, CI => n383, CO => n378, S => 
                           n379);
   U354 : ADFULD1 port map( A => n412, B => n389, CI => n387, CO => n380, S => 
                           n381);
   U355 : ADFULD1 port map( A => n391, B => n416, CI => n414, CO => n382, S => 
                           n383);
   U356 : ADFULD1 port map( A => n395, B => n397, CI => n399, CO => n384, S => 
                           n385);
   U357 : ADFULD1 port map( A => n418, B => n422, CI => n393, CO => n386, S => 
                           n387);
   U358 : ADFULD1 port map( A => n424, B => n426, CI => n420, CO => n388, S => 
                           n389);
   U359 : ADFULD1 port map( A => n428, B => n1171, CI => n401, CO => n390, S =>
                           n391);
   U360 : ADFULD1 port map( A => n1129, B => n1189, CI => n1141, CO => n392, S 
                           => n393);
   U361 : ADFULD1 port map( A => n1231, B => n1111, CI => n1105, CO => n394, S 
                           => n395);
   U362 : ADFULD1 port map( A => n1255, B => n1119, CI => n1101, CO => n396, S 
                           => n397);
   U363 : ADFULD1 port map( A => n1281, B => n1155, CI => n1209, CO => n398, S 
                           => n399);
   U365 : ADFULD1 port map( A => n432, B => n407, CI => n405, CO => n402, S => 
                           n403);
   U366 : ADFULD1 port map( A => n409, B => n436, CI => n434, CO => n404, S => 
                           n405);
   U367 : ADFULD1 port map( A => n438, B => n413, CI => n411, CO => n406, S => 
                           n407);
   U368 : ADFULD1 port map( A => n440, B => n417, CI => n415, CO => n408, S => 
                           n409);
   U369 : ADFULD1 port map( A => n444, B => n419, CI => n442, CO => n410, S => 
                           n411);
   U370 : ADFULD1 port map( A => n421, B => n423, CI => n425, CO => n412, S => 
                           n413);
   U371 : ADFULD1 port map( A => n448, B => n446, CI => n427, CO => n414, S => 
                           n415);
   U372 : ADFULD1 port map( A => n452, B => n429, CI => n450, CO => n416, S => 
                           n417);
   U373 : ADFULD1 port map( A => n1232, B => n1190, CI => n454, CO => n418, S 
                           => n419);
   U374 : ADFULD1 port map( A => n1142, B => n1256, CI => n1172, CO => n420, S 
                           => n421);
   U375 : ADFULD1 port map( A => n1112, B => n1130, CI => n1120, CO => n422, S 
                           => n423);
   U376 : ADFULD1 port map( A => n1282, B => n1156, CI => n1210, CO => n424, S 
                           => n425);
   U377 : ADFULD1 port map( A => n1106, B => n1340, CI => n1310, CO => n426, S 
                           => n427);
   U379 : ADFULD1 port map( A => n458, B => n435, CI => n433, CO => n430, S => 
                           n431);
   U380 : ADFULD1 port map( A => n437, B => n439, CI => n460, CO => n432, S => 
                           n433);
   U381 : ADFULD1 port map( A => n441, B => n464, CI => n462, CO => n434, S => 
                           n435);
   U382 : ADFULD1 port map( A => n466, B => n445, CI => n443, CO => n436, S => 
                           n437);
   U383 : ADFULD1 port map( A => n449, B => n451, CI => n468, CO => n438, S => 
                           n439);
   U384 : ADFULD1 port map( A => n453, B => n447, CI => n470, CO => n440, S => 
                           n441);
   U385 : ADFULD1 port map( A => n474, B => n472, CI => n476, CO => n442, S => 
                           n443);
   U386 : ADFULD1 port map( A => n455, B => n480, CI => n478, CO => n444, S => 
                           n445);
   U387 : ADFULD1 port map( A => n1131, B => n1191, CI => n1173, CO => n446, S 
                           => n447);
   U388 : ADFULD1 port map( A => n1113, B => n1233, CI => n1121, CO => n448, S 
                           => n449);
   U389 : ADFULD1 port map( A => n1283, B => n1143, CI => n1257, CO => n450, S 
                           => n451);
   U390 : ADFULD1 port map( A => n1107, B => n1157, CI => n1211, CO => n452, S 
                           => n453);
   U392 : ADFULD1 port map( A => n484, B => n461, CI => n459, CO => n456, S => 
                           n457);
   U393 : ADFULD1 port map( A => n486, B => n488, CI => n463, CO => n458, S => 
                           n459);
   U394 : ADFULD1 port map( A => n467, B => n469, CI => n465, CO => n460, S => 
                           n461);
   U395 : ADFULD1 port map( A => n492, B => n494, CI => n490, CO => n462, S => 
                           n463);
   U396 : ADFULD1 port map( A => n475, B => n477, CI => n471, CO => n464, S => 
                           n465);
   U397 : ADFULD1 port map( A => n479, B => n500, CI => n473, CO => n466, S => 
                           n467);
   U398 : ADFULD1 port map( A => n498, B => n502, CI => n496, CO => n468, S => 
                           n469);
   U399 : ADFULD1 port map( A => n504, B => n1192, CI => n481, CO => n470, S =>
                           n471);
   U400 : ADFULD1 port map( A => n1144, B => n1234, CI => n1158, CO => n472, S 
                           => n473);
   U401 : ADFULD1 port map( A => n1258, B => n1132, CI => n1122, CO => n474, S 
                           => n475);
   U402 : ADFULD1 port map( A => n1284, B => n1174, CI => n1212, CO => n476, S 
                           => n477);
   U403 : ADFULD1 port map( A => n1114, B => n1342, CI => n1312, CO => n478, S 
                           => n479);
   U405 : ADFULD1 port map( A => n508, B => n487, CI => n485, CO => n482, S => 
                           n483);
   U406 : ADFULD1 port map( A => n510, B => n512, CI => n489, CO => n484, S => 
                           n485);
   U407 : ADFULD1 port map( A => n493, B => n514, CI => n491, CO => n486, S => 
                           n487);
   U408 : ADFULD1 port map( A => n516, B => n518, CI => n495, CO => n488, S => 
                           n489);
   U409 : ADFULD1 port map( A => n501, B => n503, CI => n497, CO => n490, S => 
                           n491);
   U410 : ADFULD1 port map( A => n522, B => n524, CI => n499, CO => n492, S => 
                           n493);
   U411 : ADFULD1 port map( A => n526, B => n505, CI => n520, CO => n494, S => 
                           n495);
   U412 : ADFULD1 port map( A => n1235, B => n1259, CI => n528, CO => n496, S 
                           => n497);
   U413 : ADFULD1 port map( A => n1159, B => n1285, CI => n1193, CO => n498, S 
                           => n499);
   U414 : ADFULD1 port map( A => n1123, B => n1145, CI => n1133, CO => n500, S 
                           => n501);
   U415 : ADFULD1 port map( A => n1115, B => n1175, CI => n1213, CO => n502, S 
                           => n503);
   U417 : ADFULD1 port map( A => n532, B => n511, CI => n509, CO => n506, S => 
                           n507);
   U418 : ADFULD1 port map( A => n513, B => n536, CI => n534, CO => n508, S => 
                           n509);
   U419 : ADFULD1 port map( A => n517, B => n538, CI => n515, CO => n510, S => 
                           n511);
   U420 : ADFULD1 port map( A => n540, B => n542, CI => n519, CO => n512, S => 
                           n513);
   U421 : ADFULD1 port map( A => n525, B => n521, CI => n523, CO => n514, S => 
                           n515);
   U422 : ADFULD1 port map( A => n544, B => n546, CI => n527, CO => n516, S => 
                           n517);
   U423 : ADFULD1 port map( A => n529, B => n550, CI => n548, CO => n518, S => 
                           n519);
   U424 : ADFULD1 port map( A => n1194, B => n1260, CI => n1236, CO => n520, S 
                           => n521);
   U425 : ADFULD1 port map( A => n1134, B => n1286, CI => n1160, CO => n522, S 
                           => n523);
   U426 : ADFULD1 port map( A => n1124, B => n1176, CI => n1214, CO => n524, S 
                           => n525);
   U427 : ADFULD1 port map( A => n1146, B => n1344, CI => n1314, CO => n526, S 
                           => n527);
   U429 : ADFULD1 port map( A => n554, B => n535, CI => n533, CO => n530, S => 
                           n531);
   U430 : ADFULD1 port map( A => n556, B => n539, CI => n537, CO => n532, S => 
                           n533);
   U431 : ADFULD1 port map( A => n541, B => n560, CI => n558, CO => n534, S => 
                           n535);
   U432 : ADFULD1 port map( A => n562, B => n545, CI => n543, CO => n536, S => 
                           n537);
   U433 : ADFULD1 port map( A => n549, B => n564, CI => n547, CO => n538, S => 
                           n539);
   U434 : ADFULD1 port map( A => n566, B => n570, CI => n568, CO => n540, S => 
                           n541);
   U435 : ADFULD1 port map( A => n572, B => n1195, CI => n551, CO => n542, S =>
                           n543);
   U436 : ADFULD1 port map( A => n1135, B => n1237, CI => n1147, CO => n544, S 
                           => n545);
   U437 : ADFULD1 port map( A => n1287, B => n1161, CI => n1261, CO => n546, S 
                           => n547);
   U438 : ADFULD1 port map( A => n1125, B => n1177, CI => n1215, CO => n548, S 
                           => n549);
   U440 : ADFULD1 port map( A => n576, B => n557, CI => n555, CO => n552, S => 
                           n553);
   U441 : ADFULD1 port map( A => n559, B => n561, CI => n578, CO => n554, S => 
                           n555);
   U442 : ADFULD1 port map( A => n563, B => n582, CI => n580, CO => n556, S => 
                           n557);
   U443 : ADFULD1 port map( A => n565, B => n569, CI => n584, CO => n558, S => 
                           n559);
   U444 : ADFULD1 port map( A => n571, B => n586, CI => n567, CO => n560, S => 
                           n561);
   U445 : ADFULD1 port map( A => n590, B => n573, CI => n588, CO => n562, S => 
                           n563);
   U446 : ADFULD1 port map( A => n1196, B => n1238, CI => n592, CO => n564, S 
                           => n565);
   U447 : ADFULD1 port map( A => n1148, B => n1262, CI => n1162, CO => n566, S 
                           => n567);
   U448 : ADFULD1 port map( A => n1288, B => n1178, CI => n1216, CO => n568, S 
                           => n569);
   U449 : ADFULD1 port map( A => n1136, B => n1346, CI => n1316, CO => n570, S 
                           => n571);
   U451 : ADFULD1 port map( A => n596, B => n579, CI => n577, CO => n574, S => 
                           n575);
   U452 : ADFULD1 port map( A => n581, B => n583, CI => n598, CO => n576, S => 
                           n577);
   U453 : ADFULD1 port map( A => n585, B => n602, CI => n600, CO => n578, S => 
                           n579);
   U454 : ADFULD1 port map( A => n591, B => n589, CI => n604, CO => n580, S => 
                           n581);
   U455 : ADFULD1 port map( A => n606, B => n608, CI => n587, CO => n582, S => 
                           n583);
   U456 : ADFULD1 port map( A => n593, B => n612, CI => n610, CO => n584, S => 
                           n585);
   U457 : ADFULD1 port map( A => n1163, B => n1239, CI => n1197, CO => n586, S 
                           => n587);
   U458 : ADFULD1 port map( A => n1263, B => n1149, CI => n1137, CO => n588, S 
                           => n589);
   U459 : ADFULD1 port map( A => n1289, B => n1179, CI => n1217, CO => n590, S 
                           => n591);
   U461 : ADFULD1 port map( A => n616, B => n599, CI => n597, CO => n594, S => 
                           n595);
   U462 : ADFULD1 port map( A => n601, B => n603, CI => n618, CO => n596, S => 
                           n597);
   U463 : ADFULD1 port map( A => n622, B => n605, CI => n620, CO => n598, S => 
                           n599);
   U464 : ADFULD1 port map( A => n609, B => n611, CI => n607, CO => n600, S => 
                           n601);
   U465 : ADFULD1 port map( A => n626, B => n628, CI => n624, CO => n602, S => 
                           n603);
   U466 : ADFULD1 port map( A => n630, B => n1240, CI => n613, CO => n604, S =>
                           n605);
   U467 : ADFULD1 port map( A => n1150, B => n1264, CI => n1180, CO => n606, S 
                           => n607);
   U468 : ADFULD1 port map( A => n1290, B => n1198, CI => n1218, CO => n608, S 
                           => n609);
   U469 : ADFULD1 port map( A => n1164, B => n1348, CI => n1318, CO => n610, S 
                           => n611);
   U471 : ADFULD1 port map( A => n634, B => n619, CI => n617, CO => n614, S => 
                           n615);
   U472 : ADFULD1 port map( A => n621, B => n623, CI => n636, CO => n616, S => 
                           n617);
   U473 : ADFULD1 port map( A => n640, B => n625, CI => n638, CO => n618, S => 
                           n619);
   U474 : ADFULD1 port map( A => n627, B => n644, CI => n629, CO => n620, S => 
                           n621);
   U475 : ADFULD1 port map( A => n646, B => n631, CI => n642, CO => n622, S => 
                           n623);
   U476 : ADFULD1 port map( A => n1241, B => n1265, CI => n648, CO => n624, S 
                           => n625);
   U477 : ADFULD1 port map( A => n1291, B => n1181, CI => n1165, CO => n626, S 
                           => n627);
   U478 : ADFULD1 port map( A => n1151, B => n1199, CI => n1219, CO => n628, S 
                           => n629);
   U480 : ADFULD1 port map( A => n652, B => n637, CI => n635, CO => n632, S => 
                           n633);
   U481 : ADFULD1 port map( A => n639, B => n641, CI => n654, CO => n634, S => 
                           n635);
   U482 : ADFULD1 port map( A => n658, B => n645, CI => n656, CO => n636, S => 
                           n637);
   U483 : ADFULD1 port map( A => n647, B => n660, CI => n643, CO => n638, S => 
                           n639);
   U484 : ADFULD1 port map( A => n649, B => n664, CI => n662, CO => n640, S => 
                           n641);
   U485 : ADFULD1 port map( A => n1182, B => n1292, CI => n1242, CO => n642, S 
                           => n643);
   U486 : ADFULD1 port map( A => n1166, B => n1266, CI => n1220, CO => n644, S 
                           => n645);
   U487 : ADFULD1 port map( A => n1200, B => n1350, CI => n1320, CO => n646, S 
                           => n647);
   U489 : ADFULD1 port map( A => n668, B => n655, CI => n653, CO => n650, S => 
                           n651);
   U490 : ADFULD1 port map( A => n670, B => n659, CI => n657, CO => n652, S => 
                           n653);
   U491 : ADFULD1 port map( A => n663, B => n661, CI => n672, CO => n654, S => 
                           n655);
   U492 : ADFULD1 port map( A => n676, B => n678, CI => n674, CO => n656, S => 
                           n657);
   U493 : ADFULD1 port map( A => n680, B => n1267, CI => n665, CO => n658, S =>
                           n659);
   U494 : ADFULD1 port map( A => n1183, B => n1167, CI => n1243, CO => n660, S 
                           => n661);
   U495 : ADFULD1 port map( A => n1293, B => n1201, CI => n1221, CO => n662, S 
                           => n663);
   U497 : ADFULD1 port map( A => n684, B => n671, CI => n669, CO => n666, S => 
                           n667);
   U498 : ADFULD1 port map( A => n686, B => n688, CI => n673, CO => n668, S => 
                           n669);
   U499 : ADFULD1 port map( A => n677, B => n679, CI => n675, CO => n670, S => 
                           n671);
   U500 : ADFULD1 port map( A => n692, B => n681, CI => n690, CO => n672, S => 
                           n673);
   U501 : ADFULD1 port map( A => n1244, B => n1294, CI => n694, CO => n674, S 
                           => n675);
   U502 : ADFULD1 port map( A => n1184, B => n1268, CI => n1222, CO => n676, S 
                           => n677);
   U503 : ADFULD1 port map( A => n1202, B => n1352, CI => n1322, CO => n678, S 
                           => n679);
   U505 : ADFULD1 port map( A => n698, B => n687, CI => n685, CO => n682, S => 
                           n683);
   U506 : ADFULD1 port map( A => n700, B => n702, CI => n689, CO => n684, S => 
                           n685);
   U507 : ADFULD1 port map( A => n691, B => n704, CI => n693, CO => n686, S => 
                           n687);
   U508 : ADFULD1 port map( A => n695, B => n708, CI => n706, CO => n688, S => 
                           n689);
   U509 : ADFULD1 port map( A => n1185, B => n1245, CI => n1203, CO => n690, S 
                           => n691);
   U510 : ADFULD1 port map( A => n1295, B => n1269, CI => n1223, CO => n692, S 
                           => n693);
   U512 : ADFULD1 port map( A => n712, B => n701, CI => n699, CO => n696, S => 
                           n697);
   U513 : ADFULD1 port map( A => n703, B => n705, CI => n714, CO => n698, S => 
                           n699);
   U514 : ADFULD1 port map( A => n716, B => n718, CI => n707, CO => n700, S => 
                           n701);
   U515 : ADFULD1 port map( A => n720, B => n1270, CI => n709, CO => n702, S =>
                           n703);
   U516 : ADFULD1 port map( A => n1246, B => n1296, CI => n1224, CO => n704, S 
                           => n705);
   U517 : ADFULD1 port map( A => n1204, B => n1354, CI => n1324, CO => n706, S 
                           => n707);
   U519 : ADFULD1 port map( A => n724, B => n715, CI => n713, CO => n710, S => 
                           n711);
   U520 : ADFULD1 port map( A => n717, B => n719, CI => n726, CO => n712, S => 
                           n713);
   U521 : ADFULD1 port map( A => n730, B => n721, CI => n728, CO => n714, S => 
                           n715);
   U522 : ADFULD1 port map( A => n1205, B => n1247, CI => n732, CO => n716, S 
                           => n717);
   U523 : ADFULD1 port map( A => n1271, B => n1297, CI => n1225, CO => n718, S 
                           => n719);
   U525 : ADFULD1 port map( A => n736, B => n727, CI => n725, CO => n722, S => 
                           n723);
   U526 : ADFULD1 port map( A => n729, B => n731, CI => n738, CO => n724, S => 
                           n725);
   U527 : ADFULD1 port map( A => n733, B => n742, CI => n740, CO => n726, S => 
                           n727);
   U528 : ADFULD1 port map( A => n1272, B => n1298, CI => n1226, CO => n728, S 
                           => n729);
   U529 : ADFULD1 port map( A => n1248, B => n1356, CI => n1326, CO => n730, S 
                           => n731);
   U531 : ADFULD1 port map( A => n746, B => n739, CI => n737, CO => n734, S => 
                           n735);
   U532 : ADFULD1 port map( A => n748, B => n750, CI => n741, CO => n736, S => 
                           n737);
   U533 : ADFULD1 port map( A => n752, B => n1299, CI => n743, CO => n738, S =>
                           n739);
   U534 : ADFULD1 port map( A => n1273, B => n1249, CI => n1227, CO => n740, S 
                           => n741);
   U536 : ADFULD1 port map( A => n756, B => n749, CI => n747, CO => n744, S => 
                           n745);
   U537 : ADFULD1 port map( A => n758, B => n753, CI => n751, CO => n746, S => 
                           n747);
   U538 : ADFULD1 port map( A => n1274, B => n1300, CI => n760, CO => n748, S 
                           => n749);
   U539 : ADFULD1 port map( A => n1250, B => n1358, CI => n1328, CO => n750, S 
                           => n751);
   U541 : ADFULD1 port map( A => n764, B => n759, CI => n757, CO => n754, S => 
                           n755);
   U542 : ADFULD1 port map( A => n761, B => n768, CI => n766, CO => n756, S => 
                           n757);
   U543 : ADFULD1 port map( A => n1275, B => n1251, CI => n1301, CO => n758, S 
                           => n759);
   U545 : ADFULD1 port map( A => n767, B => n772, CI => n765, CO => n762, S => 
                           n763);
   U546 : ADFULD1 port map( A => n774, B => n1302, CI => n769, CO => n764, S =>
                           n765);
   U547 : ADFULD1 port map( A => n1276, B => n1360, CI => n1330, CO => n766, S 
                           => n767);
   U549 : ADFULD1 port map( A => n778, B => n775, CI => n773, CO => n770, S => 
                           n771);
   U550 : ADFULD1 port map( A => n1277, B => n1303, CI => n780, CO => n772, S 
                           => n773);
   U552 : ADFULD1 port map( A => n781, B => n784, CI => n779, CO => n776, S => 
                           n777);
   U553 : ADFULD1 port map( A => n1304, B => n1362, CI => n1332, CO => n778, S 
                           => n779);
   U555 : ADFULD1 port map( A => n788, B => n1305, CI => n785, CO => n782, S =>
                           n783);
   U557 : ADFULD1 port map( A => n1334, B => n1364, CI => n790, CO => n786, S 
                           => n787);
   U561 : NOR2M1D1 port map( A1 => n104, A2 => n105, Z => n1081);
   U562 : MUXB2DL port map( A0 => n104, A1 => n105, SL => n794, Z => n1097);
   U563 : MUXB2DL port map( A0 => b(1), A1 => n1548, SL => n106, Z => n794);
   U564 : MUXB2DL port map( A0 => n104, A1 => n105, SL => n795, Z => n1098);
   U565 : NAN2M1D1 port map( A1 => n106, A2 => b(0), Z => n795);
   U566 : NOR2M1D1 port map( A1 => n99, A2 => n101, Z => n1082);
   U567 : MUXB2DL port map( A0 => n99, A1 => n101, SL => n796, Z => n1099);
   U568 : MUXB2DL port map( A0 => b(3), A1 => n1546, SL => n103, Z => n796);
   U569 : MUXB2DL port map( A0 => n99, A1 => n101, SL => n797, Z => n1100);
   U570 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n103, Z => n797);
   U571 : MUXB2DL port map( A0 => n99, A1 => n101, SL => n798, Z => n1101);
   U572 : MUXB2DL port map( A0 => b(1), A1 => n1548, SL => n103, Z => n798);
   U573 : MUXB2DL port map( A0 => n99, A1 => n101, SL => n799, Z => n1102);
   U574 : NAN2M1D1 port map( A1 => n103, A2 => b(0), Z => n799);
   U575 : NOR2M1D1 port map( A1 => n94, A2 => n96, Z => n1083);
   U576 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n800, Z => n1103);
   U577 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n98, Z => n800);
   U578 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n801, Z => n1104);
   U579 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n98, Z => n801);
   U580 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n802, Z => n1105);
   U581 : MUXB2DL port map( A0 => b(3), A1 => n1546, SL => n98, Z => n802);
   U582 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n803, Z => n1106);
   U583 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n98, Z => n803);
   U584 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n804, Z => n1107);
   U585 : MUXB2DL port map( A0 => b(1), A1 => n1548, SL => n98, Z => n804);
   U586 : MUXB2DL port map( A0 => n94, A1 => n96, SL => n805, Z => n1108);
   U587 : NAN2M1D1 port map( A1 => n98, A2 => b(0), Z => n805);
   U588 : NOR2M1D1 port map( A1 => n89, A2 => n91, Z => n1084);
   U589 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n806, Z => n1109);
   U590 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n93, Z => n806);
   U591 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n807, Z => n1110);
   U592 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n93, Z => n807);
   U593 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n808, Z => n1111);
   U594 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n93, Z => n808);
   U595 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n809, Z => n1112);
   U596 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n93, Z => n809);
   U597 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n810, Z => n1113);
   U598 : MUXB2DL port map( A0 => b(3), A1 => n1546, SL => n93, Z => n810);
   U599 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n811, Z => n1114);
   U600 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n93, Z => n811);
   U601 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n812, Z => n1115);
   U602 : MUXB2DL port map( A0 => b(1), A1 => n1548, SL => n93, Z => n812);
   U603 : MUXB2DL port map( A0 => n89, A1 => n91, SL => n813, Z => n1116);
   U604 : NAN2M1D1 port map( A1 => n93, A2 => n1548, Z => n813);
   U605 : NOR2M1D1 port map( A1 => n84, A2 => n86, Z => n1085);
   U606 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n814, Z => n1117);
   U607 : MUXB2DL port map( A0 => n1538, A1 => b(8), SL => n88, Z => n814);
   U608 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n815, Z => n1118);
   U609 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n88, Z => n815);
   U610 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n816, Z => n1119);
   U611 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n88, Z => n816);
   U612 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n817, Z => n1120);
   U613 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n88, Z => n817);
   U614 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n818, Z => n1121);
   U615 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n88, Z => n818);
   U616 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n819, Z => n1122);
   U617 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n88, Z => n819);
   U618 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n820, Z => n1123);
   U619 : MUXB2DL port map( A0 => b(3), A1 => n1546, SL => n88, Z => n820);
   U620 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n821, Z => n1124);
   U621 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n88, Z => n821);
   U622 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n822, Z => n1125);
   U623 : MUXB2DL port map( A0 => b(1), A1 => n1548, SL => n88, Z => n822);
   U624 : MUXB2DL port map( A0 => n84, A1 => n86, SL => n823, Z => n1126);
   U625 : NAN2M1D1 port map( A1 => n88, A2 => n1548, Z => n823);
   U626 : NOR2M1D1 port map( A1 => n79, A2 => n81, Z => n1086);
   U627 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n824, Z => n1127);
   U628 : MUXB2DL port map( A0 => n1540, A1 => n1539, SL => n83, Z => n824);
   U629 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n825, Z => n1128);
   U630 : MUXB2DL port map( A0 => n1539, A1 => n1538, SL => n83, Z => n825);
   U631 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n826, Z => n1129);
   U632 : MUXB2DL port map( A0 => n1538, A1 => b(8), SL => n83, Z => n826);
   U633 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n827, Z => n1130);
   U634 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n83, Z => n827);
   U635 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n828, Z => n1131);
   U636 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n83, Z => n828);
   U637 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n829, Z => n1132);
   U638 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n83, Z => n829);
   U639 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n830, Z => n1133);
   U640 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n83, Z => n830);
   U641 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n831, Z => n1134);
   U642 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n83, Z => n831);
   U643 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n832, Z => n1135);
   U644 : MUXB2DL port map( A0 => b(3), A1 => n1546, SL => n83, Z => n832);
   U645 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n833, Z => n1136);
   U646 : MUXB2DL port map( A0 => n1546, A1 => b(1), SL => n83, Z => n833);
   U647 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n834, Z => n1137);
   U648 : MUXB2DL port map( A0 => b(1), A1 => n1548, SL => n83, Z => n834);
   U649 : MUXB2DL port map( A0 => n79, A1 => n81, SL => n835, Z => n1138);
   U650 : NAN2M1D1 port map( A1 => n83, A2 => b(0), Z => n835);
   U651 : NOR2M1D1 port map( A1 => n73, A2 => n76, Z => n1087);
   U652 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n836, Z => n1139);
   U653 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n78, Z => n836);
   U654 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n837, Z => n1140);
   U655 : MUXB2DL port map( A0 => b(12), A1 => n1540, SL => n78, Z => n837);
   U656 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n838, Z => n1141);
   U657 : MUXB2DL port map( A0 => n1540, A1 => n1539, SL => n78, Z => n838);
   U658 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n839, Z => n1142);
   U659 : MUXB2DL port map( A0 => n1539, A1 => n1538, SL => n78, Z => n839);
   U660 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n840, Z => n1143);
   U661 : MUXB2DL port map( A0 => n1538, A1 => b(8), SL => n78, Z => n840);
   U662 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n841, Z => n1144);
   U663 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n78, Z => n841);
   U664 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n842, Z => n1145);
   U665 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n78, Z => n842);
   U666 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n843, Z => n1146);
   U667 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n78, Z => n843);
   U668 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n844, Z => n1147);
   U669 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n78, Z => n844);
   U670 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n845, Z => n1148);
   U671 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n78, Z => n845);
   U672 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n846, Z => n1149);
   U673 : MUXB2DL port map( A0 => b(3), A1 => n1546, SL => n78, Z => n846);
   U674 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n847, Z => n1150);
   U675 : MUXB2DL port map( A0 => n1546, A1 => b(1), SL => n78, Z => n847);
   U676 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n848, Z => n1151);
   U677 : MUXB2DL port map( A0 => b(1), A1 => n1548, SL => n78, Z => n848);
   U678 : MUXB2DL port map( A0 => n73, A1 => n76, SL => n849, Z => n1152);
   U679 : NAN2M1D1 port map( A1 => n78, A2 => n1548, Z => n849);
   U680 : NOR2M1D1 port map( A1 => n66, A2 => n69, Z => n1088);
   U681 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n850, Z => n1153);
   U682 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n71, Z => n850);
   U683 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n851, Z => n1154);
   U684 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n71, Z => n851);
   U685 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n852, Z => n1155);
   U686 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n71, Z => n852);
   U687 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n853, Z => n1156);
   U688 : MUXB2DL port map( A0 => b(12), A1 => n1540, SL => n71, Z => n853);
   U689 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n854, Z => n1157);
   U690 : MUXB2DL port map( A0 => n1540, A1 => n1539, SL => n71, Z => n854);
   U691 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n855, Z => n1158);
   U692 : MUXB2DL port map( A0 => n1539, A1 => n1538, SL => n71, Z => n855);
   U693 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n856, Z => n1159);
   U694 : MUXB2DL port map( A0 => n1538, A1 => b(8), SL => n71, Z => n856);
   U695 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n857, Z => n1160);
   U696 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n71, Z => n857);
   U697 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n858, Z => n1161);
   U698 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n71, Z => n858);
   U699 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n859, Z => n1162);
   U700 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n71, Z => n859);
   U701 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n860, Z => n1163);
   U702 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n71, Z => n860);
   U703 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n861, Z => n1164);
   U704 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n71, Z => n861);
   U705 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n862, Z => n1165);
   U706 : MUXB2DL port map( A0 => b(3), A1 => n1546, SL => n71, Z => n862);
   U707 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n863, Z => n1166);
   U708 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n71, Z => n863);
   U709 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n864, Z => n1167);
   U710 : MUXB2DL port map( A0 => b(1), A1 => n1548, SL => n71, Z => n864);
   U711 : MUXB2DL port map( A0 => n66, A1 => n69, SL => n865, Z => n1168);
   U712 : NAN2M1D1 port map( A1 => n71, A2 => b(0), Z => n865);
   U713 : NOR2M1D1 port map( A1 => n58, A2 => n61, Z => n1089);
   U714 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n866, Z => n1169);
   U715 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n63, Z => n866);
   U716 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n867, Z => n1170);
   U717 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n63, Z => n867);
   U718 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n868, Z => n1171);
   U719 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n63, Z => n868);
   U720 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n869, Z => n1172);
   U721 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n63, Z => n869);
   U722 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n870, Z => n1173);
   U723 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n63, Z => n870);
   U724 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n871, Z => n1174);
   U725 : MUXB2DL port map( A0 => b(12), A1 => n1540, SL => n63, Z => n871);
   U726 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n872, Z => n1175);
   U727 : MUXB2DL port map( A0 => n1540, A1 => n1539, SL => n63, Z => n872);
   U728 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n873, Z => n1176);
   U729 : MUXB2DL port map( A0 => n1539, A1 => n1538, SL => n63, Z => n873);
   U730 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n874, Z => n1177);
   U731 : MUXB2DL port map( A0 => n1538, A1 => b(8), SL => n63, Z => n874);
   U732 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n875, Z => n1178);
   U733 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n63, Z => n875);
   U734 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n876, Z => n1179);
   U735 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n63, Z => n876);
   U736 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n877, Z => n1180);
   U737 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n63, Z => n877);
   U738 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n878, Z => n1181);
   U739 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n63, Z => n878);
   U740 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n879, Z => n1182);
   U741 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n63, Z => n879);
   U742 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n880, Z => n1183);
   U743 : MUXB2DL port map( A0 => b(3), A1 => n1546, SL => n63, Z => n880);
   U744 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n881, Z => n1184);
   U745 : MUXB2DL port map( A0 => n1546, A1 => b(1), SL => n63, Z => n881);
   U746 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n882, Z => n1185);
   U747 : MUXB2DL port map( A0 => b(1), A1 => n1548, SL => n63, Z => n882);
   U748 : MUXB2DL port map( A0 => n58, A1 => n61, SL => n883, Z => n1186);
   U749 : NAN2M1D1 port map( A1 => n63, A2 => b(0), Z => n883);
   U750 : NOR2M1D1 port map( A1 => n50, A2 => n53, Z => n1090);
   U751 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n884, Z => n1187);
   U752 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n56, Z => n884);
   U753 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n885, Z => n1188);
   U754 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n56, Z => n885);
   U755 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n886, Z => n1189);
   U756 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n56, Z => n886);
   U757 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n887, Z => n1190);
   U758 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n56, Z => n887);
   U759 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n888, Z => n1191);
   U760 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n56, Z => n888);
   U761 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n889, Z => n1192);
   U762 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n56, Z => n889);
   U763 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n890, Z => n1193);
   U764 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n56, Z => n890);
   U765 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n891, Z => n1194);
   U766 : MUXB2DL port map( A0 => b(12), A1 => n1540, SL => n56, Z => n891);
   U767 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n892, Z => n1195);
   U768 : MUXB2DL port map( A0 => n1540, A1 => n1539, SL => n56, Z => n892);
   U769 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n893, Z => n1196);
   U770 : MUXB2DL port map( A0 => n1539, A1 => n1538, SL => n56, Z => n893);
   U771 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n894, Z => n1197);
   U772 : MUXB2DL port map( A0 => n1538, A1 => b(8), SL => n56, Z => n894);
   U773 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n895, Z => n1198);
   U774 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n56, Z => n895);
   U775 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n896, Z => n1199);
   U776 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n56, Z => n896);
   U777 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n897, Z => n1200);
   U778 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n56, Z => n897);
   U779 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n898, Z => n1201);
   U780 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n56, Z => n898);
   U781 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n899, Z => n1202);
   U782 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n56, Z => n899);
   U783 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n900, Z => n1203);
   U784 : MUXB2DL port map( A0 => b(3), A1 => n1546, SL => n56, Z => n900);
   U785 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n901, Z => n1204);
   U786 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n56, Z => n901);
   U787 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n902, Z => n1205);
   U788 : MUXB2DL port map( A0 => b(1), A1 => b(0), SL => n56, Z => n902);
   U789 : MUXB2DL port map( A0 => n50, A1 => n53, SL => n903, Z => n1206);
   U790 : NAN2M1D1 port map( A1 => n56, A2 => n1548, Z => n903);
   U791 : NOR2M1D1 port map( A1 => n42, A2 => n45, Z => n1091);
   U792 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n904, Z => n1207);
   U793 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n48, Z => n904);
   U794 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n905, Z => n1208);
   U795 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n48, Z => n905);
   U796 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n906, Z => n1209);
   U797 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n48, Z => n906);
   U798 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n907, Z => n1210);
   U799 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n48, Z => n907);
   U800 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n908, Z => n1211);
   U801 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n48, Z => n908);
   U802 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n909, Z => n1212);
   U803 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n48, Z => n909);
   U804 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n910, Z => n1213);
   U805 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n48, Z => n910);
   U806 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n911, Z => n1214);
   U807 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n48, Z => n911);
   U808 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n912, Z => n1215);
   U809 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n48, Z => n912);
   U810 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n913, Z => n1216);
   U811 : MUXB2DL port map( A0 => b(12), A1 => n1540, SL => n48, Z => n913);
   U812 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n914, Z => n1217);
   U813 : MUXB2DL port map( A0 => n1540, A1 => n1539, SL => n48, Z => n914);
   U814 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n915, Z => n1218);
   U815 : MUXB2DL port map( A0 => n1539, A1 => n1538, SL => n48, Z => n915);
   U816 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n916, Z => n1219);
   U817 : MUXB2DL port map( A0 => n1538, A1 => b(8), SL => n48, Z => n916);
   U818 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n917, Z => n1220);
   U819 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n48, Z => n917);
   U820 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n918, Z => n1221);
   U821 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n48, Z => n918);
   U822 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n919, Z => n1222);
   U823 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n48, Z => n919);
   U824 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n920, Z => n1223);
   U825 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n48, Z => n920);
   U826 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n921, Z => n1224);
   U827 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n48, Z => n921);
   U828 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n922, Z => n1225);
   U829 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n48, Z => n922);
   U830 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n923, Z => n1226);
   U831 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n48, Z => n923);
   U832 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n924, Z => n1227);
   U833 : MUXB2DL port map( A0 => b(1), A1 => b(0), SL => n48, Z => n924);
   U834 : MUXB2DL port map( A0 => n42, A1 => n45, SL => n925, Z => n1228);
   U835 : NAN2M1D1 port map( A1 => n48, A2 => b(0), Z => n925);
   U836 : NOR2M1D1 port map( A1 => n1519, A2 => n38, Z => n1092);
   U837 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n926, Z => n1229);
   U838 : MUXB2DL port map( A0 => b(23), A1 => b(22), SL => n1541, Z => n926);
   U839 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n927, Z => n1230);
   U840 : MUXB2DL port map( A0 => b(22), A1 => b(21), SL => n1541, Z => n927);
   U841 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n928, Z => n1231);
   U842 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n1541, Z => n928);
   U843 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n929, Z => n1232);
   U844 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n1541, Z => n929);
   U845 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n930, Z => n1233);
   U846 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n1541, Z => n930);
   U847 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n931, Z => n1234);
   U848 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n1541, Z => n931);
   U849 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n932, Z => n1235);
   U850 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n1541, Z => n932);
   U851 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n933, Z => n1236);
   U852 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n1541, Z => n933);
   U853 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n934, Z => n1237);
   U854 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n1541, Z => n934);
   U855 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n935, Z => n1238);
   U856 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n1541, Z => n935);
   U857 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n936, Z => n1239);
   U858 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n1541, Z => n936);
   U859 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n937, Z => n1240);
   U860 : MUXB2DL port map( A0 => b(12), A1 => n1540, SL => n1541, Z => n937);
   U861 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n938, Z => n1241);
   U862 : MUXB2DL port map( A0 => n1540, A1 => n1539, SL => n1541, Z => n938);
   U863 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n939, Z => n1242);
   U864 : MUXB2DL port map( A0 => n1539, A1 => n1538, SL => n1541, Z => n939);
   U865 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n940, Z => n1243);
   U866 : MUXB2DL port map( A0 => n1538, A1 => b(8), SL => n1541, Z => n940);
   U867 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n941, Z => n1244);
   U868 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n1541, Z => n941);
   U869 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n942, Z => n1245);
   U870 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n1541, Z => n942);
   U871 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n943, Z => n1246);
   U872 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n1541, Z => n943);
   U873 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n944, Z => n1247);
   U874 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n1541, Z => n944);
   U875 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n945, Z => n1248);
   U876 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n1541, Z => n945);
   U877 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n946, Z => n1249);
   U878 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n1541, Z => n946);
   U879 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n947, Z => n1250);
   U880 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n1541, Z => n947);
   U881 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n948, Z => n1251);
   U882 : MUXB2DL port map( A0 => b(1), A1 => b(0), SL => n1541, Z => n948);
   U883 : MUXB2DL port map( A0 => n1519, A1 => n38, SL => n949, Z => n1252);
   U884 : NAN2M1D1 port map( A1 => n1541, A2 => b(0), Z => n949);
   U886 : MUXB2DL port map( A0 => n1543, A1 => n30, SL => n950, Z => n1253);
   U887 : MUXB2DL port map( A0 => b(25), A1 => b(24), SL => n1542, Z => n950);
   U888 : MUXB2DL port map( A0 => n1543, A1 => n30, SL => n951, Z => n1254);
   U889 : MUXB2DL port map( A0 => b(24), A1 => b(23), SL => n1542, Z => n951);
   U890 : MUXB2DL port map( A0 => n1543, A1 => n30, SL => n952, Z => n1255);
   U891 : MUXB2DL port map( A0 => b(23), A1 => b(22), SL => n1542, Z => n952);
   U892 : MUXB2DL port map( A0 => n1543, A1 => n30, SL => n953, Z => n1256);
   U893 : MUXB2DL port map( A0 => b(22), A1 => b(21), SL => n1542, Z => n953);
   U894 : MUXB2DL port map( A0 => n1543, A1 => n30, SL => n954, Z => n1257);
   U895 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n1542, Z => n954);
   U896 : MUXB2DL port map( A0 => n1543, A1 => n30, SL => n955, Z => n1258);
   U897 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n1542, Z => n955);
   U898 : MUXB2DL port map( A0 => n1543, A1 => n30, SL => n956, Z => n1259);
   U899 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n1542, Z => n956);
   U900 : MUXB2DL port map( A0 => n1543, A1 => n30, SL => n957, Z => n1260);
   U901 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n1542, Z => n957);
   U902 : MUXB2DL port map( A0 => n1543, A1 => n30, SL => n958, Z => n1261);
   U903 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n1542, Z => n958);
   U904 : MUXB2DL port map( A0 => n1543, A1 => n30, SL => n959, Z => n1262);
   U905 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n1542, Z => n959);
   U906 : MUXB2DL port map( A0 => n1543, A1 => n30, SL => n960, Z => n1263);
   U907 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n1542, Z => n960);
   U908 : MUXB2DL port map( A0 => n1543, A1 => n30, SL => n961, Z => n1264);
   U909 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n1542, Z => n961);
   U910 : MUXB2DL port map( A0 => n1543, A1 => n30, SL => n962, Z => n1265);
   U911 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n1542, Z => n962);
   U912 : MUXB2DL port map( A0 => n1543, A1 => n30, SL => n963, Z => n1266);
   U913 : MUXB2DL port map( A0 => b(12), A1 => n1540, SL => n1542, Z => n963);
   U914 : MUXB2DL port map( A0 => n1543, A1 => n30, SL => n964, Z => n1267);
   U915 : MUXB2DL port map( A0 => n1540, A1 => n1539, SL => n1542, Z => n964);
   U916 : MUXB2DL port map( A0 => n1543, A1 => n30, SL => n965, Z => n1268);
   U917 : MUXB2DL port map( A0 => n1539, A1 => n1538, SL => n1542, Z => n965);
   U918 : MUXB2DL port map( A0 => n1543, A1 => n30, SL => n966, Z => n1269);
   U919 : MUXB2DL port map( A0 => n1538, A1 => b(8), SL => n1542, Z => n966);
   U920 : MUXB2DL port map( A0 => n1543, A1 => n30, SL => n967, Z => n1270);
   U921 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n1542, Z => n967);
   U922 : MUXB2DL port map( A0 => n1543, A1 => n30, SL => n968, Z => n1271);
   U923 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n1542, Z => n968);
   U924 : MUXB2DL port map( A0 => n1543, A1 => n30, SL => n969, Z => n1272);
   U925 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n1542, Z => n969);
   U926 : MUXB2DL port map( A0 => n1543, A1 => n30, SL => n970, Z => n1273);
   U927 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n1542, Z => n970);
   U928 : MUXB2DL port map( A0 => n1543, A1 => n30, SL => n971, Z => n1274);
   U929 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n1542, Z => n971);
   U930 : MUXB2DL port map( A0 => n1543, A1 => n30, SL => n972, Z => n1275);
   U931 : MUXB2DL port map( A0 => b(3), A1 => b(2), SL => n1542, Z => n972);
   U932 : MUXB2DL port map( A0 => n1543, A1 => n30, SL => n973, Z => n1276);
   U933 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n1542, Z => n973);
   U934 : MUXB2DL port map( A0 => n1543, A1 => n30, SL => n974, Z => n1277);
   U935 : MUXB2DL port map( A0 => b(1), A1 => b(0), SL => n1542, Z => n974);
   U936 : MUXB2DL port map( A0 => n1543, A1 => n30, SL => n975, Z => n1278);
   U937 : NAN2M1D1 port map( A1 => n1542, A2 => b(0), Z => n975);
   U938 : NOR2M1D1 port map( A1 => n1518, A2 => n22, Z => n1094);
   U939 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n976, Z => n1279);
   U940 : MUXB2DL port map( A0 => b(27), A1 => b(26), SL => n1544, Z => n976);
   U941 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n977, Z => n1280);
   U942 : MUXB2DL port map( A0 => b(26), A1 => b(25), SL => n1544, Z => n977);
   U943 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n978, Z => n1281);
   U944 : MUXB2DL port map( A0 => b(25), A1 => b(24), SL => n1544, Z => n978);
   U945 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n979, Z => n1282);
   U946 : MUXB2DL port map( A0 => b(24), A1 => b(23), SL => n1544, Z => n979);
   U947 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n980, Z => n1283);
   U948 : MUXB2DL port map( A0 => b(23), A1 => b(22), SL => n1544, Z => n980);
   U949 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n981, Z => n1284);
   U950 : MUXB2DL port map( A0 => b(22), A1 => b(21), SL => n1544, Z => n981);
   U951 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n982, Z => n1285);
   U952 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n1544, Z => n982);
   U953 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n983, Z => n1286);
   U954 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n1544, Z => n983);
   U955 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n984, Z => n1287);
   U956 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n1544, Z => n984);
   U957 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n985, Z => n1288);
   U958 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n1544, Z => n985);
   U959 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n986, Z => n1289);
   U960 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n1544, Z => n986);
   U961 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n987, Z => n1290);
   U962 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n1544, Z => n987);
   U963 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n988, Z => n1291);
   U964 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n1544, Z => n988);
   U965 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n989, Z => n1292);
   U966 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n1544, Z => n989);
   U967 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n990, Z => n1293);
   U968 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n1544, Z => n990);
   U969 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n991, Z => n1294);
   U970 : MUXB2DL port map( A0 => b(12), A1 => n1540, SL => n1544, Z => n991);
   U971 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n992, Z => n1295);
   U972 : MUXB2DL port map( A0 => n1540, A1 => n1539, SL => n1544, Z => n992);
   U973 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n993, Z => n1296);
   U974 : MUXB2DL port map( A0 => n1539, A1 => n1538, SL => n1544, Z => n993);
   U975 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n994, Z => n1297);
   U976 : MUXB2DL port map( A0 => n1538, A1 => b(8), SL => n1544, Z => n994);
   U977 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n995, Z => n1298);
   U978 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n1544, Z => n995);
   U979 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n996, Z => n1299);
   U980 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n1544, Z => n996);
   U981 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n997, Z => n1300);
   U982 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n1544, Z => n997);
   U983 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n998, Z => n1301);
   U984 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n1544, Z => n998);
   U985 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n999, Z => n1302);
   U986 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n1544, Z => n999);
   U987 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n1000, Z => n1303);
   U988 : MUXB2DL port map( A0 => b(3), A1 => n1546, SL => n1544, Z => n1000);
   U989 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n1001, Z => n1304);
   U990 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n1544, Z => n1001);
   U991 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n1002, Z => n1305);
   U992 : MUXB2DL port map( A0 => b(1), A1 => n1548, SL => n1544, Z => n1002);
   U993 : MUXB2DL port map( A0 => n1518, A1 => n22, SL => n1003, Z => n1306);
   U994 : NAN2M1D1 port map( A1 => n1544, A2 => b(0), Z => n1003);
   U995 : NOR2M1D1 port map( A1 => n1517, A2 => n14, Z => n1095);
   U996 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1004, Z => n1307);
   U997 : MUXB2DL port map( A0 => b(29), A1 => b(28), SL => n1545, Z => n1004);
   U998 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1005, Z => n1308);
   U999 : MUXB2DL port map( A0 => b(28), A1 => b(27), SL => n1545, Z => n1005);
   U1000 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1006, Z => n1309);
   U1001 : MUXB2DL port map( A0 => b(27), A1 => b(26), SL => n1545, Z => n1006)
                           ;
   U1002 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1007, Z => n1310);
   U1003 : MUXB2DL port map( A0 => b(26), A1 => b(25), SL => n1545, Z => n1007)
                           ;
   U1004 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1008, Z => n1311);
   U1005 : MUXB2DL port map( A0 => b(25), A1 => b(24), SL => n1545, Z => n1008)
                           ;
   U1006 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1009, Z => n1312);
   U1007 : MUXB2DL port map( A0 => b(24), A1 => b(23), SL => n1545, Z => n1009)
                           ;
   U1008 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1010, Z => n1313);
   U1009 : MUXB2DL port map( A0 => b(23), A1 => b(22), SL => n1545, Z => n1010)
                           ;
   U1010 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1011, Z => n1314);
   U1011 : MUXB2DL port map( A0 => b(22), A1 => b(21), SL => n1545, Z => n1011)
                           ;
   U1012 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1012, Z => n1315);
   U1013 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n1545, Z => n1012)
                           ;
   U1014 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1013, Z => n1316);
   U1015 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n1545, Z => n1013)
                           ;
   U1016 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1014, Z => n1317);
   U1017 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n1545, Z => n1014)
                           ;
   U1018 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1015, Z => n1318);
   U1019 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n1545, Z => n1015)
                           ;
   U1020 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1016, Z => n1319);
   U1021 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n1545, Z => n1016)
                           ;
   U1022 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1017, Z => n1320);
   U1023 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n1545, Z => n1017)
                           ;
   U1024 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1018, Z => n1321);
   U1025 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n1545, Z => n1018)
                           ;
   U1026 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1019, Z => n1322);
   U1027 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n1545, Z => n1019)
                           ;
   U1028 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1020, Z => n1323);
   U1029 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n1545, Z => n1020)
                           ;
   U1030 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1021, Z => n1324);
   U1031 : MUXB2DL port map( A0 => b(12), A1 => n1540, SL => n1545, Z => n1021)
                           ;
   U1032 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1022, Z => n1325);
   U1033 : MUXB2DL port map( A0 => n1540, A1 => n1539, SL => n1545, Z => n1022)
                           ;
   U1034 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1023, Z => n1326);
   U1035 : MUXB2DL port map( A0 => n1539, A1 => n1538, SL => n1545, Z => n1023)
                           ;
   U1036 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1024, Z => n1327);
   U1037 : MUXB2DL port map( A0 => n1538, A1 => b(8), SL => n1545, Z => n1024);
   U1038 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1025, Z => n1328);
   U1039 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n1545, Z => n1025);
   U1040 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1026, Z => n1329);
   U1041 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n1545, Z => n1026);
   U1042 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1027, Z => n1330);
   U1043 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n1545, Z => n1027);
   U1044 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1028, Z => n1331);
   U1045 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n1545, Z => n1028);
   U1046 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1029, Z => n1332);
   U1047 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n1545, Z => n1029);
   U1048 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1030, Z => n1333);
   U1049 : MUXB2DL port map( A0 => b(3), A1 => n1546, SL => n1545, Z => n1030);
   U1050 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1031, Z => n1334);
   U1051 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n1545, Z => n1031);
   U1052 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1032, Z => n1335);
   U1053 : MUXB2DL port map( A0 => b(1), A1 => n1548, SL => n1545, Z => n1032);
   U1054 : MUXB2DL port map( A0 => n1517, A1 => n14, SL => n1033, Z => n1336);
   U1055 : NAN2M1D1 port map( A1 => n1545, A2 => b(0), Z => n1033);
   U1056 : NOR2M1D1 port map( A1 => n3, A2 => n6, Z => n1096);
   U1057 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1034, Z => n1337);
   U1058 : MUXB2DL port map( A0 => b(31), A1 => b(30), SL => n8, Z => n1034);
   U1059 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1035, Z => n1338);
   U1060 : MUXB2DL port map( A0 => b(30), A1 => b(29), SL => n8, Z => n1035);
   U1061 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1036, Z => n1339);
   U1062 : MUXB2DL port map( A0 => b(29), A1 => b(28), SL => n8, Z => n1036);
   U1063 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1037, Z => n1340);
   U1064 : MUXB2DL port map( A0 => b(28), A1 => b(27), SL => n8, Z => n1037);
   U1065 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1038, Z => n1341);
   U1066 : MUXB2DL port map( A0 => b(27), A1 => b(26), SL => n8, Z => n1038);
   U1067 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1039, Z => n1342);
   U1068 : MUXB2DL port map( A0 => b(26), A1 => b(25), SL => n8, Z => n1039);
   U1069 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1040, Z => n1343);
   U1070 : MUXB2DL port map( A0 => b(25), A1 => b(24), SL => n8, Z => n1040);
   U1071 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1041, Z => n1344);
   U1072 : MUXB2DL port map( A0 => b(24), A1 => b(23), SL => n8, Z => n1041);
   U1073 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1042, Z => n1345);
   U1074 : MUXB2DL port map( A0 => b(23), A1 => b(22), SL => n8, Z => n1042);
   U1075 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1043, Z => n1346);
   U1076 : MUXB2DL port map( A0 => b(22), A1 => b(21), SL => n8, Z => n1043);
   U1077 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1044, Z => n1347);
   U1078 : MUXB2DL port map( A0 => b(21), A1 => b(20), SL => n8, Z => n1044);
   U1079 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1045, Z => n1348);
   U1080 : MUXB2DL port map( A0 => b(20), A1 => b(19), SL => n8, Z => n1045);
   U1081 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1046, Z => n1349);
   U1082 : MUXB2DL port map( A0 => b(19), A1 => b(18), SL => n8, Z => n1046);
   U1083 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1047, Z => n1350);
   U1084 : MUXB2DL port map( A0 => b(18), A1 => b(17), SL => n8, Z => n1047);
   U1085 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1048, Z => n1351);
   U1086 : MUXB2DL port map( A0 => b(17), A1 => b(16), SL => n8, Z => n1048);
   U1087 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1049, Z => n1352);
   U1088 : MUXB2DL port map( A0 => b(16), A1 => b(15), SL => n8, Z => n1049);
   U1089 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1050, Z => n1353);
   U1090 : MUXB2DL port map( A0 => b(15), A1 => b(14), SL => n8, Z => n1050);
   U1091 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1051, Z => n1354);
   U1092 : MUXB2DL port map( A0 => b(14), A1 => b(13), SL => n8, Z => n1051);
   U1093 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1052, Z => n1355);
   U1094 : MUXB2DL port map( A0 => b(13), A1 => b(12), SL => n8, Z => n1052);
   U1095 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1053, Z => n1356);
   U1096 : MUXB2DL port map( A0 => b(12), A1 => n1540, SL => n8, Z => n1053);
   U1097 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1054, Z => n1357);
   U1098 : MUXB2DL port map( A0 => n1540, A1 => n1539, SL => n8, Z => n1054);
   U1099 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1055, Z => n1358);
   U1100 : MUXB2DL port map( A0 => n1539, A1 => n1538, SL => n8, Z => n1055);
   U1101 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1056, Z => n1359);
   U1102 : MUXB2DL port map( A0 => n1538, A1 => b(8), SL => n8, Z => n1056);
   U1103 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1057, Z => n1360);
   U1104 : MUXB2DL port map( A0 => b(8), A1 => b(7), SL => n8, Z => n1057);
   U1105 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1058, Z => n1361);
   U1106 : MUXB2DL port map( A0 => b(7), A1 => b(6), SL => n8, Z => n1058);
   U1107 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1059, Z => n1362);
   U1108 : MUXB2DL port map( A0 => b(6), A1 => b(5), SL => n8, Z => n1059);
   U1109 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1060, Z => n1363);
   U1110 : MUXB2DL port map( A0 => b(5), A1 => b(4), SL => n8, Z => n1060);
   U1111 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1061, Z => n1364);
   U1112 : MUXB2DL port map( A0 => b(4), A1 => b(3), SL => n8, Z => n1061);
   U1113 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1062, Z => n1365);
   U1114 : MUXB2DL port map( A0 => b(3), A1 => n1546, SL => n8, Z => n1062);
   U1115 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1063, Z => n1366);
   U1116 : MUXB2DL port map( A0 => b(2), A1 => b(1), SL => n8, Z => n1063);
   U1117 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1064, Z => n1367);
   U1118 : MUXB2DL port map( A0 => b(1), A1 => n1548, SL => n8, Z => n1064);
   U1119 : MUXB2DL port map( A0 => n3, A1 => n6, SL => n1065, Z => n1368);
   U1120 : NAN2M1D1 port map( A1 => n8, A2 => n1548, Z => n1065);
   U1121 : OAI21D1 port map( A1 => a(29), A2 => a(30), B => n1066, Z => n104);
   U1123 : EXNOR2D1 port map( A1 => a(29), A2 => a(30), Z => n106);
   U1125 : OAI21D1 port map( A1 => a(27), A2 => a(28), B => n1067, Z => n99);
   U1127 : EXNOR2D1 port map( A1 => a(27), A2 => a(28), Z => n103);
   U1129 : OAI21D1 port map( A1 => a(25), A2 => a(26), B => n1068, Z => n94);
   U1131 : EXNOR2D1 port map( A1 => a(25), A2 => a(26), Z => n98);
   U1135 : EXNOR2D1 port map( A1 => a(23), A2 => a(24), Z => n93);
   U1186 : ADHALFDL port map( A => n1278, B => n1093, CO => n780, S => n781);
   U1187 : OAI21D1 port map( A1 => a(1), A2 => a(2), B => n1080, Z => n1517);
   U1188 : OAI21D1 port map( A1 => a(3), A2 => a(4), B => n1079, Z => n1518);
   U1189 : OAI21D1 port map( A1 => a(7), A2 => a(8), B => n1077, Z => n1519);
   U1190 : AND2D1 port map( A1 => n1522, A2 => n305, Z => product(0));
   U1191 : AO21D1 port map( A1 => n215, A2 => n187, B => n188, Z => n1521);
   U1192 : OR2D1 port map( A1 => n1368, A2 => n1096, Z => n1522);
   U1193 : OA21M20D1 port map( A1 => n1523, A2 => n197, B => n194, Z => n190);
   U1194 : INVD1 port map( A => n215, Z => n214);
   U1195 : INVD1 port map( A => n233, Z => n232);
   U1196 : NAN2D1 port map( A1 => n313, A2 => n231, Z => n162);
   U1197 : INVD1 port map( A => n242, Z => n241);
   U1198 : INVD1 port map( A => n255, Z => n254);
   U1199 : INVD1 port map( A => n230, Z => n313);
   U1200 : INVD1 port map( A => n231, Z => n229);
   U1201 : INVD1 port map( A => n264, Z => n263);
   U1202 : NAN2D1 port map( A1 => n223, A2 => n1528, Z => n216);
   U1203 : INVD1 port map( A => n221, Z => n219);
   U1204 : NAN2D1 port map( A1 => n1530, A2 => n1529, Z => n243);
   U1205 : INVD1 port map( A => n248, Z => n246);
   U1206 : NAN2D1 port map( A1 => n1524, A2 => n1527, Z => n265);
   U1207 : INVD1 port map( A => n270, Z => n268);
   U1208 : NOR2D1 port map( A1 => n258, A2 => n261, Z => n256);
   U1209 : NOR2D1 port map( A1 => n236, A2 => n239, Z => n234);
   U1210 : NOR2D1 port map( A1 => n189, A2 => n201, Z => n187);
   U1211 : INVD1 port map( A => n209, Z => n211);
   U1212 : INVD1 port map( A => n206, Z => n204);
   U1213 : INVD1 port map( A => n275, Z => n273);
   U1214 : OR2D1 port map( A1 => n553, A2 => n574, Z => n1523);
   U1215 : NAN2D1 port map( A1 => n1523, A2 => n1526, Z => n189);
   U1216 : INVD1 port map( A => n199, Z => n197);
   U1217 : INVD1 port map( A => n253, Z => n251);
   U1218 : NAN2D1 port map( A1 => n667, A2 => n682, Z => n231);
   U1219 : NOR2D1 port map( A1 => n225, A2 => n230, Z => n223);
   U1220 : NAN2D1 port map( A1 => n1525, A2 => n310, Z => n201);
   U1221 : NOR2D1 port map( A1 => n683, A2 => n696, Z => n236);
   U1222 : NAN2D1 port map( A1 => n553, A2 => n574, Z => n194);
   U1223 : INVD1 port map( A => n208, Z => n310);
   U1224 : NOR2D1 port map( A1 => n667, A2 => n682, Z => n230);
   U1225 : NAN2D1 port map( A1 => n683, A2 => n696, Z => n237);
   U1226 : NAN2D1 port map( A1 => n1523, A2 => n194, Z => n156);
   U1227 : NAN2D1 port map( A1 => n1526, A2 => n199, Z => n157);
   U1228 : NAN2D1 port map( A1 => n1525, A2 => n206, Z => n158);
   U1229 : NAN2D1 port map( A1 => n310, A2 => n209, Z => n159);
   U1230 : NAN2D1 port map( A1 => n312, A2 => n226, Z => n161);
   U1231 : INVD1 port map( A => n225, Z => n312);
   U1232 : NAN2D1 port map( A1 => n1528, A2 => n221, Z => n160);
   U1233 : NAN2D1 port map( A1 => n314, A2 => n237, Z => n163);
   U1234 : INVD1 port map( A => n236, Z => n314);
   U1235 : NAN2D1 port map( A1 => n1530, A2 => n248, Z => n165);
   U1236 : NAN2D1 port map( A1 => n315, A2 => n240, Z => n164);
   U1237 : INVD1 port map( A => n239, Z => n315);
   U1238 : NAN2D1 port map( A1 => n1529, A2 => n253, Z => n166);
   U1239 : NAN2D1 port map( A1 => n318, A2 => n259, Z => n167);
   U1240 : INVD1 port map( A => n258, Z => n318);
   U1241 : NAN2D1 port map( A1 => n319, A2 => n262, Z => n168);
   U1242 : INVD1 port map( A => n261, Z => n319);
   U1243 : INVD1 port map( A => n277, Z => n276);
   U1244 : NAN2D1 port map( A1 => n1524, A2 => n270, Z => n169);
   U1245 : NAN2D1 port map( A1 => n1527, A2 => n275, Z => n170);
   U1246 : INVD1 port map( A => n286, Z => n285);
   U1247 : OR2D1 port map( A1 => n755, A2 => n762, Z => n1524);
   U1248 : NAN2D1 port map( A1 => n755, A2 => n762, Z => n270);
   U1249 : NOR2D1 port map( A1 => n280, A2 => n283, Z => n278);
   U1250 : OA21M20D1 port map( A1 => n1531, A2 => n294, B => n293, Z => n289);
   U1251 : NOR2D1 port map( A1 => n651, A2 => n666, Z => n225);
   U1252 : OA21M20D1 port map( A1 => n1532, A2 => n302, B => n301, Z => n297);
   U1253 : OR2D1 port map( A1 => n595, A2 => n614, Z => n1525);
   U1254 : NOR2D1 port map( A1 => n771, A2 => n776, Z => n280);
   U1255 : NOR2D1 port map( A1 => n745, A2 => n754, Z => n261);
   U1256 : NOR2D1 port map( A1 => n735, A2 => n744, Z => n258);
   U1257 : NAN2D1 port map( A1 => n763, A2 => n770, Z => n275);
   U1258 : OR2D1 port map( A1 => n575, A2 => n594, Z => n1526);
   U1259 : NAN2D1 port map( A1 => n575, A2 => n594, Z => n199);
   U1260 : NAN2D1 port map( A1 => n723, A2 => n734, Z => n253);
   U1261 : NAN2D1 port map( A1 => n651, A2 => n666, Z => n226);
   U1262 : OR2D1 port map( A1 => n763, A2 => n770, Z => n1527);
   U1263 : NAN2D1 port map( A1 => n595, A2 => n614, Z => n206);
   U1264 : OR2D1 port map( A1 => n633, A2 => n650, Z => n1528);
   U1265 : NAN2D1 port map( A1 => n745, A2 => n754, Z => n262);
   U1266 : OR2D1 port map( A1 => n723, A2 => n734, Z => n1529);
   U1267 : NAN2D1 port map( A1 => n615, A2 => n632, Z => n209);
   U1268 : OR2D1 port map( A1 => n711, A2 => n722, Z => n1530);
   U1269 : NAN2D1 port map( A1 => n771, A2 => n776, Z => n281);
   U1270 : NOR2D1 port map( A1 => n615, A2 => n632, Z => n208);
   U1271 : NAN2D1 port map( A1 => n735, A2 => n744, Z => n259);
   U1272 : NOR2D1 port map( A1 => n697, A2 => n710, Z => n239);
   U1273 : NAN2D1 port map( A1 => n633, A2 => n650, Z => n221);
   U1274 : NAN2D1 port map( A1 => n711, A2 => n722, Z => n248);
   U1275 : NAN2D1 port map( A1 => n697, A2 => n710, Z => n240);
   U1276 : NAN2D1 port map( A1 => n322, A2 => n281, Z => n171);
   U1277 : INVD1 port map( A => n280, Z => n322);
   U1278 : NAN2D1 port map( A1 => n323, A2 => n284, Z => n172);
   U1279 : INVD1 port map( A => n283, Z => n323);
   U1280 : NAN2D1 port map( A1 => n324, A2 => n288, Z => n173);
   U1281 : INVD1 port map( A => n287, Z => n324);
   U1282 : NAN2D1 port map( A1 => n1531, A2 => n293, Z => n174);
   U1283 : NAN2D1 port map( A1 => n326, A2 => n296, Z => n175);
   U1284 : INVD1 port map( A => n295, Z => n326);
   U1285 : NAN2D1 port map( A1 => n1532, A2 => n301, Z => n176);
   U1286 : OR2D1 port map( A1 => n787, A2 => n789, Z => n1531);
   U1287 : OR2D1 port map( A1 => n793, A2 => n1366, Z => n1532);
   U1288 : NOR2D1 port map( A1 => n777, A2 => n782, Z => n283);
   U1289 : NAN2D1 port map( A1 => n787, A2 => n789, Z => n293);
   U1290 : NAN2D1 port map( A1 => n793, A2 => n1366, Z => n301);
   U1291 : NAN2D1 port map( A1 => n777, A2 => n782, Z => n284);
   U1292 : NOR2D1 port map( A1 => n783, A2 => n786, Z => n287);
   U1293 : NOR2D1 port map( A1 => n791, A2 => n792, Z => n295);
   U1294 : NAN2D1 port map( A1 => n783, A2 => n786, Z => n288);
   U1295 : NAN2D1 port map( A1 => n791, A2 => n792, Z => n296);
   U1296 : NAN2D1 port map( A1 => n1368, A2 => n1096, Z => n305);
   U1297 : NOR2D1 port map( A1 => n303, A2 => n305, Z => n302);
   U1298 : EXOR2D1 port map( A1 => n178, A2 => n155, Z => product(31));
   U1299 : EXOR2D1 port map( A1 => n329, A2 => n344, Z => n155);
   U1300 : ADHALFDL port map( A => n1335, B => n1365, CO => n790, S => n791);
   U1301 : INVD1 port map( A => n1533, Z => n1545);
   U1302 : ADHALFDL port map( A => n1336, B => n1095, CO => n792, S => n793);
   U1303 : NOR2D1 port map( A1 => n1537, A2 => n30, Z => n1093);
   U1304 : INVD1 port map( A => n1535, Z => n1544);
   U1305 : ADHALFDL port map( A => n1331, B => n1361, CO => n774, S => n775);
   U1306 : INVD1 port map( A => n1534, Z => n1542);
   U1307 : ADHALFDL port map( A => n1252, B => n1092, CO => n768, S => n769);
   U1308 : INVD1 port map( A => n1536, Z => n1541);
   U1309 : ADHALFDL port map( A => n1333, B => n1363, CO => n784, S => n785);
   U1310 : ADHALFDL port map( A => n1306, B => n1094, CO => n788, S => n789);
   U1311 : INVD1 port map( A => n1537, Z => n1543);
   U1312 : ADHALFDL port map( A => n1206, B => n1090, CO => n732, S => n733);
   U1313 : ADHALFDL port map( A => n1168, B => n1088, CO => n680, S => n681);
   U1314 : ADHALFDL port map( A => n1152, B => n1087, CO => n648, S => n649);
   U1315 : ADHALFDL port map( A => n1228, B => n1091, CO => n752, S => n753);
   U1316 : ADHALFDL port map( A => n1186, B => n1089, CO => n708, S => n709);
   U1317 : ADHALFDL port map( A => n1138, B => n1086, CO => n612, S => n613);
   U1318 : INVD1 port map( A => n1367, Z => n303);
   U1319 : ADHALFDL port map( A => n1126, B => n1085, CO => n572, S => n573);
   U1320 : ADHALFDL port map( A => n1116, B => n1084, CO => n528, S => n529);
   U1321 : ADHALFDL port map( A => n1108, B => n1083, CO => n480, S => n481);
   U1322 : ADHALFDL port map( A => n1102, B => n1082, CO => n428, S => n429);
   U1323 : ADHALFDL port map( A => n1098, B => n1081, CO => n372, S => n373);
   U1324 : ADHALFDL port map( A => n1329, B => n1359, CO => n760, S => n761);
   U1325 : EXOR2D1 port map( A1 => a(1), A2 => a(2), Z => n1533);
   U1326 : ADHALFDL port map( A => n1323, B => n1353, CO => n694, S => n695);
   U1327 : EXOR2D1 port map( A1 => a(5), A2 => a(6), Z => n1534);
   U1328 : EXOR2D1 port map( A1 => a(3), A2 => a(4), Z => n1535);
   U1329 : EXOR2D1 port map( A1 => a(7), A2 => a(8), Z => n1536);
   U1330 : ADHALFDL port map( A => n1317, B => n1347, CO => n592, S => n593);
   U1331 : ADHALFDL port map( A => n1327, B => n1357, CO => n742, S => n743);
   U1332 : ADHALFDL port map( A => n1319, B => n1349, CO => n630, S => n631);
   U1333 : ADHALFDL port map( A => n1321, B => n1351, CO => n664, S => n665);
   U1334 : ADHALFDL port map( A => n1325, B => n1355, CO => n720, S => n721);
   U1335 : OA21D1 port map( A1 => a(5), A2 => a(6), B => n1078, Z => n1537);
   U1336 : INVD1 port map( A => a(3), Z => n1080);
   U1337 : EXNOR2D1 port map( A1 => a(11), A2 => a(12), Z => n56);
   U1338 : INVD1 port map( A => a(7), Z => n1078);
   U1339 : NAN2D1 port map( A1 => a(0), A2 => n6, Z => n3);
   U1340 : INVD1 port map( A => a(1), Z => n6);
   U1341 : INVD1 port map( A => a(9), Z => n1077);
   U1342 : EXNOR2D1 port map( A1 => a(13), A2 => a(14), Z => n63);
   U1343 : EXNOR2D1 port map( A1 => a(15), A2 => a(16), Z => n71);
   U1344 : INVD1 port map( A => a(5), Z => n1079);
   U1345 : EXNOR2D1 port map( A1 => a(9), A2 => a(10), Z => n48);
   U1346 : EXNOR2D1 port map( A1 => a(17), A2 => a(18), Z => n78);
   U1347 : AO21D1 port map( A1 => a(1), A2 => a(2), B => n1080, Z => n14);
   U1348 : INVD1 port map( A => n1547, Z => n1546);
   U1349 : INVD1 port map( A => n1549, Z => n1548);
   U1350 : AO21D1 port map( A1 => a(5), A2 => a(6), B => n1078, Z => n30);
   U1351 : EXNOR2D1 port map( A1 => a(19), A2 => a(20), Z => n83);
   U1352 : INVD1 port map( A => a(0), Z => n8);
   U1353 : AO21D1 port map( A1 => a(11), A2 => a(12), B => n1075, Z => n53);
   U1354 : INVD1 port map( A => a(13), Z => n1075);
   U1355 : ADHALFDL port map( A => n1315, B => n1345, CO => n550, S => n551);
   U1356 : AO21D1 port map( A1 => a(3), A2 => a(4), B => n1079, Z => n22);
   U1357 : AO21D1 port map( A1 => a(7), A2 => a(8), B => n1077, Z => n38);
   U1358 : OAI21D1 port map( A1 => a(11), A2 => a(12), B => n1075, Z => n50);
   U1359 : AO21D1 port map( A1 => a(13), A2 => a(14), B => n1074, Z => n61);
   U1360 : AO21D1 port map( A1 => a(15), A2 => a(16), B => n1073, Z => n69);
   U1361 : INVD1 port map( A => a(15), Z => n1074);
   U1362 : OAI21D1 port map( A1 => a(13), A2 => a(14), B => n1074, Z => n58);
   U1363 : INVD1 port map( A => a(17), Z => n1073);
   U1364 : OAI21D1 port map( A1 => a(15), A2 => a(16), B => n1073, Z => n66);
   U1365 : AO21D1 port map( A1 => a(9), A2 => a(10), B => n1076, Z => n45);
   U1366 : INVD1 port map( A => a(11), Z => n1076);
   U1367 : OAI21D1 port map( A1 => a(17), A2 => a(18), B => n1072, Z => n73);
   U1368 : INVD1 port map( A => a(19), Z => n1072);
   U1369 : OAI21D1 port map( A1 => a(9), A2 => a(10), B => n1076, Z => n42);
   U1370 : AO21D1 port map( A1 => a(17), A2 => a(18), B => n1072, Z => n76);
   U1371 : EXNOR2D1 port map( A1 => a(21), A2 => a(22), Z => n88);
   U1372 : OAI21D1 port map( A1 => a(19), A2 => a(20), B => n1071, Z => n79);
   U1373 : INVD1 port map( A => a(21), Z => n1071);
   U1374 : AO21D1 port map( A1 => a(19), A2 => a(20), B => n1071, Z => n81);
   U1375 : OAI21D1 port map( A1 => a(21), A2 => a(22), B => n1070, Z => n84);
   U1376 : INVD1 port map( A => a(23), Z => n1070);
   U1377 : AO21D1 port map( A1 => a(21), A2 => a(22), B => n1070, Z => n86);
   U1378 : ADHALFDL port map( A => n1313, B => n1343, CO => n504, S => n505);
   U1379 : OAI21D1 port map( A1 => a(23), A2 => a(24), B => n1069, Z => n89);
   U1380 : ADHALFDL port map( A => n1311, B => n1341, CO => n454, S => n455);
   U1381 : INVD1 port map( A => a(25), Z => n1069);
   U1382 : AO21D1 port map( A1 => a(23), A2 => a(24), B => n1069, Z => n91);
   U1383 : ADHALFDL port map( A => n1309, B => n1339, CO => n400, S => n401);
   U1384 : AO21D1 port map( A1 => a(25), A2 => a(26), B => n1068, Z => n96);
   U1385 : INVD1 port map( A => a(27), Z => n1068);
   U1386 : EXOR2D1 port map( A1 => n1307, A2 => n1337, Z => n343);
   U1387 : AO21D1 port map( A1 => a(27), A2 => a(28), B => n1067, Z => n101);
   U1388 : INVD1 port map( A => a(29), Z => n1067);
   U1389 : AO21D1 port map( A1 => a(29), A2 => a(30), B => n1066, Z => n105);
   U1390 : INVD1 port map( A => b(2), Z => n1547);
   U1391 : INVD1 port map( A => b(0), Z => n1549);
   U1392 : BUFD1 port map( A => b(9), Z => n1538);
   U1393 : BUFD1 port map( A => b(10), Z => n1539);
   U1394 : BUFD1 port map( A => b(11), Z => n1540);
   U1395 : INVD1 port map( A => a(31), Z => n1066);

end hier_filter_none_5;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_gp_custom.all;

architecture hier_filter_none_5 of gp_custom is

   component NOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN4D1
      port( A1, A2, A3, A4 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AO22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2DL
      port( A0, A1, SL : in std_logic;  Z : out std_logic);
   end component;
   
   component AO31D1
      port( A1, A2, A3, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22M10D1
      port( B1, B2, A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3M1D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211D1
      port( A1, A2, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2D1
      port( A0, A1, SL : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFRPQ1
      port( D, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component DFERPQ1
      port( D, CEB, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFSPQ1
      port( D, CK, SB : in std_logic;  Q : out std_logic);
   end component;
   
   component gp_custom_DW_mult_tc_9
      port( a, b : in std_logic_vector (31 downto 0);  product : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component gp_custom_DW_mult_tc_8
      port( a, b : in std_logic_vector (31 downto 0);  product : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component gp_custom_DW_mult_tc_7
      port( a, b : in std_logic_vector (31 downto 0);  product : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component gp_custom_DW_mult_tc_6
      port( a, b : in std_logic_vector (31 downto 0);  product : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component gp_custom_DW_mult_tc_5
      port( a, b : in std_logic_vector (31 downto 0);  product : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component OA21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI32D1
      port( A1, A2, A3, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal N62, N63, N64, avs_readdata_31_port, avs_readdata_30_port, 
      avs_readdata_29_port, avs_readdata_28_port, avs_readdata_27_port, 
      avs_readdata_26_port, avs_readdata_25_port, avs_readdata_24_port, 
      avs_readdata_23_port, avs_readdata_22_port, avs_readdata_21_port, 
      avs_readdata_20_port, avs_readdata_19_port, avs_readdata_18_port, 
      avs_readdata_17_port, avs_readdata_16_port, avs_readdata_15_port, 
      avs_readdata_14_port, avs_readdata_13_port, avs_readdata_12_port, 
      avs_readdata_11_port, avs_readdata_10_port, avs_readdata_9_port, 
      avs_readdata_8_port, avs_readdata_7_port, avs_readdata_6_port, 
      avs_readdata_5_port, avs_readdata_4_port, avs_readdata_3_port, 
      avs_readdata_2_port, avs_readdata_1_port, avs_readdata_0_port, 
      stop_sim_port, out_buf_255_port, out_buf_254_port, out_buf_253_port, 
      out_buf_252_port, out_buf_251_port, out_buf_250_port, out_buf_249_port, 
      out_buf_248_port, out_buf_247_port, out_buf_246_port, out_buf_245_port, 
      out_buf_244_port, out_buf_243_port, out_buf_242_port, out_buf_241_port, 
      out_buf_240_port, out_buf_239_port, out_buf_238_port, out_buf_237_port, 
      out_buf_236_port, out_buf_235_port, out_buf_234_port, out_buf_233_port, 
      out_buf_232_port, out_buf_231_port, out_buf_230_port, out_buf_229_port, 
      out_buf_228_port, out_buf_227_port, out_buf_226_port, out_buf_225_port, 
      out_buf_224_port, out_buf_223_port, out_buf_222_port, out_buf_221_port, 
      out_buf_220_port, out_buf_219_port, out_buf_218_port, out_buf_217_port, 
      out_buf_216_port, out_buf_215_port, out_buf_214_port, out_buf_213_port, 
      out_buf_212_port, out_buf_211_port, out_buf_210_port, out_buf_209_port, 
      out_buf_208_port, out_buf_207_port, out_buf_206_port, out_buf_205_port, 
      out_buf_204_port, out_buf_203_port, out_buf_202_port, out_buf_201_port, 
      out_buf_200_port, out_buf_199_port, out_buf_198_port, out_buf_197_port, 
      out_buf_196_port, out_buf_195_port, out_buf_194_port, out_buf_193_port, 
      out_buf_192_port, out_buf_191_port, out_buf_190_port, out_buf_189_port, 
      out_buf_188_port, out_buf_187_port, out_buf_186_port, out_buf_185_port, 
      out_buf_184_port, out_buf_183_port, out_buf_182_port, out_buf_181_port, 
      out_buf_180_port, out_buf_179_port, out_buf_178_port, out_buf_177_port, 
      out_buf_176_port, out_buf_175_port, out_buf_174_port, out_buf_173_port, 
      out_buf_172_port, out_buf_171_port, out_buf_170_port, out_buf_169_port, 
      out_buf_168_port, out_buf_167_port, out_buf_166_port, out_buf_165_port, 
      out_buf_164_port, out_buf_163_port, out_buf_162_port, out_buf_161_port, 
      out_buf_160_port, out_buf_159_port, out_buf_158_port, out_buf_157_port, 
      out_buf_156_port, out_buf_155_port, out_buf_154_port, out_buf_153_port, 
      out_buf_152_port, out_buf_151_port, out_buf_150_port, out_buf_149_port, 
      out_buf_148_port, out_buf_147_port, out_buf_146_port, out_buf_145_port, 
      out_buf_144_port, out_buf_143_port, out_buf_142_port, out_buf_141_port, 
      out_buf_140_port, out_buf_139_port, out_buf_138_port, out_buf_137_port, 
      out_buf_136_port, out_buf_135_port, out_buf_134_port, out_buf_133_port, 
      out_buf_132_port, out_buf_131_port, out_buf_130_port, out_buf_129_port, 
      out_buf_128_port, out_buf_127_port, out_buf_126_port, out_buf_125_port, 
      out_buf_124_port, out_buf_123_port, out_buf_122_port, out_buf_121_port, 
      out_buf_120_port, out_buf_119_port, out_buf_118_port, out_buf_117_port, 
      out_buf_116_port, out_buf_115_port, out_buf_114_port, out_buf_113_port, 
      out_buf_112_port, out_buf_111_port, out_buf_110_port, out_buf_109_port, 
      out_buf_108_port, out_buf_107_port, out_buf_106_port, out_buf_105_port, 
      out_buf_104_port, out_buf_103_port, out_buf_102_port, out_buf_101_port, 
      out_buf_100_port, out_buf_99_port, out_buf_98_port, out_buf_97_port, 
      out_buf_96_port, out_buf_95_port, out_buf_94_port, out_buf_93_port, 
      out_buf_92_port, out_buf_91_port, out_buf_90_port, out_buf_89_port, 
      out_buf_88_port, out_buf_87_port, out_buf_86_port, out_buf_85_port, 
      out_buf_84_port, out_buf_83_port, out_buf_82_port, out_buf_81_port, 
      out_buf_80_port, out_buf_79_port, out_buf_78_port, out_buf_77_port, 
      out_buf_76_port, out_buf_75_port, out_buf_74_port, out_buf_73_port, 
      out_buf_72_port, out_buf_71_port, out_buf_70_port, out_buf_69_port, 
      out_buf_68_port, out_buf_67_port, out_buf_66_port, out_buf_65_port, 
      out_buf_64_port, out_buf_63_port, out_buf_62_port, out_buf_61_port, 
      out_buf_60_port, out_buf_59_port, out_buf_58_port, out_buf_57_port, 
      out_buf_56_port, out_buf_55_port, out_buf_54_port, out_buf_53_port, 
      out_buf_52_port, out_buf_51_port, out_buf_50_port, out_buf_49_port, 
      out_buf_48_port, out_buf_47_port, out_buf_46_port, out_buf_45_port, 
      out_buf_44_port, out_buf_43_port, out_buf_42_port, out_buf_41_port, 
      out_buf_40_port, out_buf_39_port, out_buf_38_port, out_buf_37_port, 
      out_buf_36_port, out_buf_35_port, out_buf_34_port, out_buf_33_port, 
      out_buf_32_port, out_buf_31_port, out_buf_30_port, out_buf_29_port, 
      out_buf_28_port, out_buf_27_port, out_buf_26_port, out_buf_25_port, 
      out_buf_24_port, out_buf_23_port, out_buf_22_port, out_buf_21_port, 
      out_buf_20_port, out_buf_19_port, out_buf_18_port, out_buf_17_port, 
      out_buf_16_port, out_buf_15_port, out_buf_14_port, out_buf_13_port, 
      out_buf_12_port, out_buf_11_port, out_buf_10_port, out_buf_9_port, 
      out_buf_8_port, out_buf_7_port, out_buf_6_port, out_buf_5_port, 
      out_buf_4_port, out_buf_3_port, out_buf_2_port, out_buf_1_port, 
      out_buf_0_port, coeff_memory_0_31_port, coeff_memory_0_30_port, 
      coeff_memory_0_29_port, coeff_memory_0_28_port, coeff_memory_0_27_port, 
      coeff_memory_0_26_port, coeff_memory_0_25_port, coeff_memory_0_24_port, 
      coeff_memory_0_23_port, coeff_memory_0_22_port, coeff_memory_0_21_port, 
      coeff_memory_0_20_port, coeff_memory_0_19_port, coeff_memory_0_18_port, 
      coeff_memory_0_17_port, coeff_memory_0_16_port, coeff_memory_0_15_port, 
      coeff_memory_0_14_port, coeff_memory_0_13_port, coeff_memory_0_12_port, 
      coeff_memory_0_11_port, coeff_memory_0_10_port, coeff_memory_0_9_port, 
      coeff_memory_0_8_port, coeff_memory_0_7_port, coeff_memory_0_6_port, 
      coeff_memory_0_5_port, coeff_memory_0_4_port, coeff_memory_0_3_port, 
      coeff_memory_0_2_port, coeff_memory_0_1_port, coeff_memory_0_0_port, 
      coeff_memory_1_31_port, coeff_memory_1_30_port, coeff_memory_1_29_port, 
      coeff_memory_1_28_port, coeff_memory_1_27_port, coeff_memory_1_26_port, 
      coeff_memory_1_25_port, coeff_memory_1_24_port, coeff_memory_1_23_port, 
      coeff_memory_1_22_port, coeff_memory_1_21_port, coeff_memory_1_20_port, 
      coeff_memory_1_19_port, coeff_memory_1_18_port, coeff_memory_1_17_port, 
      coeff_memory_1_16_port, coeff_memory_1_15_port, coeff_memory_1_14_port, 
      coeff_memory_1_13_port, coeff_memory_1_12_port, coeff_memory_1_11_port, 
      coeff_memory_1_10_port, coeff_memory_1_9_port, coeff_memory_1_8_port, 
      coeff_memory_1_7_port, coeff_memory_1_6_port, coeff_memory_1_5_port, 
      coeff_memory_1_4_port, coeff_memory_1_3_port, coeff_memory_1_2_port, 
      coeff_memory_1_1_port, coeff_memory_1_0_port, coeff_memory_2_31_port, 
      coeff_memory_2_30_port, coeff_memory_2_29_port, coeff_memory_2_28_port, 
      coeff_memory_2_27_port, coeff_memory_2_26_port, coeff_memory_2_25_port, 
      coeff_memory_2_24_port, coeff_memory_2_23_port, coeff_memory_2_22_port, 
      coeff_memory_2_21_port, coeff_memory_2_20_port, coeff_memory_2_19_port, 
      coeff_memory_2_18_port, coeff_memory_2_17_port, coeff_memory_2_16_port, 
      coeff_memory_2_15_port, coeff_memory_2_14_port, coeff_memory_2_13_port, 
      coeff_memory_2_12_port, coeff_memory_2_11_port, coeff_memory_2_10_port, 
      coeff_memory_2_9_port, coeff_memory_2_8_port, coeff_memory_2_7_port, 
      coeff_memory_2_6_port, coeff_memory_2_5_port, coeff_memory_2_4_port, 
      coeff_memory_2_3_port, coeff_memory_2_2_port, coeff_memory_2_1_port, 
      coeff_memory_2_0_port, coeff_memory_3_31_port, coeff_memory_3_30_port, 
      coeff_memory_3_29_port, coeff_memory_3_28_port, coeff_memory_3_27_port, 
      coeff_memory_3_26_port, coeff_memory_3_25_port, coeff_memory_3_24_port, 
      coeff_memory_3_23_port, coeff_memory_3_22_port, coeff_memory_3_21_port, 
      coeff_memory_3_20_port, coeff_memory_3_19_port, coeff_memory_3_18_port, 
      coeff_memory_3_17_port, coeff_memory_3_16_port, coeff_memory_3_15_port, 
      coeff_memory_3_14_port, coeff_memory_3_13_port, coeff_memory_3_12_port, 
      coeff_memory_3_11_port, coeff_memory_3_10_port, coeff_memory_3_9_port, 
      coeff_memory_3_8_port, coeff_memory_3_7_port, coeff_memory_3_6_port, 
      coeff_memory_3_5_port, coeff_memory_3_4_port, coeff_memory_3_3_port, 
      coeff_memory_3_2_port, coeff_memory_3_1_port, coeff_memory_3_0_port, 
      coeff_memory_4_31_port, coeff_memory_4_30_port, coeff_memory_4_29_port, 
      coeff_memory_4_28_port, coeff_memory_4_27_port, coeff_memory_4_26_port, 
      coeff_memory_4_25_port, coeff_memory_4_24_port, coeff_memory_4_23_port, 
      coeff_memory_4_22_port, coeff_memory_4_21_port, coeff_memory_4_20_port, 
      coeff_memory_4_19_port, coeff_memory_4_18_port, coeff_memory_4_17_port, 
      coeff_memory_4_16_port, coeff_memory_4_15_port, coeff_memory_4_14_port, 
      coeff_memory_4_13_port, coeff_memory_4_12_port, coeff_memory_4_11_port, 
      coeff_memory_4_10_port, coeff_memory_4_9_port, coeff_memory_4_8_port, 
      coeff_memory_4_7_port, coeff_memory_4_6_port, coeff_memory_4_5_port, 
      coeff_memory_4_4_port, coeff_memory_4_3_port, coeff_memory_4_2_port, 
      coeff_memory_4_1_port, coeff_memory_4_0_port, operand_regs_255_port, 
      operand_regs_254_port, operand_regs_253_port, operand_regs_252_port, 
      operand_regs_251_port, operand_regs_250_port, operand_regs_249_port, 
      operand_regs_248_port, operand_regs_247_port, operand_regs_246_port, 
      operand_regs_245_port, operand_regs_244_port, operand_regs_243_port, 
      operand_regs_242_port, operand_regs_241_port, operand_regs_240_port, 
      operand_regs_239_port, operand_regs_238_port, operand_regs_237_port, 
      operand_regs_236_port, operand_regs_235_port, operand_regs_234_port, 
      operand_regs_233_port, operand_regs_232_port, operand_regs_231_port, 
      operand_regs_230_port, operand_regs_229_port, operand_regs_228_port, 
      operand_regs_227_port, operand_regs_226_port, operand_regs_225_port, 
      operand_regs_224_port, operand_regs_223_port, operand_regs_222_port, 
      operand_regs_221_port, operand_regs_220_port, operand_regs_219_port, 
      operand_regs_218_port, operand_regs_217_port, operand_regs_216_port, 
      operand_regs_215_port, operand_regs_214_port, operand_regs_213_port, 
      operand_regs_212_port, operand_regs_211_port, operand_regs_210_port, 
      operand_regs_209_port, operand_regs_208_port, operand_regs_207_port, 
      operand_regs_206_port, operand_regs_205_port, operand_regs_204_port, 
      operand_regs_203_port, operand_regs_202_port, operand_regs_201_port, 
      operand_regs_200_port, operand_regs_199_port, operand_regs_198_port, 
      operand_regs_197_port, operand_regs_196_port, operand_regs_195_port, 
      operand_regs_194_port, operand_regs_193_port, operand_regs_192_port, 
      operand_regs_191_port, operand_regs_190_port, operand_regs_189_port, 
      operand_regs_188_port, operand_regs_187_port, operand_regs_186_port, 
      operand_regs_185_port, operand_regs_184_port, operand_regs_183_port, 
      operand_regs_182_port, operand_regs_181_port, operand_regs_180_port, 
      operand_regs_179_port, operand_regs_178_port, operand_regs_177_port, 
      operand_regs_176_port, operand_regs_175_port, operand_regs_174_port, 
      operand_regs_173_port, operand_regs_172_port, operand_regs_171_port, 
      operand_regs_170_port, operand_regs_169_port, operand_regs_168_port, 
      operand_regs_167_port, operand_regs_166_port, operand_regs_165_port, 
      operand_regs_164_port, operand_regs_163_port, operand_regs_162_port, 
      operand_regs_161_port, operand_regs_160_port, operand_regs_159_port, 
      operand_regs_158_port, operand_regs_157_port, operand_regs_156_port, 
      operand_regs_155_port, operand_regs_154_port, operand_regs_153_port, 
      operand_regs_152_port, operand_regs_151_port, operand_regs_150_port, 
      operand_regs_149_port, operand_regs_148_port, operand_regs_147_port, 
      operand_regs_146_port, operand_regs_145_port, operand_regs_144_port, 
      operand_regs_143_port, operand_regs_142_port, operand_regs_141_port, 
      operand_regs_140_port, operand_regs_139_port, operand_regs_138_port, 
      operand_regs_137_port, operand_regs_136_port, operand_regs_135_port, 
      operand_regs_134_port, operand_regs_133_port, operand_regs_132_port, 
      operand_regs_131_port, operand_regs_130_port, operand_regs_129_port, 
      operand_regs_128_port, operand_regs_127_port, operand_regs_126_port, 
      operand_regs_125_port, operand_regs_124_port, operand_regs_123_port, 
      operand_regs_122_port, operand_regs_121_port, operand_regs_120_port, 
      operand_regs_119_port, operand_regs_118_port, operand_regs_117_port, 
      operand_regs_116_port, operand_regs_115_port, operand_regs_114_port, 
      operand_regs_113_port, operand_regs_112_port, operand_regs_111_port, 
      operand_regs_110_port, operand_regs_109_port, operand_regs_108_port, 
      operand_regs_107_port, operand_regs_106_port, operand_regs_105_port, 
      operand_regs_104_port, operand_regs_103_port, operand_regs_102_port, 
      operand_regs_101_port, operand_regs_100_port, operand_regs_99_port, 
      operand_regs_98_port, operand_regs_97_port, operand_regs_96_port, 
      operand_regs_95_port, operand_regs_94_port, operand_regs_93_port, 
      operand_regs_92_port, operand_regs_91_port, operand_regs_90_port, 
      operand_regs_89_port, operand_regs_88_port, operand_regs_87_port, 
      operand_regs_86_port, operand_regs_85_port, operand_regs_84_port, 
      operand_regs_83_port, operand_regs_82_port, operand_regs_81_port, 
      operand_regs_80_port, operand_regs_79_port, operand_regs_78_port, 
      operand_regs_77_port, operand_regs_76_port, operand_regs_75_port, 
      operand_regs_74_port, operand_regs_73_port, operand_regs_72_port, 
      operand_regs_71_port, operand_regs_70_port, operand_regs_69_port, 
      operand_regs_68_port, operand_regs_67_port, operand_regs_66_port, 
      operand_regs_65_port, operand_regs_64_port, operand_regs_63_port, 
      operand_regs_62_port, operand_regs_61_port, operand_regs_60_port, 
      operand_regs_59_port, operand_regs_58_port, operand_regs_57_port, 
      operand_regs_56_port, operand_regs_55_port, operand_regs_54_port, 
      operand_regs_53_port, operand_regs_52_port, operand_regs_51_port, 
      operand_regs_50_port, operand_regs_49_port, operand_regs_48_port, 
      operand_regs_47_port, operand_regs_46_port, operand_regs_45_port, 
      operand_regs_44_port, operand_regs_43_port, operand_regs_42_port, 
      operand_regs_41_port, operand_regs_40_port, operand_regs_39_port, 
      operand_regs_38_port, operand_regs_37_port, operand_regs_36_port, 
      operand_regs_35_port, operand_regs_34_port, operand_regs_33_port, 
      operand_regs_32_port, operand_regs_31_port, operand_regs_30_port, 
      operand_regs_29_port, operand_regs_28_port, operand_regs_27_port, 
      operand_regs_26_port, operand_regs_25_port, operand_regs_24_port, 
      operand_regs_23_port, operand_regs_22_port, operand_regs_21_port, 
      operand_regs_20_port, operand_regs_19_port, operand_regs_18_port, 
      operand_regs_17_port, operand_regs_16_port, operand_regs_15_port, 
      operand_regs_14_port, operand_regs_13_port, operand_regs_12_port, 
      operand_regs_11_port, operand_regs_10_port, operand_regs_9_port, 
      operand_regs_8_port, operand_regs_7_port, operand_regs_6_port, 
      operand_regs_5_port, operand_regs_4_port, operand_regs_3_port, 
      operand_regs_2_port, operand_regs_1_port, operand_regs_0_port, in_trigger
      , out_trigger, coeff_load, operand_load, read_comp_res, filt_mult_inputs,
      N66, comp_res_159_port, comp_res_158_port, comp_res_157_port, 
      comp_res_156_port, comp_res_155_port, comp_res_154_port, 
      comp_res_153_port, comp_res_152_port, comp_res_151_port, 
      comp_res_150_port, comp_res_149_port, comp_res_148_port, 
      comp_res_147_port, comp_res_146_port, comp_res_145_port, 
      comp_res_144_port, comp_res_143_port, comp_res_142_port, 
      comp_res_141_port, comp_res_140_port, comp_res_139_port, 
      comp_res_138_port, comp_res_137_port, comp_res_136_port, 
      comp_res_135_port, comp_res_134_port, comp_res_133_port, 
      comp_res_132_port, comp_res_131_port, comp_res_130_port, 
      comp_res_129_port, comp_res_128_port, comp_res_127_port, 
      comp_res_126_port, comp_res_125_port, comp_res_124_port, 
      comp_res_123_port, comp_res_122_port, comp_res_121_port, 
      comp_res_120_port, comp_res_119_port, comp_res_118_port, 
      comp_res_117_port, comp_res_116_port, comp_res_115_port, 
      comp_res_114_port, comp_res_113_port, comp_res_112_port, 
      comp_res_111_port, comp_res_110_port, comp_res_109_port, 
      comp_res_108_port, comp_res_107_port, comp_res_106_port, 
      comp_res_105_port, comp_res_104_port, comp_res_103_port, 
      comp_res_102_port, comp_res_101_port, comp_res_100_port, comp_res_99_port
      , comp_res_98_port, comp_res_97_port, comp_res_96_port, comp_res_95_port,
      comp_res_94_port, comp_res_93_port, comp_res_92_port, comp_res_91_port, 
      comp_res_90_port, comp_res_89_port, comp_res_88_port, comp_res_87_port, 
      comp_res_86_port, comp_res_85_port, comp_res_84_port, comp_res_83_port, 
      comp_res_82_port, comp_res_81_port, comp_res_80_port, comp_res_79_port, 
      comp_res_78_port, comp_res_77_port, comp_res_76_port, comp_res_75_port, 
      comp_res_74_port, comp_res_73_port, comp_res_72_port, comp_res_71_port, 
      comp_res_70_port, comp_res_69_port, comp_res_68_port, comp_res_67_port, 
      comp_res_66_port, comp_res_65_port, comp_res_64_port, comp_res_63_port, 
      comp_res_62_port, comp_res_61_port, comp_res_60_port, comp_res_59_port, 
      comp_res_58_port, comp_res_57_port, comp_res_56_port, comp_res_55_port, 
      comp_res_54_port, comp_res_53_port, comp_res_52_port, comp_res_51_port, 
      comp_res_50_port, comp_res_49_port, comp_res_48_port, comp_res_47_port, 
      comp_res_46_port, comp_res_45_port, comp_res_44_port, comp_res_43_port, 
      comp_res_42_port, comp_res_41_port, comp_res_40_port, comp_res_39_port, 
      comp_res_38_port, comp_res_37_port, comp_res_36_port, comp_res_35_port, 
      comp_res_34_port, comp_res_33_port, comp_res_32_port, comp_res_31_port, 
      comp_res_30_port, comp_res_29_port, comp_res_28_port, comp_res_27_port, 
      comp_res_26_port, comp_res_25_port, comp_res_24_port, comp_res_23_port, 
      comp_res_22_port, comp_res_21_port, comp_res_20_port, comp_res_19_port, 
      comp_res_18_port, comp_res_17_port, comp_res_16_port, comp_res_15_port, 
      comp_res_14_port, comp_res_13_port, comp_res_12_port, comp_res_11_port, 
      comp_res_10_port, comp_res_9_port, comp_res_8_port, comp_res_7_port, 
      comp_res_6_port, comp_res_5_port, comp_res_4_port, comp_res_3_port, 
      comp_res_2_port, comp_res_1_port, comp_res_0_port, N1978, N1979, N1980, 
      N1981, N1982, N1983, N1984, N1985, N1986, N1987, N1988, N1989, N1990, 
      N1991, N1992, N1993, N1994, N1995, N1996, N1997, N1998, N1999, N2000, 
      N2001, N2002, N2003, N2004, N2005, N2006, N2007, N2008, N2009, 
      in_buf_255_port, in_buf_254_port, in_buf_253_port, in_buf_252_port, 
      in_buf_251_port, in_buf_250_port, in_buf_249_port, in_buf_248_port, 
      in_buf_247_port, in_buf_246_port, in_buf_245_port, in_buf_244_port, 
      in_buf_243_port, in_buf_242_port, in_buf_241_port, in_buf_240_port, 
      in_buf_239_port, in_buf_238_port, in_buf_237_port, in_buf_236_port, 
      in_buf_235_port, in_buf_234_port, in_buf_233_port, in_buf_232_port, 
      in_buf_231_port, in_buf_230_port, in_buf_229_port, in_buf_228_port, 
      in_buf_227_port, in_buf_226_port, in_buf_225_port, in_buf_224_port, 
      in_buf_223_port, in_buf_222_port, in_buf_221_port, in_buf_220_port, 
      in_buf_219_port, in_buf_218_port, in_buf_217_port, in_buf_216_port, 
      in_buf_215_port, in_buf_214_port, in_buf_213_port, in_buf_212_port, 
      in_buf_211_port, in_buf_210_port, in_buf_209_port, in_buf_208_port, 
      in_buf_207_port, in_buf_206_port, in_buf_205_port, in_buf_204_port, 
      in_buf_203_port, in_buf_202_port, in_buf_201_port, in_buf_200_port, 
      in_buf_199_port, in_buf_198_port, in_buf_197_port, in_buf_196_port, 
      in_buf_195_port, in_buf_194_port, in_buf_193_port, in_buf_192_port, 
      in_buf_191_port, in_buf_190_port, in_buf_189_port, in_buf_188_port, 
      in_buf_187_port, in_buf_186_port, in_buf_185_port, in_buf_184_port, 
      in_buf_183_port, in_buf_182_port, in_buf_181_port, in_buf_180_port, 
      in_buf_179_port, in_buf_178_port, in_buf_177_port, in_buf_176_port, 
      in_buf_175_port, in_buf_174_port, in_buf_173_port, in_buf_172_port, 
      in_buf_171_port, in_buf_170_port, in_buf_169_port, in_buf_168_port, 
      in_buf_167_port, in_buf_166_port, in_buf_165_port, in_buf_164_port, 
      in_buf_163_port, in_buf_162_port, in_buf_161_port, in_buf_160_port, 
      in_buf_159_port, in_buf_158_port, in_buf_157_port, in_buf_156_port, 
      in_buf_155_port, in_buf_154_port, in_buf_153_port, in_buf_152_port, 
      in_buf_151_port, in_buf_150_port, in_buf_149_port, in_buf_148_port, 
      in_buf_147_port, in_buf_146_port, in_buf_145_port, in_buf_144_port, 
      in_buf_143_port, in_buf_142_port, in_buf_141_port, in_buf_140_port, 
      in_buf_139_port, in_buf_138_port, in_buf_137_port, in_buf_136_port, 
      in_buf_135_port, in_buf_134_port, in_buf_133_port, in_buf_132_port, 
      in_buf_131_port, in_buf_130_port, in_buf_129_port, in_buf_128_port, 
      in_buf_127_port, in_buf_126_port, in_buf_125_port, in_buf_124_port, 
      in_buf_123_port, in_buf_122_port, in_buf_121_port, in_buf_120_port, 
      in_buf_119_port, in_buf_118_port, in_buf_117_port, in_buf_116_port, 
      in_buf_115_port, in_buf_114_port, in_buf_113_port, in_buf_112_port, 
      in_buf_111_port, in_buf_110_port, in_buf_109_port, in_buf_108_port, 
      in_buf_107_port, in_buf_106_port, in_buf_105_port, in_buf_104_port, 
      in_buf_103_port, in_buf_102_port, in_buf_101_port, in_buf_100_port, 
      in_buf_99_port, in_buf_98_port, in_buf_97_port, in_buf_96_port, 
      in_buf_95_port, in_buf_94_port, in_buf_93_port, in_buf_92_port, 
      in_buf_91_port, in_buf_90_port, in_buf_89_port, in_buf_88_port, 
      in_buf_87_port, in_buf_86_port, in_buf_85_port, in_buf_84_port, 
      in_buf_83_port, in_buf_82_port, in_buf_81_port, in_buf_80_port, 
      in_buf_79_port, in_buf_78_port, in_buf_77_port, in_buf_76_port, 
      in_buf_75_port, in_buf_74_port, in_buf_73_port, in_buf_72_port, 
      in_buf_71_port, in_buf_70_port, in_buf_69_port, in_buf_68_port, 
      in_buf_67_port, in_buf_66_port, in_buf_65_port, in_buf_64_port, 
      in_buf_63_port, in_buf_62_port, in_buf_61_port, in_buf_60_port, 
      in_buf_59_port, in_buf_58_port, in_buf_57_port, in_buf_56_port, 
      in_buf_55_port, in_buf_54_port, in_buf_53_port, in_buf_52_port, 
      in_buf_51_port, in_buf_50_port, in_buf_49_port, in_buf_48_port, 
      in_buf_47_port, in_buf_46_port, in_buf_45_port, in_buf_44_port, 
      in_buf_43_port, in_buf_42_port, in_buf_41_port, in_buf_40_port, 
      in_buf_39_port, in_buf_38_port, in_buf_37_port, in_buf_36_port, 
      in_buf_35_port, in_buf_34_port, in_buf_33_port, in_buf_32_port, 
      in_buf_31_port, in_buf_30_port, in_buf_29_port, in_buf_28_port, 
      in_buf_27_port, in_buf_26_port, in_buf_25_port, in_buf_24_port, 
      in_buf_23_port, in_buf_22_port, in_buf_21_port, in_buf_20_port, 
      in_buf_19_port, in_buf_18_port, in_buf_17_port, in_buf_16_port, 
      in_buf_15_port, in_buf_14_port, in_buf_13_port, in_buf_12_port, 
      in_buf_11_port, in_buf_10_port, in_buf_9_port, in_buf_8_port, 
      in_buf_7_port, in_buf_6_port, in_buf_5_port, in_buf_4_port, in_buf_3_port
      , in_buf_2_port, in_buf_1_port, in_buf_0_port, N2010, N2011, N2012, N2013
      , N2014, N2015, N2016, N2017, N2018, N2019, N2020, N2021, N2022, N2023, 
      N2024, N2025, N2026, N2027, N2028, N2029, N2030, N2031, N2032, N2033, 
      N2034, N2035, N2036, N2037, N2038, N2039, N2040, N2041, in_busy, out_busy
      , in_counter_2_port, in_counter_1_port, in_counter_0_port, odd, odd1, 
      N2850, N2851, N2852, N2853, N2854, N2855, N2856, N2857, N2858, N2859, 
      N2860, N2861, N2862, N2863, N2864, N2865, N2867, N2868, N2869, N2870, 
      N2871, N2872, N2873, N2874, N2875, N2876, N2877, N2878, N2879, N2880, 
      N2881, N2882, N2888, N2889, N2890, N2891, N2892, N2893, N2894, N2895, 
      N2896, N2897, N2898, N2899, N2900, N2901, N2902, N2903, N2913, N2914, 
      N2915, N2916, N2917, N2918, N2919, N2920, N2921, N2922, N2923, N2924, 
      N2925, N2926, N2927, N2928, N2929, N2930, N2931, N2932, N2933, N2934, 
      N2935, N2936, N2937, N2938, N2939, N2940, N2941, N2942, N2943, N2944, 
      N2945, N2946, N2947, N2948, N2949, N2950, N2951, N2952, N2953, N2954, 
      N2955, N2956, N2957, N2958, N2959, N2960, N2961, N2962, N2963, N2964, 
      N2965, N2966, N2967, N2968, N2969, N2970, N2971, N2972, N2973, N2974, 
      N2975, N2976, N2977, N2978, N2979, N2980, N2981, N2982, N2983, N2984, 
      N2985, N2986, N2987, N2988, N2989, N2990, N2991, N2992, N2993, N2994, 
      N2995, N2996, N2997, N2998, N2999, N3000, N3001, N3002, N3003, N3004, 
      N3005, N3006, N3007, N3008, N3009, N3010, N3011, N3012, N3013, N3014, 
      N3015, N3016, N3017, N3018, N3019, N3020, N3021, N3022, N3023, N3024, 
      N3025, N3026, N3027, N3028, N3029, N3030, N3031, N3032, N3033, N3034, 
      N3035, N3036, N3037, N3038, N3039, N3040, N3041, N3042, N3043, N3044, 
      N3045, N3046, N3047, N3048, N3049, N3050, N3051, N3052, N3053, N3054, 
      N3055, N3056, N3057, N3058, N3059, N3060, N3061, N3062, N3063, N3064, 
      N3065, N3066, N3067, N3068, N3069, N3070, N3071, N3072, N3073, N3074, 
      N3075, N3076, N3077, N3078, N3079, N3080, N3081, N3082, N3083, N3084, 
      N3085, N3086, N3087, N3088, N3089, N3090, N3091, N3092, N3093, N3094, 
      N3095, N3096, N3097, N3098, N3099, N3100, N3101, N3102, N3103, N3104, 
      N3105, N3106, N3107, N3108, N3109, N3110, N3111, N3112, N3113, N3114, 
      N3115, N3116, N3117, N3118, N3119, N3120, N3121, N3122, N3123, N3124, 
      N3125, N3126, N3127, N3128, N3129, N3130, N3131, N3132, N3133, N3134, 
      N3135, N3136, N3137, N3138, N3139, N3140, N3141, N3142, N3143, N3144, 
      N3145, N3146, N3147, N3148, N3149, N3150, N3151, N3152, N3153, N3154, 
      N3155, N3156, N3157, N3158, N3159, N3160, N3161, N3162, N3163, N3164, 
      N3165, N3166, N3167, N3168, N3233, N3234, N3235, N3236, N3237, N3238, 
      N3239, N3240, N3241, N3242, N3243, N3244, N3245, N3246, N3247, N3248, 
      N3249, N3250, N3251, N3252, N3253, N3254, N3255, N3256, N3257, N3258, 
      N3259, N3260, N3261, N3262, N3263, N3264, N3265, N3266, N3267, N3268, 
      N3269, N3270, N3271, N3272, N3273, N3274, N3275, N3276, N3277, N3278, 
      N3279, N3280, N3281, N3282, N3283, N3284, N3285, N3286, N3287, N3288, 
      N3289, N3290, N3291, N3292, N3293, N3294, N3295, N3296, N3297, N3298, 
      N3299, N3300, N3301, N3302, N3303, N3304, N3305, N3306, N3307, N3308, 
      N3309, N3310, N3311, N3312, N3313, N3314, N3315, N3316, N3317, N3318, 
      N3319, N3320, N3321, N3322, N3323, N3324, N3325, N3326, N3327, N3328, 
      N3329, N3330, N3331, N3332, N3333, N3334, N3335, N3336, N3337, N3338, 
      N3339, N3340, N3341, N3342, N3343, N3344, N3345, N3346, N3347, N3348, 
      N3349, N3350, N3351, N3352, N3353, N3354, N3355, N3356, N3357, N3358, 
      N3359, N3360, N3361, N3362, N3363, N3364, N3365, N3366, N3367, N3368, 
      N3369, N3370, N3371, N3372, N3373, N3374, N3375, N3376, N3377, N3378, 
      N3379, N3380, N3381, N3382, N3383, N3384, N3385, N3386, N3387, N3388, 
      N3389, N3390, N3391, N3392, n4, n5, n10, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, 
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n5900, n6000,
      n6100, n6300, n6400, n65, n70, n72, n73, n74, n76, n77, n78, n79, n81, 
      n84, n85, n86, n87, n88, n89, n91, n92, n95, n96, n100, n101, n104, n110,
      n111, n114, n115, n118, n119, n120, n154, n155, n156, n157, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, 
      n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, 
      n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, 
      n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, 
      n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, 
      n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, 
      n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, 
      n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, 
      n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, 
      n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, 
      n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, 
      n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, 
      n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, 
      n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, 
      n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, 
      n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, 
      n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, 
      n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, 
      n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, 
      n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, 
      n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, 
      n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, 
      n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, 
      n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, 
      n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, 
      n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, 
      n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, 
      n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, 
      n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n5901, n591, 
      n592, n593, n594, n595, n596, n597, n598, n599, n6001, n601, n602, n603, 
      n604, n605, n606, n607, n608, n609, n6101, n611, n612, n613, n614, n615, 
      n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, 
      n628, n629, n6301, n631, n632, n633, n634, n635, n636, n637, n638, n639, 
      n6401, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, 
      n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, 
      n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, 
      n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, 
      n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, 
      n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, 
      n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, 
      n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, 
      n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, 
      n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, 
      n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, 
      n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, 
      n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, 
      n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, 
      n808, n809, n810, n811, n812, n813, n_1160, n_1161, n_1162, n_1163, 
      n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, 
      n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, 
      n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, 
      n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, 
      n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, 
      n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, 
      n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, 
      n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, 
      n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, 
      n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, 
      n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, 
      n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, 
      n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, 
      n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, 
      n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, 
      n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, 
      n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, 
      n_1317, n_1318, n_1319 : std_logic;

begin
   avs_readdata <= ( avs_readdata_31_port, avs_readdata_30_port, 
      avs_readdata_29_port, avs_readdata_28_port, avs_readdata_27_port, 
      avs_readdata_26_port, avs_readdata_25_port, avs_readdata_24_port, 
      avs_readdata_23_port, avs_readdata_22_port, avs_readdata_21_port, 
      avs_readdata_20_port, avs_readdata_19_port, avs_readdata_18_port, 
      avs_readdata_17_port, avs_readdata_16_port, avs_readdata_15_port, 
      avs_readdata_14_port, avs_readdata_13_port, avs_readdata_12_port, 
      avs_readdata_11_port, avs_readdata_10_port, avs_readdata_9_port, 
      avs_readdata_8_port, avs_readdata_7_port, avs_readdata_6_port, 
      avs_readdata_5_port, avs_readdata_4_port, avs_readdata_3_port, 
      avs_readdata_2_port, avs_readdata_1_port, avs_readdata_0_port );
   clk_out <= clk;
   stop_sim <= stop_sim_port;
   
   U3 : OAI22D1 port map( A1 => N63, A2 => n4, B1 => n5, B2 => n813, Z => n201)
                           ;
   U4 : AOI21D1 port map( A1 => out_busy, A2 => n810, B => n801, Z => n5);
   U7 : AOI22D1 port map( A1 => N1978, A2 => n268, B1 => N2010, B2 => n698, Z 
                           => n10);
   U9 : AOI22D1 port map( A1 => N2011, A2 => n12, B1 => avs_readdata_30_port, 
                           B2 => n700, Z => n15);
   U12 : AOI22D1 port map( A1 => N1980, A2 => n268, B1 => N2012, B2 => n698, Z 
                           => n16);
   U14 : AOI22D1 port map( A1 => N2013, A2 => n698, B1 => avs_readdata_28_port,
                           B2 => n700, Z => n18);
   U17 : AOI22D1 port map( A1 => N1982, A2 => n268, B1 => N2014, B2 => n698, Z 
                           => n19);
   U19 : AOI22D1 port map( A1 => N2015, A2 => n698, B1 => avs_readdata_26_port,
                           B2 => n700, Z => n21);
   U22 : AOI22D1 port map( A1 => N1984, A2 => n268, B1 => N2016, B2 => n698, Z 
                           => n22);
   U24 : AOI22D1 port map( A1 => N2017, A2 => n698, B1 => avs_readdata_24_port,
                           B2 => n700, Z => n24);
   U27 : AOI22D1 port map( A1 => N1986, A2 => n268, B1 => N2018, B2 => n698, Z 
                           => n25);
   U29 : AOI22D1 port map( A1 => N2019, A2 => n12, B1 => avs_readdata_22_port, 
                           B2 => n700, Z => n27);
   U32 : AOI22D1 port map( A1 => N1988, A2 => n268, B1 => N2020, B2 => n698, Z 
                           => n28);
   U34 : AOI22D1 port map( A1 => N2021, A2 => n12, B1 => avs_readdata_20_port, 
                           B2 => n700, Z => n30);
   U37 : AOI22D1 port map( A1 => N1990, A2 => n268, B1 => N2022, B2 => n698, Z 
                           => n31);
   U39 : AOI22D1 port map( A1 => N2023, A2 => n12, B1 => avs_readdata_18_port, 
                           B2 => n700, Z => n33);
   U42 : AOI22D1 port map( A1 => N1992, A2 => n268, B1 => N2024, B2 => n698, Z 
                           => n34);
   U44 : AOI22D1 port map( A1 => N2025, A2 => n12, B1 => avs_readdata_16_port, 
                           B2 => n700, Z => n36);
   U47 : AOI22D1 port map( A1 => N1994, A2 => n268, B1 => N2026, B2 => n698, Z 
                           => n37);
   U49 : AOI22D1 port map( A1 => N2027, A2 => n12, B1 => avs_readdata_14_port, 
                           B2 => n700, Z => n39);
   U52 : AOI22D1 port map( A1 => N1996, A2 => n268, B1 => N2028, B2 => n12, Z 
                           => n40);
   U54 : AOI22D1 port map( A1 => N2029, A2 => n12, B1 => avs_readdata_12_port, 
                           B2 => n700, Z => n42);
   U57 : AOI22D1 port map( A1 => N1998, A2 => n268, B1 => N2030, B2 => n12, Z 
                           => n43);
   U59 : AOI22D1 port map( A1 => N2031, A2 => n12, B1 => avs_readdata_10_port, 
                           B2 => n700, Z => n45);
   U62 : AOI22D1 port map( A1 => N2000, A2 => n268, B1 => N2032, B2 => n12, Z 
                           => n46);
   U64 : AOI22D1 port map( A1 => N2033, A2 => n12, B1 => avs_readdata_8_port, 
                           B2 => n700, Z => n48);
   U67 : AOI22D1 port map( A1 => N2002, A2 => n268, B1 => N2034, B2 => n698, Z 
                           => n49);
   U69 : AOI22D1 port map( A1 => N2035, A2 => n12, B1 => avs_readdata_6_port, 
                           B2 => n700, Z => n51);
   U72 : AOI22D1 port map( A1 => N2004, A2 => n268, B1 => N2036, B2 => n698, Z 
                           => n52);
   U74 : AOI22D1 port map( A1 => N2037, A2 => n12, B1 => avs_readdata_4_port, 
                           B2 => n700, Z => n54);
   U77 : AOI22D1 port map( A1 => N2006, A2 => n268, B1 => N2038, B2 => n698, Z 
                           => n55);
   U79 : AOI22D1 port map( A1 => N2039, A2 => n12, B1 => avs_readdata_2_port, 
                           B2 => n700, Z => n57);
   U82 : AOI22D1 port map( A1 => N2008, A2 => n268, B1 => N2040, B2 => n698, Z 
                           => n58);
   U84 : AOI22D1 port map( A1 => N2041, A2 => n698, B1 => avs_readdata_0_port, 
                           B2 => n700, Z => n6100);
   U94 : AOI21D1 port map( A1 => n798, A2 => in_trigger, B => n72, Z => n70);
   U95 : OAI22D1 port map( A1 => n6400, A2 => n73, B1 => n74, B2 => n802, Z => 
                           n72);
   U96 : AOI22D1 port map( A1 => in_busy, A2 => n307, B1 => out_busy, B2 => 
                           n306, Z => n73);
   U97 : EXNOR2D1 port map( A1 => n811, A2 => n76, Z => n234);
   U98 : AOI22D1 port map( A1 => n77, A2 => out_busy, B1 => n811, B2 => n802, Z
                           => n76);
   U100 : OAI22D1 port map( A1 => n813, A2 => n4, B1 => n79, B2 => n696, Z => 
                           n235);
   U103 : OAI32D1 port map( A1 => n801, A2 => N62, A3 => n811, B1 => n810, B2 
                           => n81, Z => n236);
   U105 : OAI32D1 port map( A1 => n812, A2 => n811, A3 => n78, B1 => out_busy, 
                           B2 => n802, Z => n81);
   U111 : OAI211D1 port map( A1 => n808, A2 => n84, B => n85, C => n86, Z => 
                           n237);
   U113 : OAI22D1 port map( A1 => n800, A2 => n88, B1 => n89, B2 => n809, Z => 
                           n238);
   U115 : EXNOR2D1 port map( A1 => in_busy, A2 => n161, Z => n239);
   U117 : AOI22D1 port map( A1 => avs_writedata(0), A2 => n797, B1 => 
                           out_trigger, B2 => n74, Z => n92);
   U122 : AOI22D1 port map( A1 => avs_writedata(0), A2 => n798, B1 => 
                           in_trigger, B2 => n96, Z => n95);
   U125 : EXNOR2D1 port map( A1 => n811, A2 => n697, Z => n154);
   U126 : EXNOR2D1 port map( A1 => n803, A2 => in_busy, Z => n156);
   U130 : AOI22D1 port map( A1 => odd, A2 => n91, B1 => n101, B2 => in_busy, Z 
                           => n100);
   U131 : OAI21D1 port map( A1 => in_counter_1_port, A2 => n806, B => n804, Z 
                           => n91);
   U200 : OA21M20D1 port map( A1 => n806, A2 => in_trigger, B => n176, Z => 
                           n161);
   mult_21_C241 : gp_custom_DW_mult_tc_5 port map( a(31) => N2944, a(30) => 
                           N2943, a(29) => N2942, a(28) => N2941, a(27) => 
                           N2940, a(26) => N2939, a(25) => N2938, a(24) => 
                           N2937, a(23) => N2936, a(22) => N2935, a(21) => 
                           N2934, a(20) => N2933, a(19) => N2932, a(18) => 
                           N2931, a(17) => N2930, a(16) => N2929, a(15) => 
                           N2928, a(14) => N2927, a(13) => N2926, a(12) => 
                           N2925, a(11) => N2924, a(10) => N2923, a(9) => N2922
                           , a(8) => N2921, a(7) => N2920, a(6) => N2919, a(5) 
                           => N2918, a(4) => N2917, a(3) => N2916, a(2) => 
                           N2915, a(1) => N2914, a(0) => N2913, b(31) => N3104,
                           b(30) => N3103, b(29) => N3102, b(28) => N3101, 
                           b(27) => N3100, b(26) => N3099, b(25) => N3098, 
                           b(24) => N3097, b(23) => N3096, b(22) => N3095, 
                           b(21) => N3094, b(20) => N3093, b(19) => N3092, 
                           b(18) => N3091, b(17) => N3090, b(16) => N3089, 
                           b(15) => N3088, b(14) => N3087, b(13) => N3086, 
                           b(12) => N3085, b(11) => N3084, b(10) => N3083, b(9)
                           => N3082, b(8) => N3081, b(7) => N3080, b(6) => 
                           N3079, b(5) => N3078, b(4) => N3077, b(3) => N3076, 
                           b(2) => N3075, b(1) => N3074, b(0) => N3073, 
                           product(63) => n_1160, product(62) => n_1161, 
                           product(61) => n_1162, product(60) => n_1163, 
                           product(59) => n_1164, product(58) => n_1165, 
                           product(57) => n_1166, product(56) => n_1167, 
                           product(55) => n_1168, product(54) => n_1169, 
                           product(53) => n_1170, product(52) => n_1171, 
                           product(51) => n_1172, product(50) => n_1173, 
                           product(49) => n_1174, product(48) => n_1175, 
                           product(47) => n_1176, product(46) => n_1177, 
                           product(45) => n_1178, product(44) => n_1179, 
                           product(43) => n_1180, product(42) => n_1181, 
                           product(41) => n_1182, product(40) => n_1183, 
                           product(39) => n_1184, product(38) => n_1185, 
                           product(37) => n_1186, product(36) => n_1187, 
                           product(35) => n_1188, product(34) => n_1189, 
                           product(33) => n_1190, product(32) => n_1191, 
                           product(31) => N3264, product(30) => N3263, 
                           product(29) => N3262, product(28) => N3261, 
                           product(27) => N3260, product(26) => N3259, 
                           product(25) => N3258, product(24) => N3257, 
                           product(23) => N3256, product(22) => N3255, 
                           product(21) => N3254, product(20) => N3253, 
                           product(19) => N3252, product(18) => N3251, 
                           product(17) => N3250, product(16) => N3249, 
                           product(15) => N3248, product(14) => N3247, 
                           product(13) => N3246, product(12) => N3245, 
                           product(11) => N3244, product(10) => N3243, 
                           product(9) => N3242, product(8) => N3241, product(7)
                           => N3240, product(6) => N3239, product(5) => N3238, 
                           product(4) => N3237, product(3) => N3236, product(2)
                           => N3235, product(1) => N3234, product(0) => N3233);
   mult_21_C243 : gp_custom_DW_mult_tc_6 port map( a(31) => N2976, a(30) => 
                           N2975, a(29) => N2974, a(28) => N2973, a(27) => 
                           N2972, a(26) => N2971, a(25) => N2970, a(24) => 
                           N2969, a(23) => N2968, a(22) => N2967, a(21) => 
                           N2966, a(20) => N2965, a(19) => N2964, a(18) => 
                           N2963, a(17) => N2962, a(16) => N2961, a(15) => 
                           N2960, a(14) => N2959, a(13) => N2958, a(12) => 
                           N2957, a(11) => N2956, a(10) => N2955, a(9) => N2954
                           , a(8) => N2953, a(7) => N2952, a(6) => N2951, a(5) 
                           => N2950, a(4) => N2949, a(3) => N2948, a(2) => 
                           N2947, a(1) => N2946, a(0) => N2945, b(31) => N3136,
                           b(30) => N3135, b(29) => N3134, b(28) => N3133, 
                           b(27) => N3132, b(26) => N3131, b(25) => N3130, 
                           b(24) => N3129, b(23) => N3128, b(22) => N3127, 
                           b(21) => N3126, b(20) => N3125, b(19) => N3124, 
                           b(18) => N3123, b(17) => N3122, b(16) => N3121, 
                           b(15) => N3120, b(14) => N3119, b(13) => N3118, 
                           b(12) => N3117, b(11) => N3116, b(10) => N3115, b(9)
                           => N3114, b(8) => N3113, b(7) => N3112, b(6) => 
                           N3111, b(5) => N3110, b(4) => N3109, b(3) => N3108, 
                           b(2) => N3107, b(1) => N3106, b(0) => N3105, 
                           product(63) => n_1192, product(62) => n_1193, 
                           product(61) => n_1194, product(60) => n_1195, 
                           product(59) => n_1196, product(58) => n_1197, 
                           product(57) => n_1198, product(56) => n_1199, 
                           product(55) => n_1200, product(54) => n_1201, 
                           product(53) => n_1202, product(52) => n_1203, 
                           product(51) => n_1204, product(50) => n_1205, 
                           product(49) => n_1206, product(48) => n_1207, 
                           product(47) => n_1208, product(46) => n_1209, 
                           product(45) => n_1210, product(44) => n_1211, 
                           product(43) => n_1212, product(42) => n_1213, 
                           product(41) => n_1214, product(40) => n_1215, 
                           product(39) => n_1216, product(38) => n_1217, 
                           product(37) => n_1218, product(36) => n_1219, 
                           product(35) => n_1220, product(34) => n_1221, 
                           product(33) => n_1222, product(32) => n_1223, 
                           product(31) => N3296, product(30) => N3295, 
                           product(29) => N3294, product(28) => N3293, 
                           product(27) => N3292, product(26) => N3291, 
                           product(25) => N3290, product(24) => N3289, 
                           product(23) => N3288, product(22) => N3287, 
                           product(21) => N3286, product(20) => N3285, 
                           product(19) => N3284, product(18) => N3283, 
                           product(17) => N3282, product(16) => N3281, 
                           product(15) => N3280, product(14) => N3279, 
                           product(13) => N3278, product(12) => N3277, 
                           product(11) => N3276, product(10) => N3275, 
                           product(9) => N3274, product(8) => N3273, product(7)
                           => N3272, product(6) => N3271, product(5) => N3270, 
                           product(4) => N3269, product(3) => N3268, product(2)
                           => N3267, product(1) => N3266, product(0) => N3265);
   mult_21_C245 : gp_custom_DW_mult_tc_7 port map( a(31) => N3008, a(30) => 
                           N3007, a(29) => N3006, a(28) => N3005, a(27) => 
                           N3004, a(26) => N3003, a(25) => N3002, a(24) => 
                           N3001, a(23) => N3000, a(22) => N2999, a(21) => 
                           N2998, a(20) => N2997, a(19) => N2996, a(18) => 
                           N2995, a(17) => N2994, a(16) => N2993, a(15) => 
                           N2992, a(14) => N2991, a(13) => N2990, a(12) => 
                           N2989, a(11) => N2988, a(10) => N2987, a(9) => N2986
                           , a(8) => N2985, a(7) => N2984, a(6) => N2983, a(5) 
                           => N2982, a(4) => N2981, a(3) => N2980, a(2) => 
                           N2979, a(1) => N2978, a(0) => N2977, b(31) => N3168,
                           b(30) => N3167, b(29) => N3166, b(28) => N3165, 
                           b(27) => N3164, b(26) => N3163, b(25) => N3162, 
                           b(24) => N3161, b(23) => N3160, b(22) => N3159, 
                           b(21) => N3158, b(20) => N3157, b(19) => N3156, 
                           b(18) => N3155, b(17) => N3154, b(16) => N3153, 
                           b(15) => N3152, b(14) => N3151, b(13) => N3150, 
                           b(12) => N3149, b(11) => N3148, b(10) => N3147, b(9)
                           => N3146, b(8) => N3145, b(7) => N3144, b(6) => 
                           N3143, b(5) => N3142, b(4) => N3141, b(3) => N3140, 
                           b(2) => N3139, b(1) => N3138, b(0) => N3137, 
                           product(63) => n_1224, product(62) => n_1225, 
                           product(61) => n_1226, product(60) => n_1227, 
                           product(59) => n_1228, product(58) => n_1229, 
                           product(57) => n_1230, product(56) => n_1231, 
                           product(55) => n_1232, product(54) => n_1233, 
                           product(53) => n_1234, product(52) => n_1235, 
                           product(51) => n_1236, product(50) => n_1237, 
                           product(49) => n_1238, product(48) => n_1239, 
                           product(47) => n_1240, product(46) => n_1241, 
                           product(45) => n_1242, product(44) => n_1243, 
                           product(43) => n_1244, product(42) => n_1245, 
                           product(41) => n_1246, product(40) => n_1247, 
                           product(39) => n_1248, product(38) => n_1249, 
                           product(37) => n_1250, product(36) => n_1251, 
                           product(35) => n_1252, product(34) => n_1253, 
                           product(33) => n_1254, product(32) => n_1255, 
                           product(31) => N3328, product(30) => N3327, 
                           product(29) => N3326, product(28) => N3325, 
                           product(27) => N3324, product(26) => N3323, 
                           product(25) => N3322, product(24) => N3321, 
                           product(23) => N3320, product(22) => N3319, 
                           product(21) => N3318, product(20) => N3317, 
                           product(19) => N3316, product(18) => N3315, 
                           product(17) => N3314, product(16) => N3313, 
                           product(15) => N3312, product(14) => N3311, 
                           product(13) => N3310, product(12) => N3309, 
                           product(11) => N3308, product(10) => N3307, 
                           product(9) => N3306, product(8) => N3305, product(7)
                           => N3304, product(6) => N3303, product(5) => N3302, 
                           product(4) => N3301, product(3) => N3300, product(2)
                           => N3299, product(1) => N3298, product(0) => N3297);
   mult_21_C247 : gp_custom_DW_mult_tc_8 port map( a(31) => N3040, a(30) => 
                           N3039, a(29) => N3038, a(28) => N3037, a(27) => 
                           N3036, a(26) => N3035, a(25) => N3034, a(24) => 
                           N3033, a(23) => N3032, a(22) => N3031, a(21) => 
                           N3030, a(20) => N3029, a(19) => N3028, a(18) => 
                           N3027, a(17) => N3026, a(16) => N3025, a(15) => 
                           N3024, a(14) => N3023, a(13) => N3022, a(12) => 
                           N3021, a(11) => N3020, a(10) => N3019, a(9) => N3018
                           , a(8) => N3017, a(7) => N3016, a(6) => N3015, a(5) 
                           => N3014, a(4) => N3013, a(3) => N3012, a(2) => 
                           N3011, a(1) => N3010, a(0) => N3009, b(31) => n312, 
                           b(30) => n311, b(29) => n310, b(28) => n305, b(27) 
                           => n303, b(26) => n302, b(25) => n299, b(24) => n298
                           , b(23) => n297, b(22) => n296, b(21) => n295, b(20)
                           => n294, b(19) => n293, b(18) => n290, b(17) => n289
                           , b(16) => n292, b(15) => n291, b(14) => n273, b(13)
                           => n272, b(12) => n271, b(11) => n274, b(10) => n285
                           , b(9) => n281, b(8) => n280, b(7) => n279, b(6) => 
                           n278, b(5) => n282, b(4) => n287, b(3) => n286, b(2)
                           => n284, b(1) => n283, b(0) => n288, product(63) => 
                           n_1256, product(62) => n_1257, product(61) => n_1258
                           , product(60) => n_1259, product(59) => n_1260, 
                           product(58) => n_1261, product(57) => n_1262, 
                           product(56) => n_1263, product(55) => n_1264, 
                           product(54) => n_1265, product(53) => n_1266, 
                           product(52) => n_1267, product(51) => n_1268, 
                           product(50) => n_1269, product(49) => n_1270, 
                           product(48) => n_1271, product(47) => n_1272, 
                           product(46) => n_1273, product(45) => n_1274, 
                           product(44) => n_1275, product(43) => n_1276, 
                           product(42) => n_1277, product(41) => n_1278, 
                           product(40) => n_1279, product(39) => n_1280, 
                           product(38) => n_1281, product(37) => n_1282, 
                           product(36) => n_1283, product(35) => n_1284, 
                           product(34) => n_1285, product(33) => n_1286, 
                           product(32) => n_1287, product(31) => N3360, 
                           product(30) => N3359, product(29) => N3358, 
                           product(28) => N3357, product(27) => N3356, 
                           product(26) => N3355, product(25) => N3354, 
                           product(24) => N3353, product(23) => N3352, 
                           product(22) => N3351, product(21) => N3350, 
                           product(20) => N3349, product(19) => N3348, 
                           product(18) => N3347, product(17) => N3346, 
                           product(16) => N3345, product(15) => N3344, 
                           product(14) => N3343, product(13) => N3342, 
                           product(12) => N3341, product(11) => N3340, 
                           product(10) => N3339, product(9) => N3338, 
                           product(8) => N3337, product(7) => N3336, product(6)
                           => N3335, product(5) => N3334, product(4) => N3333, 
                           product(3) => N3332, product(2) => N3331, product(1)
                           => N3330, product(0) => N3329);
   mult_21_C249 : gp_custom_DW_mult_tc_9 port map( a(31) => N3072, a(30) => 
                           N3071, a(29) => N3070, a(28) => N3069, a(27) => 
                           N3068, a(26) => N3067, a(25) => N3066, a(24) => 
                           N3065, a(23) => N3064, a(22) => N3063, a(21) => 
                           N3062, a(20) => N3061, a(19) => N3060, a(18) => 
                           N3059, a(17) => N3058, a(16) => N3057, a(15) => 
                           N3056, a(14) => N3055, a(13) => N3054, a(12) => 
                           N3053, a(11) => N3052, a(10) => N3051, a(9) => N3050
                           , a(8) => N3049, a(7) => N3048, a(6) => N3047, a(5) 
                           => N3046, a(4) => N3045, a(3) => N3044, a(2) => 
                           N3043, a(1) => N3042, a(0) => N3041, b(31) => n312, 
                           b(30) => n311, b(29) => n310, b(28) => n305, b(27) 
                           => n303, b(26) => n302, b(25) => n299, b(24) => n298
                           , b(23) => n297, b(22) => n296, b(21) => n295, b(20)
                           => n294, b(19) => n293, b(18) => n290, b(17) => n289
                           , b(16) => n292, b(15) => n291, b(14) => n273, b(13)
                           => n272, b(12) => n271, b(11) => n274, b(10) => n285
                           , b(9) => n281, b(8) => n280, b(7) => n279, b(6) => 
                           n278, b(5) => n282, b(4) => n287, b(3) => n286, b(2)
                           => n284, b(1) => n283, b(0) => n288, product(63) => 
                           n_1288, product(62) => n_1289, product(61) => n_1290
                           , product(60) => n_1291, product(59) => n_1292, 
                           product(58) => n_1293, product(57) => n_1294, 
                           product(56) => n_1295, product(55) => n_1296, 
                           product(54) => n_1297, product(53) => n_1298, 
                           product(52) => n_1299, product(51) => n_1300, 
                           product(50) => n_1301, product(49) => n_1302, 
                           product(48) => n_1303, product(47) => n_1304, 
                           product(46) => n_1305, product(45) => n_1306, 
                           product(44) => n_1307, product(43) => n_1308, 
                           product(42) => n_1309, product(41) => n_1310, 
                           product(40) => n_1311, product(39) => n_1312, 
                           product(38) => n_1313, product(37) => n_1314, 
                           product(36) => n_1315, product(35) => n_1316, 
                           product(34) => n_1317, product(33) => n_1318, 
                           product(32) => n_1319, product(31) => N3392, 
                           product(30) => N3391, product(29) => N3390, 
                           product(28) => N3389, product(27) => N3388, 
                           product(26) => N3387, product(25) => N3386, 
                           product(24) => N3385, product(23) => N3384, 
                           product(22) => N3383, product(21) => N3382, 
                           product(20) => N3381, product(19) => N3380, 
                           product(18) => N3379, product(17) => N3378, 
                           product(16) => N3377, product(15) => N3376, 
                           product(14) => N3375, product(13) => N3374, 
                           product(12) => N3373, product(11) => N3372, 
                           product(10) => N3371, product(9) => N3370, 
                           product(8) => N3369, product(7) => N3368, product(6)
                           => N3367, product(5) => N3366, product(4) => N3365, 
                           product(3) => N3364, product(2) => N3363, product(1)
                           => N3362, product(0) => N3361);
   comp_res_reg_4_30_inst : DFFRPQ1 port map( D => N3391, CK => clk, RB => 
                           resetn, Q => comp_res_30_port);
   comp_res_reg_4_28_inst : DFFRPQ1 port map( D => N3389, CK => clk, RB => 
                           resetn, Q => comp_res_28_port);
   comp_res_reg_4_26_inst : DFFRPQ1 port map( D => N3387, CK => clk, RB => 
                           resetn, Q => comp_res_26_port);
   comp_res_reg_4_24_inst : DFFRPQ1 port map( D => N3385, CK => clk, RB => 
                           resetn, Q => comp_res_24_port);
   comp_res_reg_4_22_inst : DFFRPQ1 port map( D => N3383, CK => clk, RB => 
                           resetn, Q => comp_res_22_port);
   comp_res_reg_4_20_inst : DFFRPQ1 port map( D => N3381, CK => clk, RB => 
                           resetn, Q => comp_res_20_port);
   comp_res_reg_4_18_inst : DFFRPQ1 port map( D => N3379, CK => clk, RB => 
                           resetn, Q => comp_res_18_port);
   comp_res_reg_4_16_inst : DFFRPQ1 port map( D => N3377, CK => clk, RB => 
                           resetn, Q => comp_res_16_port);
   comp_res_reg_4_14_inst : DFFRPQ1 port map( D => N3375, CK => clk, RB => 
                           resetn, Q => comp_res_14_port);
   comp_res_reg_4_12_inst : DFFRPQ1 port map( D => N3373, CK => clk, RB => 
                           resetn, Q => comp_res_12_port);
   comp_res_reg_4_10_inst : DFFRPQ1 port map( D => N3371, CK => clk, RB => 
                           resetn, Q => comp_res_10_port);
   comp_res_reg_4_8_inst : DFFRPQ1 port map( D => N3369, CK => clk, RB => 
                           resetn, Q => comp_res_8_port);
   comp_res_reg_4_6_inst : DFFRPQ1 port map( D => N3367, CK => clk, RB => 
                           resetn, Q => comp_res_6_port);
   comp_res_reg_4_4_inst : DFFRPQ1 port map( D => N3365, CK => clk, RB => 
                           resetn, Q => comp_res_4_port);
   comp_res_reg_4_2_inst : DFFRPQ1 port map( D => N3363, CK => clk, RB => 
                           resetn, Q => comp_res_2_port);
   comp_res_reg_4_0_inst : DFFRPQ1 port map( D => N3361, CK => clk, RB => 
                           resetn, Q => comp_res_0_port);
   comp_res_reg_4_31_inst : DFFRPQ1 port map( D => N3392, CK => clk, RB => 
                           resetn, Q => comp_res_31_port);
   comp_res_reg_4_29_inst : DFFRPQ1 port map( D => N3390, CK => clk, RB => 
                           resetn, Q => comp_res_29_port);
   comp_res_reg_4_27_inst : DFFRPQ1 port map( D => N3388, CK => clk, RB => 
                           resetn, Q => comp_res_27_port);
   comp_res_reg_4_25_inst : DFFRPQ1 port map( D => N3386, CK => clk, RB => 
                           resetn, Q => comp_res_25_port);
   comp_res_reg_4_23_inst : DFFRPQ1 port map( D => N3384, CK => clk, RB => 
                           resetn, Q => comp_res_23_port);
   comp_res_reg_4_21_inst : DFFRPQ1 port map( D => N3382, CK => clk, RB => 
                           resetn, Q => comp_res_21_port);
   comp_res_reg_4_19_inst : DFFRPQ1 port map( D => N3380, CK => clk, RB => 
                           resetn, Q => comp_res_19_port);
   comp_res_reg_4_17_inst : DFFRPQ1 port map( D => N3378, CK => clk, RB => 
                           resetn, Q => comp_res_17_port);
   comp_res_reg_4_15_inst : DFFRPQ1 port map( D => N3376, CK => clk, RB => 
                           resetn, Q => comp_res_15_port);
   comp_res_reg_4_13_inst : DFFRPQ1 port map( D => N3374, CK => clk, RB => 
                           resetn, Q => comp_res_13_port);
   comp_res_reg_4_11_inst : DFFRPQ1 port map( D => N3372, CK => clk, RB => 
                           resetn, Q => comp_res_11_port);
   comp_res_reg_4_9_inst : DFFRPQ1 port map( D => N3370, CK => clk, RB => 
                           resetn, Q => comp_res_9_port);
   comp_res_reg_4_7_inst : DFFRPQ1 port map( D => N3368, CK => clk, RB => 
                           resetn, Q => comp_res_7_port);
   comp_res_reg_4_5_inst : DFFRPQ1 port map( D => N3366, CK => clk, RB => 
                           resetn, Q => comp_res_5_port);
   comp_res_reg_4_3_inst : DFFRPQ1 port map( D => N3364, CK => clk, RB => 
                           resetn, Q => comp_res_3_port);
   comp_res_reg_4_1_inst : DFFRPQ1 port map( D => N3362, CK => clk, RB => 
                           resetn, Q => comp_res_1_port);
   comp_res_reg_3_30_inst : DFFRPQ1 port map( D => N3359, CK => clk, RB => 
                           resetn, Q => comp_res_62_port);
   comp_res_reg_3_28_inst : DFFRPQ1 port map( D => N3357, CK => clk, RB => 
                           resetn, Q => comp_res_60_port);
   comp_res_reg_3_26_inst : DFFRPQ1 port map( D => N3355, CK => clk, RB => 
                           resetn, Q => comp_res_58_port);
   comp_res_reg_3_24_inst : DFFRPQ1 port map( D => N3353, CK => clk, RB => 
                           resetn, Q => comp_res_56_port);
   comp_res_reg_3_22_inst : DFFRPQ1 port map( D => N3351, CK => clk, RB => 
                           resetn, Q => comp_res_54_port);
   comp_res_reg_3_20_inst : DFFRPQ1 port map( D => N3349, CK => clk, RB => 
                           resetn, Q => comp_res_52_port);
   comp_res_reg_3_18_inst : DFFRPQ1 port map( D => N3347, CK => clk, RB => 
                           resetn, Q => comp_res_50_port);
   comp_res_reg_3_16_inst : DFFRPQ1 port map( D => N3345, CK => clk, RB => 
                           resetn, Q => comp_res_48_port);
   comp_res_reg_3_14_inst : DFFRPQ1 port map( D => N3343, CK => clk, RB => 
                           resetn, Q => comp_res_46_port);
   comp_res_reg_3_12_inst : DFFRPQ1 port map( D => N3341, CK => clk, RB => 
                           resetn, Q => comp_res_44_port);
   comp_res_reg_3_10_inst : DFFRPQ1 port map( D => N3339, CK => clk, RB => 
                           resetn, Q => comp_res_42_port);
   comp_res_reg_3_8_inst : DFFRPQ1 port map( D => N3337, CK => clk, RB => 
                           resetn, Q => comp_res_40_port);
   comp_res_reg_3_6_inst : DFFRPQ1 port map( D => N3335, CK => clk, RB => 
                           resetn, Q => comp_res_38_port);
   comp_res_reg_3_4_inst : DFFRPQ1 port map( D => N3333, CK => clk, RB => 
                           resetn, Q => comp_res_36_port);
   comp_res_reg_3_2_inst : DFFRPQ1 port map( D => N3331, CK => clk, RB => 
                           resetn, Q => comp_res_34_port);
   comp_res_reg_2_30_inst : DFFRPQ1 port map( D => N3327, CK => clk, RB => 
                           resetn, Q => comp_res_94_port);
   comp_res_reg_2_28_inst : DFFRPQ1 port map( D => N3325, CK => clk, RB => 
                           resetn, Q => comp_res_92_port);
   comp_res_reg_2_26_inst : DFFRPQ1 port map( D => N3323, CK => clk, RB => 
                           resetn, Q => comp_res_90_port);
   comp_res_reg_2_24_inst : DFFRPQ1 port map( D => N3321, CK => clk, RB => 
                           resetn, Q => comp_res_88_port);
   comp_res_reg_2_22_inst : DFFRPQ1 port map( D => N3319, CK => clk, RB => 
                           resetn, Q => comp_res_86_port);
   comp_res_reg_2_20_inst : DFFRPQ1 port map( D => N3317, CK => clk, RB => 
                           resetn, Q => comp_res_84_port);
   comp_res_reg_2_18_inst : DFFRPQ1 port map( D => N3315, CK => clk, RB => 
                           resetn, Q => comp_res_82_port);
   comp_res_reg_2_16_inst : DFFRPQ1 port map( D => N3313, CK => clk, RB => 
                           resetn, Q => comp_res_80_port);
   comp_res_reg_2_14_inst : DFFRPQ1 port map( D => N3311, CK => clk, RB => 
                           resetn, Q => comp_res_78_port);
   comp_res_reg_2_12_inst : DFFRPQ1 port map( D => N3309, CK => clk, RB => 
                           resetn, Q => comp_res_76_port);
   comp_res_reg_2_10_inst : DFFRPQ1 port map( D => N3307, CK => clk, RB => 
                           resetn, Q => comp_res_74_port);
   comp_res_reg_2_8_inst : DFFRPQ1 port map( D => N3305, CK => clk, RB => 
                           resetn, Q => comp_res_72_port);
   comp_res_reg_2_6_inst : DFFRPQ1 port map( D => N3303, CK => clk, RB => 
                           resetn, Q => comp_res_70_port);
   comp_res_reg_2_4_inst : DFFRPQ1 port map( D => N3301, CK => clk, RB => 
                           resetn, Q => comp_res_68_port);
   comp_res_reg_2_2_inst : DFFRPQ1 port map( D => N3299, CK => clk, RB => 
                           resetn, Q => comp_res_66_port);
   comp_res_reg_1_30_inst : DFFRPQ1 port map( D => N3295, CK => clk, RB => 
                           resetn, Q => comp_res_126_port);
   comp_res_reg_1_28_inst : DFFRPQ1 port map( D => N3293, CK => clk, RB => 
                           resetn, Q => comp_res_124_port);
   comp_res_reg_1_26_inst : DFFRPQ1 port map( D => N3291, CK => clk, RB => 
                           resetn, Q => comp_res_122_port);
   comp_res_reg_1_24_inst : DFFRPQ1 port map( D => N3289, CK => clk, RB => 
                           resetn, Q => comp_res_120_port);
   comp_res_reg_1_22_inst : DFFRPQ1 port map( D => N3287, CK => clk, RB => 
                           resetn, Q => comp_res_118_port);
   comp_res_reg_1_20_inst : DFFRPQ1 port map( D => N3285, CK => clk, RB => 
                           resetn, Q => comp_res_116_port);
   comp_res_reg_1_18_inst : DFFRPQ1 port map( D => N3283, CK => clk, RB => 
                           resetn, Q => comp_res_114_port);
   comp_res_reg_1_16_inst : DFFRPQ1 port map( D => N3281, CK => clk, RB => 
                           resetn, Q => comp_res_112_port);
   comp_res_reg_1_14_inst : DFFRPQ1 port map( D => N3279, CK => clk, RB => 
                           resetn, Q => comp_res_110_port);
   comp_res_reg_1_12_inst : DFFRPQ1 port map( D => N3277, CK => clk, RB => 
                           resetn, Q => comp_res_108_port);
   comp_res_reg_1_10_inst : DFFRPQ1 port map( D => N3275, CK => clk, RB => 
                           resetn, Q => comp_res_106_port);
   comp_res_reg_1_8_inst : DFFRPQ1 port map( D => N3273, CK => clk, RB => 
                           resetn, Q => comp_res_104_port);
   comp_res_reg_1_6_inst : DFFRPQ1 port map( D => N3271, CK => clk, RB => 
                           resetn, Q => comp_res_102_port);
   comp_res_reg_1_4_inst : DFFRPQ1 port map( D => N3269, CK => clk, RB => 
                           resetn, Q => comp_res_100_port);
   comp_res_reg_1_2_inst : DFFRPQ1 port map( D => N3267, CK => clk, RB => 
                           resetn, Q => comp_res_98_port);
   comp_res_reg_0_30_inst : DFFRPQ1 port map( D => N3263, CK => clk, RB => 
                           resetn, Q => comp_res_158_port);
   comp_res_reg_0_28_inst : DFFRPQ1 port map( D => N3261, CK => clk, RB => 
                           resetn, Q => comp_res_156_port);
   comp_res_reg_0_26_inst : DFFRPQ1 port map( D => N3259, CK => clk, RB => 
                           resetn, Q => comp_res_154_port);
   comp_res_reg_0_24_inst : DFFRPQ1 port map( D => N3257, CK => clk, RB => 
                           resetn, Q => comp_res_152_port);
   comp_res_reg_0_22_inst : DFFRPQ1 port map( D => N3255, CK => clk, RB => 
                           resetn, Q => comp_res_150_port);
   comp_res_reg_0_20_inst : DFFRPQ1 port map( D => N3253, CK => clk, RB => 
                           resetn, Q => comp_res_148_port);
   comp_res_reg_0_18_inst : DFFRPQ1 port map( D => N3251, CK => clk, RB => 
                           resetn, Q => comp_res_146_port);
   comp_res_reg_0_16_inst : DFFRPQ1 port map( D => N3249, CK => clk, RB => 
                           resetn, Q => comp_res_144_port);
   comp_res_reg_0_14_inst : DFFRPQ1 port map( D => N3247, CK => clk, RB => 
                           resetn, Q => comp_res_142_port);
   comp_res_reg_0_12_inst : DFFRPQ1 port map( D => N3245, CK => clk, RB => 
                           resetn, Q => comp_res_140_port);
   comp_res_reg_0_10_inst : DFFRPQ1 port map( D => N3243, CK => clk, RB => 
                           resetn, Q => comp_res_138_port);
   comp_res_reg_0_8_inst : DFFRPQ1 port map( D => N3241, CK => clk, RB => 
                           resetn, Q => comp_res_136_port);
   comp_res_reg_0_6_inst : DFFRPQ1 port map( D => N3239, CK => clk, RB => 
                           resetn, Q => comp_res_134_port);
   comp_res_reg_0_4_inst : DFFRPQ1 port map( D => N3237, CK => clk, RB => 
                           resetn, Q => comp_res_132_port);
   comp_res_reg_0_2_inst : DFFRPQ1 port map( D => N3235, CK => clk, RB => 
                           resetn, Q => comp_res_130_port);
   comp_res_reg_3_0_inst : DFFRPQ1 port map( D => N3329, CK => clk, RB => 
                           resetn, Q => comp_res_32_port);
   comp_res_reg_2_0_inst : DFFRPQ1 port map( D => N3297, CK => clk, RB => 
                           resetn, Q => comp_res_64_port);
   comp_res_reg_1_0_inst : DFFRPQ1 port map( D => N3265, CK => clk, RB => 
                           resetn, Q => comp_res_96_port);
   comp_res_reg_0_0_inst : DFFRPQ1 port map( D => N3233, CK => clk, RB => 
                           resetn, Q => comp_res_128_port);
   in_buf_reg_7_31_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n176,
                           CK => clk, RB => resetn, Q => in_buf_31_port);
   in_buf_reg_7_29_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n176,
                           CK => clk, RB => resetn, Q => in_buf_29_port);
   in_buf_reg_7_27_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n176,
                           CK => clk, RB => resetn, Q => in_buf_27_port);
   in_buf_reg_7_25_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n176, 
                           CK => clk, RB => resetn, Q => in_buf_25_port);
   in_buf_reg_7_23_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n176, 
                           CK => clk, RB => resetn, Q => in_buf_23_port);
   in_buf_reg_7_21_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n176, 
                           CK => clk, RB => resetn, Q => in_buf_21_port);
   in_buf_reg_7_19_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n176, 
                           CK => clk, RB => resetn, Q => in_buf_19_port);
   in_buf_reg_7_17_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n176, 
                           CK => clk, RB => resetn, Q => in_buf_17_port);
   in_buf_reg_7_15_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n177,
                           CK => clk, RB => resetn, Q => in_buf_15_port);
   in_buf_reg_7_13_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n177,
                           CK => clk, RB => resetn, Q => in_buf_13_port);
   in_buf_reg_7_11_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n177,
                           CK => clk, RB => resetn, Q => in_buf_11_port);
   in_buf_reg_7_9_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n177, 
                           CK => clk, RB => resetn, Q => in_buf_9_port);
   in_buf_reg_7_7_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n177, 
                           CK => clk, RB => resetn, Q => in_buf_7_port);
   in_buf_reg_7_5_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n177, 
                           CK => clk, RB => resetn, Q => in_buf_5_port);
   in_buf_reg_7_3_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n177, 
                           CK => clk, RB => resetn, Q => in_buf_3_port);
   in_buf_reg_7_1_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n177, 
                           CK => clk, RB => resetn, Q => in_buf_1_port);
   comp_res_reg_3_31_inst : DFFRPQ1 port map( D => N3360, CK => clk, RB => 
                           resetn, Q => comp_res_63_port);
   comp_res_reg_3_29_inst : DFFRPQ1 port map( D => N3358, CK => clk, RB => 
                           resetn, Q => comp_res_61_port);
   comp_res_reg_3_27_inst : DFFRPQ1 port map( D => N3356, CK => clk, RB => 
                           resetn, Q => comp_res_59_port);
   comp_res_reg_3_25_inst : DFFRPQ1 port map( D => N3354, CK => clk, RB => 
                           resetn, Q => comp_res_57_port);
   comp_res_reg_3_23_inst : DFFRPQ1 port map( D => N3352, CK => clk, RB => 
                           resetn, Q => comp_res_55_port);
   comp_res_reg_3_21_inst : DFFRPQ1 port map( D => N3350, CK => clk, RB => 
                           resetn, Q => comp_res_53_port);
   comp_res_reg_3_19_inst : DFFRPQ1 port map( D => N3348, CK => clk, RB => 
                           resetn, Q => comp_res_51_port);
   comp_res_reg_3_17_inst : DFFRPQ1 port map( D => N3346, CK => clk, RB => 
                           resetn, Q => comp_res_49_port);
   comp_res_reg_3_15_inst : DFFRPQ1 port map( D => N3344, CK => clk, RB => 
                           resetn, Q => comp_res_47_port);
   comp_res_reg_3_13_inst : DFFRPQ1 port map( D => N3342, CK => clk, RB => 
                           resetn, Q => comp_res_45_port);
   comp_res_reg_3_11_inst : DFFRPQ1 port map( D => N3340, CK => clk, RB => 
                           resetn, Q => comp_res_43_port);
   comp_res_reg_3_9_inst : DFFRPQ1 port map( D => N3338, CK => clk, RB => 
                           resetn, Q => comp_res_41_port);
   comp_res_reg_3_7_inst : DFFRPQ1 port map( D => N3336, CK => clk, RB => 
                           resetn, Q => comp_res_39_port);
   comp_res_reg_3_5_inst : DFFRPQ1 port map( D => N3334, CK => clk, RB => 
                           resetn, Q => comp_res_37_port);
   comp_res_reg_3_3_inst : DFFRPQ1 port map( D => N3332, CK => clk, RB => 
                           resetn, Q => comp_res_35_port);
   comp_res_reg_3_1_inst : DFFRPQ1 port map( D => N3330, CK => clk, RB => 
                           resetn, Q => comp_res_33_port);
   comp_res_reg_2_31_inst : DFFRPQ1 port map( D => N3328, CK => clk, RB => 
                           resetn, Q => comp_res_95_port);
   comp_res_reg_2_29_inst : DFFRPQ1 port map( D => N3326, CK => clk, RB => 
                           resetn, Q => comp_res_93_port);
   comp_res_reg_2_27_inst : DFFRPQ1 port map( D => N3324, CK => clk, RB => 
                           resetn, Q => comp_res_91_port);
   comp_res_reg_2_25_inst : DFFRPQ1 port map( D => N3322, CK => clk, RB => 
                           resetn, Q => comp_res_89_port);
   comp_res_reg_2_23_inst : DFFRPQ1 port map( D => N3320, CK => clk, RB => 
                           resetn, Q => comp_res_87_port);
   comp_res_reg_2_21_inst : DFFRPQ1 port map( D => N3318, CK => clk, RB => 
                           resetn, Q => comp_res_85_port);
   comp_res_reg_2_19_inst : DFFRPQ1 port map( D => N3316, CK => clk, RB => 
                           resetn, Q => comp_res_83_port);
   comp_res_reg_2_17_inst : DFFRPQ1 port map( D => N3314, CK => clk, RB => 
                           resetn, Q => comp_res_81_port);
   comp_res_reg_2_15_inst : DFFRPQ1 port map( D => N3312, CK => clk, RB => 
                           resetn, Q => comp_res_79_port);
   comp_res_reg_2_13_inst : DFFRPQ1 port map( D => N3310, CK => clk, RB => 
                           resetn, Q => comp_res_77_port);
   comp_res_reg_2_11_inst : DFFRPQ1 port map( D => N3308, CK => clk, RB => 
                           resetn, Q => comp_res_75_port);
   comp_res_reg_2_9_inst : DFFRPQ1 port map( D => N3306, CK => clk, RB => 
                           resetn, Q => comp_res_73_port);
   comp_res_reg_2_7_inst : DFFRPQ1 port map( D => N3304, CK => clk, RB => 
                           resetn, Q => comp_res_71_port);
   comp_res_reg_2_5_inst : DFFRPQ1 port map( D => N3302, CK => clk, RB => 
                           resetn, Q => comp_res_69_port);
   comp_res_reg_2_3_inst : DFFRPQ1 port map( D => N3300, CK => clk, RB => 
                           resetn, Q => comp_res_67_port);
   comp_res_reg_2_1_inst : DFFRPQ1 port map( D => N3298, CK => clk, RB => 
                           resetn, Q => comp_res_65_port);
   in_buf_reg_3_31_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n168,
                           CK => clk, RB => resetn, Q => in_buf_159_port);
   in_buf_reg_3_29_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n168,
                           CK => clk, RB => resetn, Q => in_buf_157_port);
   in_buf_reg_3_27_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n168,
                           CK => clk, RB => resetn, Q => in_buf_155_port);
   in_buf_reg_3_25_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n168, 
                           CK => clk, RB => resetn, Q => in_buf_153_port);
   in_buf_reg_3_23_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n168, 
                           CK => clk, RB => resetn, Q => in_buf_151_port);
   in_buf_reg_3_21_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n168, 
                           CK => clk, RB => resetn, Q => in_buf_149_port);
   in_buf_reg_3_19_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n168, 
                           CK => clk, RB => resetn, Q => in_buf_147_port);
   in_buf_reg_3_17_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n168, 
                           CK => clk, RB => resetn, Q => in_buf_145_port);
   in_buf_reg_3_15_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n169,
                           CK => clk, RB => resetn, Q => in_buf_143_port);
   in_buf_reg_3_13_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n169,
                           CK => clk, RB => resetn, Q => in_buf_141_port);
   in_buf_reg_3_11_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n169,
                           CK => clk, RB => resetn, Q => in_buf_139_port);
   in_buf_reg_3_9_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n169, 
                           CK => clk, RB => resetn, Q => in_buf_137_port);
   in_buf_reg_3_7_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n169, 
                           CK => clk, RB => resetn, Q => in_buf_135_port);
   in_buf_reg_3_5_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n169, 
                           CK => clk, RB => resetn, Q => in_buf_133_port);
   in_buf_reg_3_3_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n169, 
                           CK => clk, RB => resetn, Q => in_buf_131_port);
   in_buf_reg_3_1_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n169, 
                           CK => clk, RB => resetn, Q => in_buf_129_port);
   in_buf_reg_2_31_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n166,
                           CK => clk, RB => resetn, Q => in_buf_191_port);
   in_buf_reg_2_29_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n166,
                           CK => clk, RB => resetn, Q => in_buf_189_port);
   in_buf_reg_2_27_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n166,
                           CK => clk, RB => resetn, Q => in_buf_187_port);
   in_buf_reg_2_25_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n166, 
                           CK => clk, RB => resetn, Q => in_buf_185_port);
   in_buf_reg_2_23_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n166, 
                           CK => clk, RB => resetn, Q => in_buf_183_port);
   in_buf_reg_2_21_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n166, 
                           CK => clk, RB => resetn, Q => in_buf_181_port);
   in_buf_reg_2_19_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n166, 
                           CK => clk, RB => resetn, Q => in_buf_179_port);
   in_buf_reg_2_17_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n166, 
                           CK => clk, RB => resetn, Q => in_buf_177_port);
   in_buf_reg_6_31_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n174,
                           CK => clk, RB => resetn, Q => in_buf_63_port);
   in_buf_reg_6_29_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n174,
                           CK => clk, RB => resetn, Q => in_buf_61_port);
   in_buf_reg_6_27_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n174,
                           CK => clk, RB => resetn, Q => in_buf_59_port);
   in_buf_reg_6_25_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n174, 
                           CK => clk, RB => resetn, Q => in_buf_57_port);
   in_buf_reg_6_23_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n174, 
                           CK => clk, RB => resetn, Q => in_buf_55_port);
   in_buf_reg_6_21_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n174, 
                           CK => clk, RB => resetn, Q => in_buf_53_port);
   in_buf_reg_6_19_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n174, 
                           CK => clk, RB => resetn, Q => in_buf_51_port);
   in_buf_reg_6_17_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n174, 
                           CK => clk, RB => resetn, Q => in_buf_49_port);
   in_buf_reg_2_15_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n167,
                           CK => clk, RB => resetn, Q => in_buf_175_port);
   in_buf_reg_2_13_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n167,
                           CK => clk, RB => resetn, Q => in_buf_173_port);
   in_buf_reg_2_11_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n167,
                           CK => clk, RB => resetn, Q => in_buf_171_port);
   in_buf_reg_2_9_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n167, 
                           CK => clk, RB => resetn, Q => in_buf_169_port);
   in_buf_reg_2_7_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n167, 
                           CK => clk, RB => resetn, Q => in_buf_167_port);
   in_buf_reg_2_5_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n167, 
                           CK => clk, RB => resetn, Q => in_buf_165_port);
   in_buf_reg_2_3_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n167, 
                           CK => clk, RB => resetn, Q => in_buf_163_port);
   in_buf_reg_2_1_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n167, 
                           CK => clk, RB => resetn, Q => in_buf_161_port);
   in_buf_reg_6_15_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n175,
                           CK => clk, RB => resetn, Q => in_buf_47_port);
   in_buf_reg_6_13_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n175,
                           CK => clk, RB => resetn, Q => in_buf_45_port);
   in_buf_reg_6_11_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n175,
                           CK => clk, RB => resetn, Q => in_buf_43_port);
   in_buf_reg_6_9_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n175, 
                           CK => clk, RB => resetn, Q => in_buf_41_port);
   in_buf_reg_6_7_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n175, 
                           CK => clk, RB => resetn, Q => in_buf_39_port);
   in_buf_reg_6_5_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n175, 
                           CK => clk, RB => resetn, Q => in_buf_37_port);
   in_buf_reg_6_3_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n175, 
                           CK => clk, RB => resetn, Q => in_buf_35_port);
   in_buf_reg_6_1_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n175, 
                           CK => clk, RB => resetn, Q => in_buf_33_port);
   in_buf_reg_5_31_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n172,
                           CK => clk, RB => resetn, Q => in_buf_95_port);
   in_buf_reg_5_29_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n172,
                           CK => clk, RB => resetn, Q => in_buf_93_port);
   in_buf_reg_5_27_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n172,
                           CK => clk, RB => resetn, Q => in_buf_91_port);
   in_buf_reg_5_25_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n172, 
                           CK => clk, RB => resetn, Q => in_buf_89_port);
   in_buf_reg_5_23_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n172, 
                           CK => clk, RB => resetn, Q => in_buf_87_port);
   in_buf_reg_5_21_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n172, 
                           CK => clk, RB => resetn, Q => in_buf_85_port);
   in_buf_reg_5_19_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n172, 
                           CK => clk, RB => resetn, Q => in_buf_83_port);
   in_buf_reg_5_17_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n172, 
                           CK => clk, RB => resetn, Q => in_buf_81_port);
   in_buf_reg_5_15_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n173,
                           CK => clk, RB => resetn, Q => in_buf_79_port);
   in_buf_reg_5_13_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n173,
                           CK => clk, RB => resetn, Q => in_buf_77_port);
   in_buf_reg_5_11_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n173,
                           CK => clk, RB => resetn, Q => in_buf_75_port);
   in_buf_reg_5_9_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n173, 
                           CK => clk, RB => resetn, Q => in_buf_73_port);
   in_buf_reg_5_7_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n173, 
                           CK => clk, RB => resetn, Q => in_buf_71_port);
   in_buf_reg_5_5_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n173, 
                           CK => clk, RB => resetn, Q => in_buf_69_port);
   in_buf_reg_5_3_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n173, 
                           CK => clk, RB => resetn, Q => in_buf_67_port);
   in_buf_reg_5_1_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n173, 
                           CK => clk, RB => resetn, Q => in_buf_65_port);
   comp_res_reg_1_31_inst : DFFRPQ1 port map( D => N3296, CK => clk, RB => 
                           resetn, Q => comp_res_127_port);
   comp_res_reg_1_29_inst : DFFRPQ1 port map( D => N3294, CK => clk, RB => 
                           resetn, Q => comp_res_125_port);
   comp_res_reg_1_27_inst : DFFRPQ1 port map( D => N3292, CK => clk, RB => 
                           resetn, Q => comp_res_123_port);
   comp_res_reg_1_25_inst : DFFRPQ1 port map( D => N3290, CK => clk, RB => 
                           resetn, Q => comp_res_121_port);
   comp_res_reg_1_23_inst : DFFRPQ1 port map( D => N3288, CK => clk, RB => 
                           resetn, Q => comp_res_119_port);
   comp_res_reg_1_21_inst : DFFRPQ1 port map( D => N3286, CK => clk, RB => 
                           resetn, Q => comp_res_117_port);
   comp_res_reg_1_19_inst : DFFRPQ1 port map( D => N3284, CK => clk, RB => 
                           resetn, Q => comp_res_115_port);
   comp_res_reg_1_17_inst : DFFRPQ1 port map( D => N3282, CK => clk, RB => 
                           resetn, Q => comp_res_113_port);
   comp_res_reg_1_15_inst : DFFRPQ1 port map( D => N3280, CK => clk, RB => 
                           resetn, Q => comp_res_111_port);
   comp_res_reg_1_13_inst : DFFRPQ1 port map( D => N3278, CK => clk, RB => 
                           resetn, Q => comp_res_109_port);
   comp_res_reg_1_11_inst : DFFRPQ1 port map( D => N3276, CK => clk, RB => 
                           resetn, Q => comp_res_107_port);
   comp_res_reg_1_9_inst : DFFRPQ1 port map( D => N3274, CK => clk, RB => 
                           resetn, Q => comp_res_105_port);
   comp_res_reg_1_7_inst : DFFRPQ1 port map( D => N3272, CK => clk, RB => 
                           resetn, Q => comp_res_103_port);
   comp_res_reg_1_5_inst : DFFRPQ1 port map( D => N3270, CK => clk, RB => 
                           resetn, Q => comp_res_101_port);
   comp_res_reg_1_3_inst : DFFRPQ1 port map( D => N3268, CK => clk, RB => 
                           resetn, Q => comp_res_99_port);
   comp_res_reg_1_1_inst : DFFRPQ1 port map( D => N3266, CK => clk, RB => 
                           resetn, Q => comp_res_97_port);
   comp_res_reg_0_31_inst : DFFRPQ1 port map( D => N3264, CK => clk, RB => 
                           resetn, Q => comp_res_159_port);
   comp_res_reg_0_29_inst : DFFRPQ1 port map( D => N3262, CK => clk, RB => 
                           resetn, Q => comp_res_157_port);
   comp_res_reg_0_27_inst : DFFRPQ1 port map( D => N3260, CK => clk, RB => 
                           resetn, Q => comp_res_155_port);
   comp_res_reg_0_25_inst : DFFRPQ1 port map( D => N3258, CK => clk, RB => 
                           resetn, Q => comp_res_153_port);
   comp_res_reg_0_23_inst : DFFRPQ1 port map( D => N3256, CK => clk, RB => 
                           resetn, Q => comp_res_151_port);
   comp_res_reg_0_21_inst : DFFRPQ1 port map( D => N3254, CK => clk, RB => 
                           resetn, Q => comp_res_149_port);
   comp_res_reg_0_19_inst : DFFRPQ1 port map( D => N3252, CK => clk, RB => 
                           resetn, Q => comp_res_147_port);
   comp_res_reg_0_17_inst : DFFRPQ1 port map( D => N3250, CK => clk, RB => 
                           resetn, Q => comp_res_145_port);
   comp_res_reg_0_15_inst : DFFRPQ1 port map( D => N3248, CK => clk, RB => 
                           resetn, Q => comp_res_143_port);
   comp_res_reg_0_13_inst : DFFRPQ1 port map( D => N3246, CK => clk, RB => 
                           resetn, Q => comp_res_141_port);
   comp_res_reg_0_11_inst : DFFRPQ1 port map( D => N3244, CK => clk, RB => 
                           resetn, Q => comp_res_139_port);
   comp_res_reg_0_9_inst : DFFRPQ1 port map( D => N3242, CK => clk, RB => 
                           resetn, Q => comp_res_137_port);
   comp_res_reg_0_7_inst : DFFRPQ1 port map( D => N3240, CK => clk, RB => 
                           resetn, Q => comp_res_135_port);
   comp_res_reg_0_5_inst : DFFRPQ1 port map( D => N3238, CK => clk, RB => 
                           resetn, Q => comp_res_133_port);
   comp_res_reg_0_3_inst : DFFRPQ1 port map( D => N3236, CK => clk, RB => 
                           resetn, Q => comp_res_131_port);
   comp_res_reg_0_1_inst : DFFRPQ1 port map( D => N3234, CK => clk, RB => 
                           resetn, Q => comp_res_129_port);
   in_buf_reg_1_31_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n164,
                           CK => clk, RB => resetn, Q => in_buf_223_port);
   in_buf_reg_1_29_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n164,
                           CK => clk, RB => resetn, Q => in_buf_221_port);
   in_buf_reg_1_27_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n164,
                           CK => clk, RB => resetn, Q => in_buf_219_port);
   in_buf_reg_1_25_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n164, 
                           CK => clk, RB => resetn, Q => in_buf_217_port);
   in_buf_reg_1_23_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n164, 
                           CK => clk, RB => resetn, Q => in_buf_215_port);
   in_buf_reg_1_21_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n164, 
                           CK => clk, RB => resetn, Q => in_buf_213_port);
   in_buf_reg_1_19_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n164, 
                           CK => clk, RB => resetn, Q => in_buf_211_port);
   in_buf_reg_1_17_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n164, 
                           CK => clk, RB => resetn, Q => in_buf_209_port);
   in_buf_reg_1_15_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n165,
                           CK => clk, RB => resetn, Q => in_buf_207_port);
   in_buf_reg_1_13_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n165,
                           CK => clk, RB => resetn, Q => in_buf_205_port);
   in_buf_reg_1_11_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n165,
                           CK => clk, RB => resetn, Q => in_buf_203_port);
   in_buf_reg_1_9_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n165, 
                           CK => clk, RB => resetn, Q => in_buf_201_port);
   in_buf_reg_1_7_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n165, 
                           CK => clk, RB => resetn, Q => in_buf_199_port);
   in_buf_reg_1_5_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n165, 
                           CK => clk, RB => resetn, Q => in_buf_197_port);
   in_buf_reg_1_3_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n165, 
                           CK => clk, RB => resetn, Q => in_buf_195_port);
   in_buf_reg_1_1_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n165, 
                           CK => clk, RB => resetn, Q => in_buf_193_port);
   in_buf_reg_4_31_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n170,
                           CK => clk, RB => resetn, Q => in_buf_127_port);
   in_buf_reg_4_29_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n170,
                           CK => clk, RB => resetn, Q => in_buf_125_port);
   in_buf_reg_4_27_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n170,
                           CK => clk, RB => resetn, Q => in_buf_123_port);
   in_buf_reg_4_25_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n170, 
                           CK => clk, RB => resetn, Q => in_buf_121_port);
   in_buf_reg_4_23_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n170, 
                           CK => clk, RB => resetn, Q => in_buf_119_port);
   in_buf_reg_4_21_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n170, 
                           CK => clk, RB => resetn, Q => in_buf_117_port);
   in_buf_reg_4_19_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n170, 
                           CK => clk, RB => resetn, Q => in_buf_115_port);
   in_buf_reg_4_17_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n170, 
                           CK => clk, RB => resetn, Q => in_buf_113_port);
   in_buf_reg_0_31_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n162,
                           CK => clk, RB => resetn, Q => in_buf_255_port);
   in_buf_reg_0_29_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n162,
                           CK => clk, RB => resetn, Q => in_buf_253_port);
   in_buf_reg_0_27_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n162,
                           CK => clk, RB => resetn, Q => in_buf_251_port);
   in_buf_reg_0_25_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n162, 
                           CK => clk, RB => resetn, Q => in_buf_249_port);
   in_buf_reg_0_23_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n162, 
                           CK => clk, RB => resetn, Q => in_buf_247_port);
   in_buf_reg_0_21_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n162, 
                           CK => clk, RB => resetn, Q => in_buf_245_port);
   in_buf_reg_0_19_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n162, 
                           CK => clk, RB => resetn, Q => in_buf_243_port);
   in_buf_reg_0_17_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n162, 
                           CK => clk, RB => resetn, Q => in_buf_241_port);
   in_buf_reg_0_15_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n163,
                           CK => clk, RB => resetn, Q => in_buf_239_port);
   in_buf_reg_0_13_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n163,
                           CK => clk, RB => resetn, Q => in_buf_237_port);
   in_buf_reg_0_11_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n163,
                           CK => clk, RB => resetn, Q => in_buf_235_port);
   in_buf_reg_0_9_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n163, 
                           CK => clk, RB => resetn, Q => in_buf_233_port);
   in_buf_reg_0_7_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n163, 
                           CK => clk, RB => resetn, Q => in_buf_231_port);
   in_buf_reg_0_5_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n163, 
                           CK => clk, RB => resetn, Q => in_buf_229_port);
   in_buf_reg_0_3_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n163, 
                           CK => clk, RB => resetn, Q => in_buf_227_port);
   in_buf_reg_0_1_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n163, 
                           CK => clk, RB => resetn, Q => in_buf_225_port);
   in_buf_reg_4_15_inst : DFERPQ1 port map( D => siso_data_in(15), CEB => n171,
                           CK => clk, RB => resetn, Q => in_buf_111_port);
   in_buf_reg_4_13_inst : DFERPQ1 port map( D => siso_data_in(13), CEB => n171,
                           CK => clk, RB => resetn, Q => in_buf_109_port);
   in_buf_reg_4_11_inst : DFERPQ1 port map( D => siso_data_in(11), CEB => n171,
                           CK => clk, RB => resetn, Q => in_buf_107_port);
   in_buf_reg_4_9_inst : DFERPQ1 port map( D => siso_data_in(9), CEB => n171, 
                           CK => clk, RB => resetn, Q => in_buf_105_port);
   in_buf_reg_4_7_inst : DFERPQ1 port map( D => siso_data_in(7), CEB => n171, 
                           CK => clk, RB => resetn, Q => in_buf_103_port);
   in_buf_reg_4_5_inst : DFERPQ1 port map( D => siso_data_in(5), CEB => n171, 
                           CK => clk, RB => resetn, Q => in_buf_101_port);
   in_buf_reg_4_3_inst : DFERPQ1 port map( D => siso_data_in(3), CEB => n171, 
                           CK => clk, RB => resetn, Q => in_buf_99_port);
   in_buf_reg_4_1_inst : DFERPQ1 port map( D => siso_data_in(1), CEB => n171, 
                           CK => clk, RB => resetn, Q => in_buf_97_port);
   in_buf_reg_7_30_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n176,
                           CK => clk, RB => resetn, Q => in_buf_30_port);
   in_buf_reg_7_28_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n176,
                           CK => clk, RB => resetn, Q => in_buf_28_port);
   in_buf_reg_7_26_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n176,
                           CK => clk, RB => resetn, Q => in_buf_26_port);
   in_buf_reg_7_24_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n176, 
                           CK => clk, RB => resetn, Q => in_buf_24_port);
   in_buf_reg_7_22_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n176, 
                           CK => clk, RB => resetn, Q => in_buf_22_port);
   in_buf_reg_7_20_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n176, 
                           CK => clk, RB => resetn, Q => in_buf_20_port);
   in_buf_reg_7_18_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n176, 
                           CK => clk, RB => resetn, Q => in_buf_18_port);
   in_buf_reg_7_16_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n176, 
                           CK => clk, RB => resetn, Q => in_buf_16_port);
   in_buf_reg_7_14_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n177,
                           CK => clk, RB => resetn, Q => in_buf_14_port);
   in_buf_reg_7_12_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n177,
                           CK => clk, RB => resetn, Q => in_buf_12_port);
   in_buf_reg_7_10_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n177,
                           CK => clk, RB => resetn, Q => in_buf_10_port);
   in_buf_reg_7_8_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n177, 
                           CK => clk, RB => resetn, Q => in_buf_8_port);
   in_buf_reg_7_6_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n177, 
                           CK => clk, RB => resetn, Q => in_buf_6_port);
   in_buf_reg_7_4_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n177, 
                           CK => clk, RB => resetn, Q => in_buf_4_port);
   in_buf_reg_7_2_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n177, 
                           CK => clk, RB => resetn, Q => in_buf_2_port);
   in_trigger_reg : DFFRPQ1 port map( D => n241, CK => clk, RB => resetn, Q => 
                           in_trigger);
   in_buf_reg_3_30_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n168,
                           CK => clk, RB => resetn, Q => in_buf_158_port);
   in_buf_reg_3_28_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n168,
                           CK => clk, RB => resetn, Q => in_buf_156_port);
   in_buf_reg_3_26_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n168,
                           CK => clk, RB => resetn, Q => in_buf_154_port);
   in_buf_reg_3_24_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n168, 
                           CK => clk, RB => resetn, Q => in_buf_152_port);
   in_buf_reg_3_22_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n168, 
                           CK => clk, RB => resetn, Q => in_buf_150_port);
   in_buf_reg_3_20_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n168, 
                           CK => clk, RB => resetn, Q => in_buf_148_port);
   in_buf_reg_3_18_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n168, 
                           CK => clk, RB => resetn, Q => in_buf_146_port);
   in_buf_reg_3_16_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n168, 
                           CK => clk, RB => resetn, Q => in_buf_144_port);
   in_buf_reg_3_14_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n169,
                           CK => clk, RB => resetn, Q => in_buf_142_port);
   in_buf_reg_3_12_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n169,
                           CK => clk, RB => resetn, Q => in_buf_140_port);
   in_buf_reg_3_10_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n169,
                           CK => clk, RB => resetn, Q => in_buf_138_port);
   in_buf_reg_3_8_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n169, 
                           CK => clk, RB => resetn, Q => in_buf_136_port);
   in_buf_reg_3_6_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n169, 
                           CK => clk, RB => resetn, Q => in_buf_134_port);
   in_buf_reg_3_4_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n169, 
                           CK => clk, RB => resetn, Q => in_buf_132_port);
   in_buf_reg_3_2_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n169, 
                           CK => clk, RB => resetn, Q => in_buf_130_port);
   in_buf_reg_2_30_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n166,
                           CK => clk, RB => resetn, Q => in_buf_190_port);
   in_buf_reg_2_28_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n166,
                           CK => clk, RB => resetn, Q => in_buf_188_port);
   in_buf_reg_2_26_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n166,
                           CK => clk, RB => resetn, Q => in_buf_186_port);
   in_buf_reg_2_24_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n166, 
                           CK => clk, RB => resetn, Q => in_buf_184_port);
   in_buf_reg_2_22_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n166, 
                           CK => clk, RB => resetn, Q => in_buf_182_port);
   in_buf_reg_2_20_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n166, 
                           CK => clk, RB => resetn, Q => in_buf_180_port);
   in_buf_reg_2_18_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n166, 
                           CK => clk, RB => resetn, Q => in_buf_178_port);
   in_buf_reg_2_16_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n166, 
                           CK => clk, RB => resetn, Q => in_buf_176_port);
   in_buf_reg_6_30_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n174,
                           CK => clk, RB => resetn, Q => in_buf_62_port);
   in_buf_reg_6_28_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n174,
                           CK => clk, RB => resetn, Q => in_buf_60_port);
   in_buf_reg_6_26_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n174,
                           CK => clk, RB => resetn, Q => in_buf_58_port);
   in_buf_reg_6_24_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n174, 
                           CK => clk, RB => resetn, Q => in_buf_56_port);
   in_buf_reg_6_22_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n174, 
                           CK => clk, RB => resetn, Q => in_buf_54_port);
   in_buf_reg_6_20_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n174, 
                           CK => clk, RB => resetn, Q => in_buf_52_port);
   in_buf_reg_6_18_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n174, 
                           CK => clk, RB => resetn, Q => in_buf_50_port);
   in_buf_reg_6_16_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n174, 
                           CK => clk, RB => resetn, Q => in_buf_48_port);
   in_buf_reg_2_14_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n167,
                           CK => clk, RB => resetn, Q => in_buf_174_port);
   in_buf_reg_2_12_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n167,
                           CK => clk, RB => resetn, Q => in_buf_172_port);
   in_buf_reg_2_10_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n167,
                           CK => clk, RB => resetn, Q => in_buf_170_port);
   in_buf_reg_2_8_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n167, 
                           CK => clk, RB => resetn, Q => in_buf_168_port);
   in_buf_reg_2_6_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n167, 
                           CK => clk, RB => resetn, Q => in_buf_166_port);
   in_buf_reg_2_4_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n167, 
                           CK => clk, RB => resetn, Q => in_buf_164_port);
   in_buf_reg_2_2_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n167, 
                           CK => clk, RB => resetn, Q => in_buf_162_port);
   in_buf_reg_6_14_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n175,
                           CK => clk, RB => resetn, Q => in_buf_46_port);
   in_buf_reg_6_12_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n175,
                           CK => clk, RB => resetn, Q => in_buf_44_port);
   in_buf_reg_6_10_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n175,
                           CK => clk, RB => resetn, Q => in_buf_42_port);
   in_buf_reg_6_8_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n175, 
                           CK => clk, RB => resetn, Q => in_buf_40_port);
   in_buf_reg_6_6_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n175, 
                           CK => clk, RB => resetn, Q => in_buf_38_port);
   in_buf_reg_6_4_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n175, 
                           CK => clk, RB => resetn, Q => in_buf_36_port);
   in_buf_reg_6_2_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n175, 
                           CK => clk, RB => resetn, Q => in_buf_34_port);
   in_buf_reg_5_30_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n172,
                           CK => clk, RB => resetn, Q => in_buf_94_port);
   in_buf_reg_5_28_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n172,
                           CK => clk, RB => resetn, Q => in_buf_92_port);
   in_buf_reg_5_26_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n172,
                           CK => clk, RB => resetn, Q => in_buf_90_port);
   in_buf_reg_5_24_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n172, 
                           CK => clk, RB => resetn, Q => in_buf_88_port);
   in_buf_reg_5_22_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n172, 
                           CK => clk, RB => resetn, Q => in_buf_86_port);
   in_buf_reg_5_20_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n172, 
                           CK => clk, RB => resetn, Q => in_buf_84_port);
   in_buf_reg_5_18_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n172, 
                           CK => clk, RB => resetn, Q => in_buf_82_port);
   in_buf_reg_5_16_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n172, 
                           CK => clk, RB => resetn, Q => in_buf_80_port);
   in_buf_reg_5_14_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n173,
                           CK => clk, RB => resetn, Q => in_buf_78_port);
   in_buf_reg_5_12_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n173,
                           CK => clk, RB => resetn, Q => in_buf_76_port);
   in_buf_reg_5_10_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n173,
                           CK => clk, RB => resetn, Q => in_buf_74_port);
   in_buf_reg_5_8_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n173, 
                           CK => clk, RB => resetn, Q => in_buf_72_port);
   in_buf_reg_5_6_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n173, 
                           CK => clk, RB => resetn, Q => in_buf_70_port);
   in_buf_reg_5_4_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n173, 
                           CK => clk, RB => resetn, Q => in_buf_68_port);
   in_buf_reg_5_2_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n173, 
                           CK => clk, RB => resetn, Q => in_buf_66_port);
   in_buf_reg_7_0_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n177, 
                           CK => clk, RB => resetn, Q => in_buf_0_port);
   in_buf_reg_1_30_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n164,
                           CK => clk, RB => resetn, Q => in_buf_222_port);
   in_buf_reg_1_28_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n164,
                           CK => clk, RB => resetn, Q => in_buf_220_port);
   in_buf_reg_1_26_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n164,
                           CK => clk, RB => resetn, Q => in_buf_218_port);
   in_buf_reg_1_24_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n164, 
                           CK => clk, RB => resetn, Q => in_buf_216_port);
   in_buf_reg_1_22_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n164, 
                           CK => clk, RB => resetn, Q => in_buf_214_port);
   in_buf_reg_1_20_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n164, 
                           CK => clk, RB => resetn, Q => in_buf_212_port);
   in_buf_reg_1_18_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n164, 
                           CK => clk, RB => resetn, Q => in_buf_210_port);
   in_buf_reg_1_16_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n164, 
                           CK => clk, RB => resetn, Q => in_buf_208_port);
   in_buf_reg_1_14_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n165,
                           CK => clk, RB => resetn, Q => in_buf_206_port);
   in_buf_reg_1_12_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n165,
                           CK => clk, RB => resetn, Q => in_buf_204_port);
   in_buf_reg_1_10_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n165,
                           CK => clk, RB => resetn, Q => in_buf_202_port);
   in_buf_reg_1_8_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n165, 
                           CK => clk, RB => resetn, Q => in_buf_200_port);
   in_buf_reg_1_6_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n165, 
                           CK => clk, RB => resetn, Q => in_buf_198_port);
   in_buf_reg_1_4_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n165, 
                           CK => clk, RB => resetn, Q => in_buf_196_port);
   in_buf_reg_1_2_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n165, 
                           CK => clk, RB => resetn, Q => in_buf_194_port);
   in_buf_reg_4_30_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n170,
                           CK => clk, RB => resetn, Q => in_buf_126_port);
   in_buf_reg_4_28_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n170,
                           CK => clk, RB => resetn, Q => in_buf_124_port);
   in_buf_reg_4_26_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n170,
                           CK => clk, RB => resetn, Q => in_buf_122_port);
   in_buf_reg_4_24_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n170, 
                           CK => clk, RB => resetn, Q => in_buf_120_port);
   in_buf_reg_4_22_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n170, 
                           CK => clk, RB => resetn, Q => in_buf_118_port);
   in_buf_reg_4_20_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n170, 
                           CK => clk, RB => resetn, Q => in_buf_116_port);
   in_buf_reg_4_18_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n170, 
                           CK => clk, RB => resetn, Q => in_buf_114_port);
   in_buf_reg_4_16_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n170, 
                           CK => clk, RB => resetn, Q => in_buf_112_port);
   in_buf_reg_0_30_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n162,
                           CK => clk, RB => resetn, Q => in_buf_254_port);
   in_buf_reg_0_28_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n162,
                           CK => clk, RB => resetn, Q => in_buf_252_port);
   in_buf_reg_0_26_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n162,
                           CK => clk, RB => resetn, Q => in_buf_250_port);
   in_buf_reg_0_24_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n162, 
                           CK => clk, RB => resetn, Q => in_buf_248_port);
   in_buf_reg_0_22_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n162, 
                           CK => clk, RB => resetn, Q => in_buf_246_port);
   in_buf_reg_0_20_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n162, 
                           CK => clk, RB => resetn, Q => in_buf_244_port);
   in_buf_reg_0_18_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n162, 
                           CK => clk, RB => resetn, Q => in_buf_242_port);
   in_buf_reg_0_16_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n162, 
                           CK => clk, RB => resetn, Q => in_buf_240_port);
   in_buf_reg_0_14_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n163,
                           CK => clk, RB => resetn, Q => in_buf_238_port);
   in_buf_reg_0_12_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n163,
                           CK => clk, RB => resetn, Q => in_buf_236_port);
   in_buf_reg_0_10_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n163,
                           CK => clk, RB => resetn, Q => in_buf_234_port);
   in_buf_reg_0_8_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n163, 
                           CK => clk, RB => resetn, Q => in_buf_232_port);
   in_buf_reg_0_6_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n163, 
                           CK => clk, RB => resetn, Q => in_buf_230_port);
   in_buf_reg_0_4_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n163, 
                           CK => clk, RB => resetn, Q => in_buf_228_port);
   in_buf_reg_0_2_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n163, 
                           CK => clk, RB => resetn, Q => in_buf_226_port);
   in_buf_reg_4_14_inst : DFERPQ1 port map( D => siso_data_in(14), CEB => n171,
                           CK => clk, RB => resetn, Q => in_buf_110_port);
   in_buf_reg_4_12_inst : DFERPQ1 port map( D => siso_data_in(12), CEB => n171,
                           CK => clk, RB => resetn, Q => in_buf_108_port);
   in_buf_reg_4_10_inst : DFERPQ1 port map( D => siso_data_in(10), CEB => n171,
                           CK => clk, RB => resetn, Q => in_buf_106_port);
   in_buf_reg_4_8_inst : DFERPQ1 port map( D => siso_data_in(8), CEB => n171, 
                           CK => clk, RB => resetn, Q => in_buf_104_port);
   in_buf_reg_4_6_inst : DFERPQ1 port map( D => siso_data_in(6), CEB => n171, 
                           CK => clk, RB => resetn, Q => in_buf_102_port);
   in_buf_reg_4_4_inst : DFERPQ1 port map( D => siso_data_in(4), CEB => n171, 
                           CK => clk, RB => resetn, Q => in_buf_100_port);
   in_buf_reg_4_2_inst : DFERPQ1 port map( D => siso_data_in(2), CEB => n171, 
                           CK => clk, RB => resetn, Q => in_buf_98_port);
   in_buf_reg_3_0_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n169, 
                           CK => clk, RB => resetn, Q => in_buf_128_port);
   in_buf_reg_2_0_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n167, 
                           CK => clk, RB => resetn, Q => in_buf_160_port);
   in_buf_reg_6_0_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n175, 
                           CK => clk, RB => resetn, Q => in_buf_32_port);
   in_buf_reg_5_0_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n173, 
                           CK => clk, RB => resetn, Q => in_buf_64_port);
   out_buf_reg_7_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_15_port)
                           ;
   out_buf_reg_7_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_14_port)
                           ;
   out_buf_reg_7_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_13_port)
                           ;
   out_buf_reg_7_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_12_port)
                           ;
   out_buf_reg_7_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_11_port)
                           ;
   out_buf_reg_7_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_10_port)
                           ;
   out_buf_reg_7_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => n246,
                           CK => clk, RB => resetn, Q => out_buf_9_port);
   out_buf_reg_7_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => n246,
                           CK => clk, RB => resetn, Q => out_buf_8_port);
   out_buf_reg_7_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => n246,
                           CK => clk, RB => resetn, Q => out_buf_7_port);
   out_buf_reg_7_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => n246,
                           CK => clk, RB => resetn, Q => out_buf_6_port);
   out_buf_reg_7_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => n246,
                           CK => clk, RB => resetn, Q => out_buf_5_port);
   out_buf_reg_7_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => n246,
                           CK => clk, RB => resetn, Q => out_buf_4_port);
   out_buf_reg_7_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => n246,
                           CK => clk, RB => resetn, Q => out_buf_3_port);
   out_buf_reg_7_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => n246,
                           CK => clk, RB => resetn, Q => out_buf_2_port);
   out_buf_reg_7_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => n246,
                           CK => clk, RB => resetn, Q => out_buf_1_port);
   out_buf_reg_7_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => n246,
                           CK => clk, RB => resetn, Q => out_buf_0_port);
   in_buf_reg_1_0_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n165, 
                           CK => clk, RB => resetn, Q => in_buf_192_port);
   out_buf_reg_3_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n253, CK => clk, RB => resetn, Q => out_buf_143_port
                           );
   out_buf_reg_3_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n253, CK => clk, RB => resetn, Q => out_buf_142_port
                           );
   out_buf_reg_3_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n253, CK => clk, RB => resetn, Q => out_buf_141_port
                           );
   out_buf_reg_3_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n253, CK => clk, RB => resetn, Q => out_buf_140_port
                           );
   out_buf_reg_3_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n253, CK => clk, RB => resetn, Q => out_buf_139_port
                           );
   out_buf_reg_3_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n253, CK => clk, RB => resetn, Q => out_buf_138_port
                           );
   out_buf_reg_3_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => n253,
                           CK => clk, RB => resetn, Q => out_buf_137_port);
   out_buf_reg_3_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => n253,
                           CK => clk, RB => resetn, Q => out_buf_136_port);
   out_buf_reg_3_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => n253,
                           CK => clk, RB => resetn, Q => out_buf_135_port);
   out_buf_reg_3_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => n253,
                           CK => clk, RB => resetn, Q => out_buf_134_port);
   out_buf_reg_3_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => n253,
                           CK => clk, RB => resetn, Q => out_buf_133_port);
   out_buf_reg_3_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => n253,
                           CK => clk, RB => resetn, Q => out_buf_132_port);
   out_buf_reg_3_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => n253,
                           CK => clk, RB => resetn, Q => out_buf_131_port);
   out_buf_reg_3_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => n253,
                           CK => clk, RB => resetn, Q => out_buf_130_port);
   out_buf_reg_3_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => n253,
                           CK => clk, RB => resetn, Q => out_buf_129_port);
   out_buf_reg_3_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => n253,
                           CK => clk, RB => resetn, Q => out_buf_128_port);
   in_buf_reg_0_0_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n163, 
                           CK => clk, RB => resetn, Q => in_buf_224_port);
   in_buf_reg_4_0_inst : DFERPQ1 port map( D => siso_data_in(0), CEB => n171, 
                           CK => clk, RB => resetn, Q => in_buf_96_port);
   out_buf_reg_2_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_175_port
                           );
   out_buf_reg_2_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_174_port
                           );
   out_buf_reg_2_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_173_port
                           );
   out_buf_reg_2_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_172_port
                           );
   out_buf_reg_2_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_171_port
                           );
   out_buf_reg_2_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_170_port
                           );
   out_buf_reg_2_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => n252,
                           CK => clk, RB => resetn, Q => out_buf_169_port);
   out_buf_reg_2_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => n252,
                           CK => clk, RB => resetn, Q => out_buf_168_port);
   out_buf_reg_2_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => n252,
                           CK => clk, RB => resetn, Q => out_buf_167_port);
   out_buf_reg_2_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => n252,
                           CK => clk, RB => resetn, Q => out_buf_166_port);
   out_buf_reg_2_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => n252,
                           CK => clk, RB => resetn, Q => out_buf_165_port);
   out_buf_reg_2_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => n252,
                           CK => clk, RB => resetn, Q => out_buf_164_port);
   out_buf_reg_2_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => n252,
                           CK => clk, RB => resetn, Q => out_buf_163_port);
   out_buf_reg_2_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => n252,
                           CK => clk, RB => resetn, Q => out_buf_162_port);
   out_buf_reg_2_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => n252,
                           CK => clk, RB => resetn, Q => out_buf_161_port);
   out_buf_reg_2_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => n252,
                           CK => clk, RB => resetn, Q => out_buf_160_port);
   out_buf_reg_6_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_47_port)
                           ;
   out_buf_reg_6_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_46_port)
                           ;
   out_buf_reg_6_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_45_port)
                           ;
   out_buf_reg_6_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_44_port)
                           ;
   out_buf_reg_6_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_43_port)
                           ;
   out_buf_reg_6_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_42_port)
                           ;
   out_buf_reg_6_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => n251,
                           CK => clk, RB => resetn, Q => out_buf_41_port);
   out_buf_reg_6_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => n251,
                           CK => clk, RB => resetn, Q => out_buf_40_port);
   out_buf_reg_6_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => n251,
                           CK => clk, RB => resetn, Q => out_buf_39_port);
   out_buf_reg_6_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => n251,
                           CK => clk, RB => resetn, Q => out_buf_38_port);
   out_buf_reg_6_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => n251,
                           CK => clk, RB => resetn, Q => out_buf_37_port);
   out_buf_reg_6_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => n251,
                           CK => clk, RB => resetn, Q => out_buf_36_port);
   out_buf_reg_6_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => n251,
                           CK => clk, RB => resetn, Q => out_buf_35_port);
   out_buf_reg_6_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => n251,
                           CK => clk, RB => resetn, Q => out_buf_34_port);
   out_buf_reg_6_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => n251,
                           CK => clk, RB => resetn, Q => out_buf_33_port);
   out_buf_reg_6_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => n251,
                           CK => clk, RB => resetn, Q => out_buf_32_port);
   out_buf_reg_7_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_31_port)
                           ;
   out_buf_reg_7_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_30_port)
                           ;
   out_buf_reg_7_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_29_port)
                           ;
   out_buf_reg_7_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_28_port)
                           ;
   out_buf_reg_7_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_27_port)
                           ;
   out_buf_reg_7_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_26_port)
                           ;
   out_buf_reg_7_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_25_port)
                           ;
   out_buf_reg_7_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_24_port)
                           ;
   out_buf_reg_7_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_23_port)
                           ;
   out_buf_reg_7_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_22_port)
                           ;
   out_buf_reg_7_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_21_port)
                           ;
   out_buf_reg_7_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_20_port)
                           ;
   out_buf_reg_7_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_19_port)
                           ;
   out_buf_reg_7_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_18_port)
                           ;
   out_buf_reg_7_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_17_port)
                           ;
   out_buf_reg_7_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n246, CK => clk, RB => resetn, Q => out_buf_16_port)
                           ;
   out_buf_reg_5_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_79_port)
                           ;
   out_buf_reg_5_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_78_port)
                           ;
   out_buf_reg_5_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_77_port)
                           ;
   out_buf_reg_5_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_76_port)
                           ;
   out_buf_reg_5_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_75_port)
                           ;
   out_buf_reg_5_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_74_port)
                           ;
   out_buf_reg_5_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => n250,
                           CK => clk, RB => resetn, Q => out_buf_73_port);
   out_buf_reg_5_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => n250,
                           CK => clk, RB => resetn, Q => out_buf_72_port);
   out_buf_reg_5_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => n250,
                           CK => clk, RB => resetn, Q => out_buf_71_port);
   out_buf_reg_5_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => n250,
                           CK => clk, RB => resetn, Q => out_buf_70_port);
   out_buf_reg_5_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => n250,
                           CK => clk, RB => resetn, Q => out_buf_69_port);
   out_buf_reg_5_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => n250,
                           CK => clk, RB => resetn, Q => out_buf_68_port);
   out_buf_reg_5_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => n250,
                           CK => clk, RB => resetn, Q => out_buf_67_port);
   out_buf_reg_5_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => n250,
                           CK => clk, RB => resetn, Q => out_buf_66_port);
   out_buf_reg_5_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => n250,
                           CK => clk, RB => resetn, Q => out_buf_65_port);
   out_buf_reg_5_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => n250,
                           CK => clk, RB => resetn, Q => out_buf_64_port);
   out_buf_reg_3_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n253, CK => clk, RB => resetn, Q => out_buf_159_port
                           );
   out_buf_reg_3_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n253, CK => clk, RB => resetn, Q => out_buf_158_port
                           );
   out_buf_reg_3_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n253, CK => clk, RB => resetn, Q => out_buf_157_port
                           );
   out_buf_reg_3_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n253, CK => clk, RB => resetn, Q => out_buf_156_port
                           );
   out_buf_reg_3_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n253, CK => clk, RB => resetn, Q => out_buf_155_port
                           );
   out_buf_reg_3_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n253, CK => clk, RB => resetn, Q => out_buf_154_port
                           );
   out_buf_reg_3_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n253, CK => clk, RB => resetn, Q => out_buf_153_port
                           );
   out_buf_reg_3_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n253, CK => clk, RB => resetn, Q => out_buf_152_port
                           );
   out_buf_reg_3_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n253, CK => clk, RB => resetn, Q => out_buf_151_port
                           );
   out_buf_reg_3_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n253, CK => clk, RB => resetn, Q => out_buf_150_port
                           );
   out_buf_reg_3_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n253, CK => clk, RB => resetn, Q => out_buf_149_port
                           );
   out_buf_reg_3_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n253, CK => clk, RB => resetn, Q => out_buf_148_port
                           );
   out_buf_reg_3_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n253, CK => clk, RB => resetn, Q => out_buf_147_port
                           );
   out_buf_reg_3_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n253, CK => clk, RB => resetn, Q => out_buf_146_port
                           );
   out_buf_reg_3_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n253, CK => clk, RB => resetn, Q => out_buf_145_port
                           );
   out_buf_reg_3_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n253, CK => clk, RB => resetn, Q => out_buf_144_port
                           );
   out_buf_reg_1_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_207_port
                           );
   out_buf_reg_1_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_206_port
                           );
   out_buf_reg_1_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_205_port
                           );
   out_buf_reg_1_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_204_port
                           );
   out_buf_reg_1_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_203_port
                           );
   out_buf_reg_1_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_202_port
                           );
   out_buf_reg_1_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => n249,
                           CK => clk, RB => resetn, Q => out_buf_201_port);
   out_buf_reg_1_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => n249,
                           CK => clk, RB => resetn, Q => out_buf_200_port);
   out_buf_reg_1_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => n249,
                           CK => clk, RB => resetn, Q => out_buf_199_port);
   out_buf_reg_1_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => n249,
                           CK => clk, RB => resetn, Q => out_buf_198_port);
   out_buf_reg_1_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => n249,
                           CK => clk, RB => resetn, Q => out_buf_197_port);
   out_buf_reg_1_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => n249,
                           CK => clk, RB => resetn, Q => out_buf_196_port);
   out_buf_reg_1_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => n249,
                           CK => clk, RB => resetn, Q => out_buf_195_port);
   out_buf_reg_1_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => n249,
                           CK => clk, RB => resetn, Q => out_buf_194_port);
   out_buf_reg_1_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => n249,
                           CK => clk, RB => resetn, Q => out_buf_193_port);
   out_buf_reg_1_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => n249,
                           CK => clk, RB => resetn, Q => out_buf_192_port);
   out_buf_reg_2_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_191_port
                           );
   out_buf_reg_2_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_190_port
                           );
   out_buf_reg_2_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_189_port
                           );
   out_buf_reg_2_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_188_port
                           );
   out_buf_reg_2_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_187_port
                           );
   out_buf_reg_2_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_186_port
                           );
   out_buf_reg_2_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_185_port
                           );
   out_buf_reg_2_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_184_port
                           );
   out_buf_reg_2_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_183_port
                           );
   out_buf_reg_2_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_182_port
                           );
   out_buf_reg_2_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_181_port
                           );
   out_buf_reg_2_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_180_port
                           );
   out_buf_reg_2_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_179_port
                           );
   out_buf_reg_2_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_178_port
                           );
   out_buf_reg_2_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_177_port
                           );
   out_buf_reg_2_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n252, CK => clk, RB => resetn, Q => out_buf_176_port
                           );
   out_buf_reg_6_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_63_port)
                           ;
   out_buf_reg_6_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_62_port)
                           ;
   out_buf_reg_6_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_61_port)
                           ;
   out_buf_reg_6_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_60_port)
                           ;
   out_buf_reg_6_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_59_port)
                           ;
   out_buf_reg_6_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_58_port)
                           ;
   out_buf_reg_6_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_57_port)
                           ;
   out_buf_reg_6_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_56_port)
                           ;
   out_buf_reg_6_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_55_port)
                           ;
   out_buf_reg_6_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_54_port)
                           ;
   out_buf_reg_6_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_53_port)
                           ;
   out_buf_reg_6_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_52_port)
                           ;
   out_buf_reg_6_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_51_port)
                           ;
   out_buf_reg_6_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_50_port)
                           ;
   out_buf_reg_6_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_49_port)
                           ;
   out_buf_reg_6_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n251, CK => clk, RB => resetn, Q => out_buf_48_port)
                           ;
   out_buf_reg_0_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_239_port
                           );
   out_buf_reg_0_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_238_port
                           );
   out_buf_reg_0_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_237_port
                           );
   out_buf_reg_0_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_236_port
                           );
   out_buf_reg_0_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_235_port
                           );
   out_buf_reg_0_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_234_port
                           );
   out_buf_reg_0_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => n248,
                           CK => clk, RB => resetn, Q => out_buf_233_port);
   out_buf_reg_0_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => n248,
                           CK => clk, RB => resetn, Q => out_buf_232_port);
   out_buf_reg_0_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => n248,
                           CK => clk, RB => resetn, Q => out_buf_231_port);
   out_buf_reg_0_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => n248,
                           CK => clk, RB => resetn, Q => out_buf_230_port);
   out_buf_reg_0_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => n248,
                           CK => clk, RB => resetn, Q => out_buf_229_port);
   out_buf_reg_0_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => n248,
                           CK => clk, RB => resetn, Q => out_buf_228_port);
   out_buf_reg_0_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => n248,
                           CK => clk, RB => resetn, Q => out_buf_227_port);
   out_buf_reg_0_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => n248,
                           CK => clk, RB => resetn, Q => out_buf_226_port);
   out_buf_reg_0_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => n248,
                           CK => clk, RB => resetn, Q => out_buf_225_port);
   out_buf_reg_0_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => n248,
                           CK => clk, RB => resetn, Q => out_buf_224_port);
   out_buf_reg_4_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_111_port
                           );
   out_buf_reg_4_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_110_port
                           );
   out_buf_reg_4_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_109_port
                           );
   out_buf_reg_4_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_108_port
                           );
   out_buf_reg_4_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_107_port
                           );
   out_buf_reg_4_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_106_port
                           );
   out_buf_reg_4_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => n247,
                           CK => clk, RB => resetn, Q => out_buf_105_port);
   out_buf_reg_4_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => n247,
                           CK => clk, RB => resetn, Q => out_buf_104_port);
   out_buf_reg_4_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => n247,
                           CK => clk, RB => resetn, Q => out_buf_103_port);
   out_buf_reg_4_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => n247,
                           CK => clk, RB => resetn, Q => out_buf_102_port);
   out_buf_reg_4_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => n247,
                           CK => clk, RB => resetn, Q => out_buf_101_port);
   out_buf_reg_4_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => n247,
                           CK => clk, RB => resetn, Q => out_buf_100_port);
   out_buf_reg_4_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => n247,
                           CK => clk, RB => resetn, Q => out_buf_99_port);
   out_buf_reg_4_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => n247,
                           CK => clk, RB => resetn, Q => out_buf_98_port);
   out_buf_reg_4_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => n247,
                           CK => clk, RB => resetn, Q => out_buf_97_port);
   out_buf_reg_4_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => n247,
                           CK => clk, RB => resetn, Q => out_buf_96_port);
   out_buf_reg_5_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_95_port)
                           ;
   out_buf_reg_5_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_94_port)
                           ;
   out_buf_reg_5_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_93_port)
                           ;
   out_buf_reg_5_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_92_port)
                           ;
   out_buf_reg_5_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_91_port)
                           ;
   out_buf_reg_5_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_90_port)
                           ;
   out_buf_reg_5_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_89_port)
                           ;
   out_buf_reg_5_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_88_port)
                           ;
   out_buf_reg_5_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_87_port)
                           ;
   out_buf_reg_5_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_86_port)
                           ;
   out_buf_reg_5_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_85_port)
                           ;
   out_buf_reg_5_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_84_port)
                           ;
   out_buf_reg_5_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_83_port)
                           ;
   out_buf_reg_5_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_82_port)
                           ;
   out_buf_reg_5_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_81_port)
                           ;
   out_buf_reg_5_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n250, CK => clk, RB => resetn, Q => out_buf_80_port)
                           ;
   out_buf_reg_1_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_223_port
                           );
   out_buf_reg_1_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_222_port
                           );
   out_buf_reg_1_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_221_port
                           );
   out_buf_reg_1_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_220_port
                           );
   out_buf_reg_1_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_219_port
                           );
   out_buf_reg_1_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_218_port
                           );
   out_buf_reg_1_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_217_port
                           );
   out_buf_reg_1_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_216_port
                           );
   out_buf_reg_1_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_215_port
                           );
   out_buf_reg_1_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_214_port
                           );
   out_buf_reg_1_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_213_port
                           );
   out_buf_reg_1_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_212_port
                           );
   out_buf_reg_1_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_211_port
                           );
   out_buf_reg_1_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_210_port
                           );
   out_buf_reg_1_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_209_port
                           );
   out_buf_reg_1_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n249, CK => clk, RB => resetn, Q => out_buf_208_port
                           );
   out_buf_reg_0_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_255_port
                           );
   out_buf_reg_0_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_254_port
                           );
   out_buf_reg_0_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_253_port
                           );
   out_buf_reg_0_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_252_port
                           );
   out_buf_reg_0_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_251_port
                           );
   out_buf_reg_0_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_250_port
                           );
   out_buf_reg_0_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_249_port
                           );
   out_buf_reg_0_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_248_port
                           );
   out_buf_reg_0_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_247_port
                           );
   out_buf_reg_0_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_246_port
                           );
   out_buf_reg_0_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_245_port
                           );
   out_buf_reg_0_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_244_port
                           );
   out_buf_reg_0_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_243_port
                           );
   out_buf_reg_0_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_242_port
                           );
   out_buf_reg_0_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_241_port
                           );
   out_buf_reg_0_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n248, CK => clk, RB => resetn, Q => out_buf_240_port
                           );
   out_buf_reg_4_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_127_port
                           );
   out_buf_reg_4_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_126_port
                           );
   out_buf_reg_4_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_125_port
                           );
   out_buf_reg_4_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_124_port
                           );
   out_buf_reg_4_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_123_port
                           );
   out_buf_reg_4_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_122_port
                           );
   out_buf_reg_4_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_121_port
                           );
   out_buf_reg_4_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_120_port
                           );
   out_buf_reg_4_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_119_port
                           );
   out_buf_reg_4_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_118_port
                           );
   out_buf_reg_4_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_117_port
                           );
   out_buf_reg_4_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_116_port
                           );
   out_buf_reg_4_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_115_port
                           );
   out_buf_reg_4_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_114_port
                           );
   out_buf_reg_4_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_113_port
                           );
   out_buf_reg_4_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB => 
                           n247, CK => clk, RB => resetn, Q => out_buf_112_port
                           );
   out_trigger_reg : DFFRPQ1 port map( D => n240, CK => clk, RB => resetn, Q =>
                           out_trigger);
   read_comp_res_reg : DFERPQ1 port map( D => avs_writedata(2), CEB => n179, CK
                           => clk, RB => resetn, Q => read_comp_res);
   in_counter_reg_0_inst : DFERPQ1 port map( D => n155, CEB => n800, CK => clk,
                           RB => resetn, Q => in_counter_0_port);
   in_counter_reg_2_inst : DFFRPQ1 port map( D => n238, CK => clk, RB => resetn
                           , Q => in_counter_2_port);
   in_counter_reg_1_inst : DFFRPQ1 port map( D => n237, CK => clk, RB => resetn
                           , Q => in_counter_1_port);
   in_busy_reg : DFFRPQ1 port map( D => n239, CK => clk, RB => resetn, Q => 
                           in_busy);
   odd_reg : DFFRPQ1 port map( D => n156, CK => clk, RB => resetn, Q => odd);
   out_busy_reg : DFFRPQ1 port map( D => n234, CK => clk, RB => resetn, Q => 
                           out_busy);
   odd_reg2 : DFFRPQ1 port map( D => n154, CK => clk, RB => resetn, Q => odd1);
   operand_load_reg : DFERPQ1 port map( D => avs_writedata(1), CEB => n179, CK 
                           => clk, RB => resetn, Q => operand_load);
   coeff_load_reg : DFERPQ1 port map( D => avs_writedata(0), CEB => n179, CK =>
                           clk, RB => resetn, Q => coeff_load);
   out_counter_reg_0_inst : DFFRPQ1 port map( D => n236, CK => clk, RB => 
                           resetn, Q => N62);
   out_counter_reg_2_inst : DFFRPQ1 port map( D => n235, CK => clk, RB => 
                           resetn, Q => N64);
   out_counter_reg_1_inst : DFFRPQ1 port map( D => n201, CK => clk, RB => 
                           resetn, Q => N63);
   operand_regs_reg_3_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           operand_regs_159_port);
   operand_regs_reg_5_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_95_port);
   operand_regs_reg_1_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_223_port);
   coeff_memory_reg_0_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB 
                           => n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_31_port);
   coeff_memory_reg_1_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB 
                           => n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_31_port);
   coeff_memory_reg_2_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_31_port);
   coeff_memory_reg_3_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_31_port);
   coeff_memory_reg_4_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_31_port);
   operand_regs_reg_2_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_191_port);
   operand_regs_reg_4_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_127_port);
   operand_regs_reg_6_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_63_port);
   operand_regs_reg_7_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB 
                           => n242, CK => clk, RB => resetn, Q => 
                           operand_regs_31_port);
   operand_regs_reg_0_31_inst : DFERPQ1 port map( D => avs_writedata(31), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_255_port);
   operand_regs_reg_3_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           operand_regs_158_port);
   operand_regs_reg_5_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_94_port);
   operand_regs_reg_3_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           operand_regs_157_port);
   operand_regs_reg_5_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_93_port);
   coeff_memory_reg_0_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB 
                           => n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_30_port);
   coeff_memory_reg_1_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB 
                           => n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_30_port);
   coeff_memory_reg_2_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_30_port);
   coeff_memory_reg_3_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_30_port);
   coeff_memory_reg_4_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_30_port);
   operand_regs_reg_2_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_190_port);
   operand_regs_reg_4_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_126_port);
   operand_regs_reg_6_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_62_port);
   operand_regs_reg_1_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_222_port);
   operand_regs_reg_7_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB 
                           => n242, CK => clk, RB => resetn, Q => 
                           operand_regs_30_port);
   operand_regs_reg_0_30_inst : DFERPQ1 port map( D => avs_writedata(30), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_254_port);
   operand_regs_reg_1_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_221_port);
   operand_regs_reg_3_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           operand_regs_156_port);
   operand_regs_reg_5_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_92_port);
   coeff_memory_reg_0_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB 
                           => n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_29_port);
   coeff_memory_reg_1_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB 
                           => n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_29_port);
   coeff_memory_reg_2_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_29_port);
   coeff_memory_reg_3_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_29_port);
   coeff_memory_reg_4_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_29_port);
   operand_regs_reg_2_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_189_port);
   operand_regs_reg_4_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_125_port);
   operand_regs_reg_6_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_61_port);
   operand_regs_reg_7_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB 
                           => n242, CK => clk, RB => resetn, Q => 
                           operand_regs_29_port);
   operand_regs_reg_0_29_inst : DFERPQ1 port map( D => avs_writedata(29), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_253_port);
   operand_regs_reg_1_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_220_port);
   operand_regs_reg_3_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           operand_regs_155_port);
   operand_regs_reg_5_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_91_port);
   coeff_memory_reg_0_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB 
                           => n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_28_port);
   coeff_memory_reg_1_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB 
                           => n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_28_port);
   coeff_memory_reg_2_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_28_port);
   coeff_memory_reg_3_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_28_port);
   coeff_memory_reg_4_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_28_port);
   operand_regs_reg_2_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_188_port);
   operand_regs_reg_4_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_124_port);
   operand_regs_reg_6_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_60_port);
   operand_regs_reg_7_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB 
                           => n242, CK => clk, RB => resetn, Q => 
                           operand_regs_28_port);
   operand_regs_reg_0_28_inst : DFERPQ1 port map( D => avs_writedata(28), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_252_port);
   avs_readdata_reg_30_inst : DFFSPQ1 port map( D => n203, CK => clk, SB => 
                           resetn, Q => avs_readdata_30_port);
   avs_readdata_reg_28_inst : DFFSPQ1 port map( D => n205, CK => clk, SB => 
                           resetn, Q => avs_readdata_28_port);
   avs_readdata_reg_26_inst : DFFSPQ1 port map( D => n207, CK => clk, SB => 
                           resetn, Q => avs_readdata_26_port);
   avs_readdata_reg_24_inst : DFFSPQ1 port map( D => n209, CK => clk, SB => 
                           resetn, Q => avs_readdata_24_port);
   avs_readdata_reg_22_inst : DFFSPQ1 port map( D => n211, CK => clk, SB => 
                           resetn, Q => avs_readdata_22_port);
   avs_readdata_reg_20_inst : DFFSPQ1 port map( D => n213, CK => clk, SB => 
                           resetn, Q => avs_readdata_20_port);
   avs_readdata_reg_18_inst : DFFSPQ1 port map( D => n215, CK => clk, SB => 
                           resetn, Q => avs_readdata_18_port);
   avs_readdata_reg_16_inst : DFFSPQ1 port map( D => n217, CK => clk, SB => 
                           resetn, Q => avs_readdata_16_port);
   avs_readdata_reg_14_inst : DFFSPQ1 port map( D => n219, CK => clk, SB => 
                           resetn, Q => avs_readdata_14_port);
   avs_readdata_reg_12_inst : DFFSPQ1 port map( D => n221, CK => clk, SB => 
                           resetn, Q => avs_readdata_12_port);
   avs_readdata_reg_10_inst : DFFSPQ1 port map( D => n223, CK => clk, SB => 
                           resetn, Q => avs_readdata_10_port);
   avs_readdata_reg_8_inst : DFFSPQ1 port map( D => n225, CK => clk, SB => 
                           resetn, Q => avs_readdata_8_port);
   avs_readdata_reg_6_inst : DFFSPQ1 port map( D => n227, CK => clk, SB => 
                           resetn, Q => avs_readdata_6_port);
   avs_readdata_reg_4_inst : DFFSPQ1 port map( D => n229, CK => clk, SB => 
                           resetn, Q => avs_readdata_4_port);
   avs_readdata_reg_2_inst : DFFSPQ1 port map( D => n231, CK => clk, SB => 
                           resetn, Q => avs_readdata_2_port);
   avs_readdata_reg_0_inst : DFFSPQ1 port map( D => n233, CK => clk, SB => 
                           resetn, Q => avs_readdata_0_port);
   operand_regs_reg_3_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           operand_regs_154_port);
   operand_regs_reg_5_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_90_port);
   operand_regs_reg_1_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_219_port);
   avs_readdata_reg_31_inst : DFFRPQ1 port map( D => n202, CK => clk, RB => 
                           resetn, Q => avs_readdata_31_port);
   avs_readdata_reg_29_inst : DFFRPQ1 port map( D => n204, CK => clk, RB => 
                           resetn, Q => avs_readdata_29_port);
   avs_readdata_reg_27_inst : DFFRPQ1 port map( D => n206, CK => clk, RB => 
                           resetn, Q => avs_readdata_27_port);
   avs_readdata_reg_25_inst : DFFRPQ1 port map( D => n208, CK => clk, RB => 
                           resetn, Q => avs_readdata_25_port);
   avs_readdata_reg_23_inst : DFFRPQ1 port map( D => n210, CK => clk, RB => 
                           resetn, Q => avs_readdata_23_port);
   avs_readdata_reg_21_inst : DFFRPQ1 port map( D => n212, CK => clk, RB => 
                           resetn, Q => avs_readdata_21_port);
   avs_readdata_reg_19_inst : DFFRPQ1 port map( D => n214, CK => clk, RB => 
                           resetn, Q => avs_readdata_19_port);
   avs_readdata_reg_17_inst : DFFRPQ1 port map( D => n216, CK => clk, RB => 
                           resetn, Q => avs_readdata_17_port);
   avs_readdata_reg_15_inst : DFFRPQ1 port map( D => n218, CK => clk, RB => 
                           resetn, Q => avs_readdata_15_port);
   avs_readdata_reg_13_inst : DFFRPQ1 port map( D => n220, CK => clk, RB => 
                           resetn, Q => avs_readdata_13_port);
   avs_readdata_reg_11_inst : DFFRPQ1 port map( D => n222, CK => clk, RB => 
                           resetn, Q => avs_readdata_11_port);
   avs_readdata_reg_9_inst : DFFRPQ1 port map( D => n224, CK => clk, RB => 
                           resetn, Q => avs_readdata_9_port);
   avs_readdata_reg_7_inst : DFFRPQ1 port map( D => n226, CK => clk, RB => 
                           resetn, Q => avs_readdata_7_port);
   avs_readdata_reg_5_inst : DFFRPQ1 port map( D => n228, CK => clk, RB => 
                           resetn, Q => avs_readdata_5_port);
   avs_readdata_reg_3_inst : DFFRPQ1 port map( D => n230, CK => clk, RB => 
                           resetn, Q => avs_readdata_3_port);
   avs_readdata_reg_1_inst : DFFRPQ1 port map( D => n232, CK => clk, RB => 
                           resetn, Q => avs_readdata_1_port);
   stop_sim_reg : DFFRPQ1 port map( D => n157, CK => clk, RB => resetn, Q => 
                           stop_sim_port);
   operand_regs_reg_1_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_218_port);
   coeff_memory_reg_0_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB 
                           => n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_27_port);
   coeff_memory_reg_1_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB 
                           => n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_27_port);
   coeff_memory_reg_2_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_27_port);
   coeff_memory_reg_3_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_27_port);
   coeff_memory_reg_4_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_27_port);
   operand_regs_reg_2_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_187_port);
   operand_regs_reg_4_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_123_port);
   operand_regs_reg_6_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_59_port);
   operand_regs_reg_7_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB 
                           => n242, CK => clk, RB => resetn, Q => 
                           operand_regs_27_port);
   operand_regs_reg_0_27_inst : DFERPQ1 port map( D => avs_writedata(27), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_251_port);
   operand_regs_reg_3_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           operand_regs_153_port);
   operand_regs_reg_5_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_89_port);
   coeff_memory_reg_0_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB 
                           => n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_26_port);
   coeff_memory_reg_1_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB 
                           => n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_26_port);
   coeff_memory_reg_2_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_26_port);
   coeff_memory_reg_3_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_26_port);
   coeff_memory_reg_4_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_26_port);
   operand_regs_reg_2_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_186_port);
   operand_regs_reg_4_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_122_port);
   operand_regs_reg_6_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_58_port);
   operand_regs_reg_7_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB 
                           => n242, CK => clk, RB => resetn, Q => 
                           operand_regs_26_port);
   operand_regs_reg_0_26_inst : DFERPQ1 port map( D => avs_writedata(26), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_250_port);
   operand_regs_reg_1_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_217_port);
   operand_regs_reg_3_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           operand_regs_152_port);
   operand_regs_reg_5_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_88_port);
   operand_regs_reg_1_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_216_port);
   coeff_memory_reg_0_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB 
                           => n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_25_port);
   coeff_memory_reg_1_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB 
                           => n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_25_port);
   coeff_memory_reg_2_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_25_port);
   coeff_memory_reg_3_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_25_port);
   coeff_memory_reg_4_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_25_port);
   operand_regs_reg_2_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_185_port);
   operand_regs_reg_4_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_121_port);
   operand_regs_reg_6_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_57_port);
   operand_regs_reg_3_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           operand_regs_151_port);
   operand_regs_reg_5_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_87_port);
   operand_regs_reg_7_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB 
                           => n242, CK => clk, RB => resetn, Q => 
                           operand_regs_25_port);
   operand_regs_reg_0_25_inst : DFERPQ1 port map( D => avs_writedata(25), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_249_port);
   operand_regs_reg_1_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_215_port);
   coeff_memory_reg_0_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB 
                           => n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_24_port);
   coeff_memory_reg_1_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB 
                           => n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_24_port);
   coeff_memory_reg_2_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_24_port);
   coeff_memory_reg_3_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_24_port);
   coeff_memory_reg_4_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_24_port);
   operand_regs_reg_2_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_184_port);
   operand_regs_reg_4_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_120_port);
   operand_regs_reg_6_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_56_port);
   operand_regs_reg_7_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB 
                           => n242, CK => clk, RB => resetn, Q => 
                           operand_regs_24_port);
   operand_regs_reg_0_24_inst : DFERPQ1 port map( D => avs_writedata(24), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_248_port);
   coeff_memory_reg_0_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB 
                           => n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_23_port);
   coeff_memory_reg_1_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB 
                           => n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_23_port);
   coeff_memory_reg_2_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_23_port);
   coeff_memory_reg_3_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_23_port);
   coeff_memory_reg_4_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_23_port);
   operand_regs_reg_2_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_183_port);
   operand_regs_reg_4_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_119_port);
   operand_regs_reg_6_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_55_port);
   operand_regs_reg_7_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB 
                           => n242, CK => clk, RB => resetn, Q => 
                           operand_regs_23_port);
   operand_regs_reg_0_23_inst : DFERPQ1 port map( D => avs_writedata(23), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_247_port);
   operand_regs_reg_3_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           operand_regs_150_port);
   operand_regs_reg_5_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_86_port);
   operand_regs_reg_3_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           operand_regs_149_port);
   operand_regs_reg_5_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_85_port);
   coeff_memory_reg_0_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB 
                           => n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_22_port);
   coeff_memory_reg_1_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB 
                           => n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_22_port);
   coeff_memory_reg_2_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_22_port);
   coeff_memory_reg_3_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_22_port);
   coeff_memory_reg_4_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_22_port);
   operand_regs_reg_2_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_182_port);
   operand_regs_reg_4_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_118_port);
   operand_regs_reg_6_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_54_port);
   operand_regs_reg_7_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB 
                           => n242, CK => clk, RB => resetn, Q => 
                           operand_regs_22_port);
   operand_regs_reg_0_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_246_port);
   operand_regs_reg_1_22_inst : DFERPQ1 port map( D => avs_writedata(22), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_214_port);
   operand_regs_reg_3_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           operand_regs_148_port);
   operand_regs_reg_5_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_84_port);
   coeff_memory_reg_0_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB 
                           => n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_21_port);
   coeff_memory_reg_1_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB 
                           => n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_21_port);
   coeff_memory_reg_2_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_21_port);
   coeff_memory_reg_3_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_21_port);
   coeff_memory_reg_4_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_21_port);
   operand_regs_reg_2_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_181_port);
   operand_regs_reg_4_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_117_port);
   operand_regs_reg_6_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_53_port);
   operand_regs_reg_1_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_213_port);
   operand_regs_reg_3_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           operand_regs_147_port);
   operand_regs_reg_5_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_83_port);
   operand_regs_reg_7_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB 
                           => n242, CK => clk, RB => resetn, Q => 
                           operand_regs_21_port);
   operand_regs_reg_0_21_inst : DFERPQ1 port map( D => avs_writedata(21), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_245_port);
   operand_regs_reg_3_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           operand_regs_144_port);
   operand_regs_reg_5_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_80_port);
   operand_regs_reg_3_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           operand_regs_146_port);
   operand_regs_reg_5_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_82_port);
   operand_regs_reg_3_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           operand_regs_143_port);
   operand_regs_reg_5_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_79_port);
   operand_regs_reg_3_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           operand_regs_139_port);
   operand_regs_reg_5_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_75_port);
   operand_regs_reg_3_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           operand_regs_145_port);
   operand_regs_reg_5_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_81_port);
   operand_regs_reg_3_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           operand_regs_142_port);
   operand_regs_reg_5_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_78_port);
   operand_regs_reg_3_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           operand_regs_141_port);
   operand_regs_reg_5_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_77_port);
   operand_regs_reg_3_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           operand_regs_140_port);
   operand_regs_reg_5_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_76_port);
   operand_regs_reg_1_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_212_port);
   coeff_memory_reg_0_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB 
                           => n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_20_port);
   coeff_memory_reg_1_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB 
                           => n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_20_port);
   coeff_memory_reg_2_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_20_port);
   coeff_memory_reg_3_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_20_port);
   coeff_memory_reg_4_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_20_port);
   operand_regs_reg_2_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_180_port);
   operand_regs_reg_4_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_116_port);
   operand_regs_reg_6_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_52_port);
   operand_regs_reg_1_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_211_port);
   operand_regs_reg_7_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB 
                           => n242, CK => clk, RB => resetn, Q => 
                           operand_regs_20_port);
   operand_regs_reg_0_20_inst : DFERPQ1 port map( D => avs_writedata(20), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_244_port);
   operand_regs_reg_1_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_208_port);
   operand_regs_reg_3_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB 
                           => n261, CK => clk, RB => resetn, Q => 
                           operand_regs_138_port);
   operand_regs_reg_5_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB 
                           => n260, CK => clk, RB => resetn, Q => 
                           operand_regs_74_port);
   coeff_memory_reg_3_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_0_port);
   coeff_memory_reg_4_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_0_port);
   operand_regs_reg_1_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_210_port);
   coeff_memory_reg_0_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_0_port);
   operand_regs_reg_6_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_32_port);
   coeff_memory_reg_0_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB 
                           => n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_19_port);
   coeff_memory_reg_1_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB 
                           => n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_19_port);
   coeff_memory_reg_2_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_19_port);
   coeff_memory_reg_3_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_19_port);
   coeff_memory_reg_4_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_19_port);
   coeff_memory_reg_1_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_0_port);
   coeff_memory_reg_2_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_0_port);
   operand_regs_reg_2_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_179_port);
   operand_regs_reg_4_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_115_port);
   operand_regs_reg_6_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_51_port);
   operand_regs_reg_2_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_160_port);
   operand_regs_reg_4_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_96_port);
   operand_regs_reg_1_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_207_port);
   operand_regs_reg_7_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB 
                           => n242, CK => clk, RB => resetn, Q => 
                           operand_regs_19_port);
   operand_regs_reg_1_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_209_port);
   operand_regs_reg_0_19_inst : DFERPQ1 port map( D => avs_writedata(19), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_243_port);
   coeff_memory_reg_0_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB 
                           => n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_18_port);
   coeff_memory_reg_1_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB 
                           => n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_18_port);
   coeff_memory_reg_2_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_18_port);
   coeff_memory_reg_3_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_18_port);
   coeff_memory_reg_4_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_18_port);
   operand_regs_reg_2_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_178_port);
   operand_regs_reg_4_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_114_port);
   operand_regs_reg_6_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_50_port);
   operand_regs_reg_3_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_137_port);
   operand_regs_reg_5_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_73_port);
   operand_regs_reg_7_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB 
                           => n242, CK => clk, RB => resetn, Q => 
                           operand_regs_18_port);
   operand_regs_reg_0_18_inst : DFERPQ1 port map( D => avs_writedata(18), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_242_port);
   operand_regs_reg_3_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_132_port);
   operand_regs_reg_5_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_68_port);
   operand_regs_reg_3_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_131_port);
   operand_regs_reg_5_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_67_port);
   operand_regs_reg_3_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_128_port);
   operand_regs_reg_5_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_64_port);
   coeff_memory_reg_0_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB 
                           => n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_10_port);
   coeff_memory_reg_1_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB 
                           => n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_10_port);
   coeff_memory_reg_2_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_10_port);
   coeff_memory_reg_3_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_10_port);
   coeff_memory_reg_4_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_10_port);
   operand_regs_reg_2_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_170_port);
   operand_regs_reg_4_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_106_port);
   operand_regs_reg_6_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_42_port);
   operand_regs_reg_0_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_234_port);
   coeff_memory_reg_0_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB 
                           => n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_17_port);
   coeff_memory_reg_1_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB 
                           => n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_17_port);
   coeff_memory_reg_2_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_17_port);
   coeff_memory_reg_3_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_17_port);
   coeff_memory_reg_4_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_17_port);
   operand_regs_reg_2_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_177_port);
   operand_regs_reg_4_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_113_port);
   operand_regs_reg_6_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_49_port);
   operand_regs_reg_3_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_133_port);
   operand_regs_reg_5_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_69_port);
   operand_regs_reg_7_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB 
                           => n242, CK => clk, RB => resetn, Q => 
                           operand_regs_17_port);
   operand_regs_reg_3_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_129_port);
   operand_regs_reg_5_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_65_port);
   operand_regs_reg_0_17_inst : DFERPQ1 port map( D => avs_writedata(17), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_241_port);
   coeff_memory_reg_0_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB 
                           => n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_16_port);
   coeff_memory_reg_1_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB 
                           => n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_16_port);
   coeff_memory_reg_2_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_16_port);
   coeff_memory_reg_3_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_16_port);
   coeff_memory_reg_4_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_16_port);
   operand_regs_reg_2_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_176_port);
   operand_regs_reg_4_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_112_port);
   operand_regs_reg_6_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_48_port);
   operand_regs_reg_3_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_130_port);
   operand_regs_reg_5_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_66_port);
   coeff_memory_reg_0_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB 
                           => n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_14_port);
   coeff_memory_reg_1_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB 
                           => n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_14_port);
   coeff_memory_reg_2_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_14_port);
   coeff_memory_reg_3_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_14_port);
   coeff_memory_reg_4_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_14_port);
   operand_regs_reg_7_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB 
                           => n242, CK => clk, RB => resetn, Q => 
                           operand_regs_16_port);
   operand_regs_reg_3_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_136_port);
   operand_regs_reg_5_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_72_port);
   operand_regs_reg_0_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_224_port);
   operand_regs_reg_0_16_inst : DFERPQ1 port map( D => avs_writedata(16), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_240_port);
   operand_regs_reg_2_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_174_port);
   operand_regs_reg_4_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_110_port);
   operand_regs_reg_6_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_46_port);
   operand_regs_reg_3_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_135_port);
   operand_regs_reg_5_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_71_port);
   operand_regs_reg_3_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => 
                           n261, CK => clk, RB => resetn, Q => 
                           operand_regs_134_port);
   operand_regs_reg_5_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => 
                           n260, CK => clk, RB => resetn, Q => 
                           operand_regs_70_port);
   operand_regs_reg_0_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_238_port);
   operand_regs_reg_1_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_203_port);
   coeff_memory_reg_0_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB 
                           => n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_13_port);
   coeff_memory_reg_1_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB 
                           => n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_13_port);
   coeff_memory_reg_2_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_13_port);
   coeff_memory_reg_3_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_13_port);
   coeff_memory_reg_4_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_13_port);
   operand_regs_reg_7_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB 
                           => n242, CK => clk, RB => resetn, Q => 
                           operand_regs_14_port);
   operand_regs_reg_2_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_173_port);
   operand_regs_reg_4_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_109_port);
   operand_regs_reg_6_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_45_port);
   coeff_memory_reg_0_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB 
                           => n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_15_port);
   coeff_memory_reg_1_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB 
                           => n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_15_port);
   coeff_memory_reg_2_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_15_port);
   coeff_memory_reg_3_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_15_port);
   coeff_memory_reg_4_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_15_port);
   operand_regs_reg_2_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_175_port);
   operand_regs_reg_4_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_111_port);
   operand_regs_reg_6_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_47_port);
   coeff_memory_reg_0_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB 
                           => n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_12_port);
   coeff_memory_reg_1_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB 
                           => n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_12_port);
   coeff_memory_reg_2_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_12_port);
   coeff_memory_reg_3_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_12_port);
   coeff_memory_reg_4_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_12_port);
   operand_regs_reg_1_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_204_port);
   operand_regs_reg_7_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB 
                           => n242, CK => clk, RB => resetn, Q => 
                           operand_regs_13_port);
   operand_regs_reg_1_14_inst : DFERPQ1 port map( D => avs_writedata(14), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_206_port);
   operand_regs_reg_0_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_237_port);
   operand_regs_reg_2_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_172_port);
   operand_regs_reg_4_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_108_port);
   operand_regs_reg_6_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_44_port);
   operand_regs_reg_1_13_inst : DFERPQ1 port map( D => avs_writedata(13), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_205_port);
   operand_regs_reg_7_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB 
                           => n242, CK => clk, RB => resetn, Q => 
                           operand_regs_15_port);
   coeff_memory_reg_0_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_9_port);
   coeff_memory_reg_1_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_9_port);
   coeff_memory_reg_2_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_9_port);
   coeff_memory_reg_3_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_9_port);
   coeff_memory_reg_4_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_9_port);
   operand_regs_reg_2_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_169_port);
   operand_regs_reg_4_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_105_port);
   operand_regs_reg_6_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_41_port);
   operand_regs_reg_0_15_inst : DFERPQ1 port map( D => avs_writedata(15), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_239_port);
   operand_regs_reg_7_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_0_port);
   operand_regs_reg_7_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB 
                           => n242, CK => clk, RB => resetn, Q => 
                           operand_regs_12_port);
   operand_regs_reg_0_12_inst : DFERPQ1 port map( D => avs_writedata(12), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_236_port);
   operand_regs_reg_0_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_233_port);
   operand_regs_reg_7_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB 
                           => n242, CK => clk, RB => resetn, Q => 
                           operand_regs_10_port);
   operand_regs_reg_1_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_196_port);
   operand_regs_reg_1_0_inst : DFERPQ1 port map( D => avs_writedata(0), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_192_port);
   coeff_memory_reg_0_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB 
                           => n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_11_port);
   coeff_memory_reg_1_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB 
                           => n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_11_port);
   coeff_memory_reg_2_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB 
                           => n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_11_port);
   coeff_memory_reg_3_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB 
                           => n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_11_port);
   coeff_memory_reg_4_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB 
                           => n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_11_port);
   operand_regs_reg_1_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_195_port);
   operand_regs_reg_2_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB 
                           => n258, CK => clk, RB => resetn, Q => 
                           operand_regs_171_port);
   operand_regs_reg_4_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB 
                           => n257, CK => clk, RB => resetn, Q => 
                           operand_regs_107_port);
   operand_regs_reg_6_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB 
                           => n256, CK => clk, RB => resetn, Q => 
                           operand_regs_43_port);
   operand_regs_reg_1_10_inst : DFERPQ1 port map( D => avs_writedata(10), CEB 
                           => n259, CK => clk, RB => resetn, Q => 
                           operand_regs_202_port);
   operand_regs_reg_7_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB 
                           => n242, CK => clk, RB => resetn, Q => 
                           operand_regs_11_port);
   operand_regs_reg_0_11_inst : DFERPQ1 port map( D => avs_writedata(11), CEB 
                           => n255, CK => clk, RB => resetn, Q => 
                           operand_regs_235_port);
   operand_regs_reg_1_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_194_port);
   operand_regs_reg_1_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_193_port);
   operand_regs_reg_7_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_9_port);
   operand_regs_reg_1_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_197_port);
   operand_regs_reg_1_9_inst : DFERPQ1 port map( D => avs_writedata(9), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_201_port);
   operand_regs_reg_1_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_200_port);
   operand_regs_reg_1_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_199_port);
   operand_regs_reg_1_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => 
                           n259, CK => clk, RB => resetn, Q => 
                           operand_regs_198_port);
   coeff_memory_reg_0_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_8_port);
   coeff_memory_reg_1_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_8_port);
   coeff_memory_reg_2_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_8_port);
   coeff_memory_reg_3_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_8_port);
   coeff_memory_reg_4_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_8_port);
   operand_regs_reg_2_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_168_port);
   operand_regs_reg_4_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_104_port);
   operand_regs_reg_6_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_40_port);
   coeff_memory_reg_0_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_4_port);
   coeff_memory_reg_1_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_4_port);
   coeff_memory_reg_2_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_4_port);
   coeff_memory_reg_3_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_4_port);
   coeff_memory_reg_4_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_4_port);
   operand_regs_reg_2_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_164_port);
   operand_regs_reg_4_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_100_port);
   operand_regs_reg_6_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_36_port);
   operand_regs_reg_7_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_8_port);
   operand_regs_reg_7_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_4_port);
   operand_regs_reg_0_8_inst : DFERPQ1 port map( D => avs_writedata(8), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_232_port);
   operand_regs_reg_0_4_inst : DFERPQ1 port map( D => avs_writedata(4), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_228_port);
   coeff_memory_reg_0_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_6_port);
   coeff_memory_reg_1_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_6_port);
   coeff_memory_reg_2_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_6_port);
   coeff_memory_reg_3_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_6_port);
   coeff_memory_reg_4_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_6_port);
   operand_regs_reg_2_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_166_port);
   operand_regs_reg_4_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_102_port);
   operand_regs_reg_6_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_38_port);
   operand_regs_reg_7_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_6_port);
   operand_regs_reg_0_6_inst : DFERPQ1 port map( D => avs_writedata(6), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_230_port);
   coeff_memory_reg_0_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_7_port);
   coeff_memory_reg_1_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_7_port);
   coeff_memory_reg_2_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_7_port);
   coeff_memory_reg_3_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_7_port);
   coeff_memory_reg_4_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_7_port);
   operand_regs_reg_2_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_167_port);
   operand_regs_reg_4_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_103_port);
   operand_regs_reg_6_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_39_port);
   coeff_memory_reg_0_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_3_port);
   coeff_memory_reg_1_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_3_port);
   coeff_memory_reg_2_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_3_port);
   coeff_memory_reg_3_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_3_port);
   coeff_memory_reg_4_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_3_port);
   operand_regs_reg_2_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_163_port);
   operand_regs_reg_4_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_99_port);
   operand_regs_reg_6_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_35_port);
   coeff_memory_reg_0_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_2_port);
   coeff_memory_reg_1_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_2_port);
   coeff_memory_reg_2_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_2_port);
   coeff_memory_reg_3_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_2_port);
   coeff_memory_reg_4_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_2_port);
   operand_regs_reg_2_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_162_port);
   operand_regs_reg_4_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_98_port);
   operand_regs_reg_6_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_34_port);
   operand_regs_reg_7_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_7_port);
   operand_regs_reg_7_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_3_port);
   operand_regs_reg_0_7_inst : DFERPQ1 port map( D => avs_writedata(7), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_231_port);
   operand_regs_reg_0_3_inst : DFERPQ1 port map( D => avs_writedata(3), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_227_port);
   operand_regs_reg_7_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_2_port);
   coeff_memory_reg_0_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_5_port);
   coeff_memory_reg_1_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_5_port);
   coeff_memory_reg_2_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_5_port);
   coeff_memory_reg_3_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_5_port);
   coeff_memory_reg_4_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_5_port);
   operand_regs_reg_2_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_165_port);
   operand_regs_reg_4_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_101_port);
   operand_regs_reg_6_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_37_port);
   operand_regs_reg_0_2_inst : DFERPQ1 port map( D => avs_writedata(2), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_226_port);
   operand_regs_reg_7_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_5_port);
   operand_regs_reg_0_5_inst : DFERPQ1 port map( D => avs_writedata(5), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_229_port);
   coeff_memory_reg_0_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => 
                           n267, CK => clk, RB => resetn, Q => 
                           coeff_memory_0_1_port);
   coeff_memory_reg_1_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => 
                           n266, CK => clk, RB => resetn, Q => 
                           coeff_memory_1_1_port);
   coeff_memory_reg_2_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => 
                           n264, CK => clk, RB => resetn, Q => 
                           coeff_memory_2_1_port);
   coeff_memory_reg_3_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => 
                           n263, CK => clk, RB => resetn, Q => 
                           coeff_memory_3_1_port);
   coeff_memory_reg_4_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => 
                           n265, CK => clk, RB => resetn, Q => 
                           coeff_memory_4_1_port);
   operand_regs_reg_2_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => 
                           n258, CK => clk, RB => resetn, Q => 
                           operand_regs_161_port);
   operand_regs_reg_4_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => 
                           n257, CK => clk, RB => resetn, Q => 
                           operand_regs_97_port);
   operand_regs_reg_6_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => 
                           n256, CK => clk, RB => resetn, Q => 
                           operand_regs_33_port);
   operand_regs_reg_7_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => 
                           n242, CK => clk, RB => resetn, Q => 
                           operand_regs_1_port);
   operand_regs_reg_0_1_inst : DFERPQ1 port map( D => avs_writedata(1), CEB => 
                           n255, CK => clk, RB => resetn, Q => 
                           operand_regs_225_port);
   filt_mult_inputs_reg : DFERPQ1 port map( D => avs_writedata(0), CEB => n178,
                           CK => clk, RB => resetn, Q => filt_mult_inputs);
   siso_req_reg : DFERPQ1 port map( D => n806, CEB => n161, CK => clk, RB => 
                           resetn, Q => siso_req);
   siso_data_out_reg_0_inst : DFERPQ1 port map( D => N2888, CEB => n811, CK => 
                           clk, RB => resetn, Q => siso_data_out(0));
   siso_data_out_reg_15_inst : DFERPQ1 port map( D => N2903, CEB => n811, CK =>
                           clk, RB => resetn, Q => siso_data_out(15));
   siso_data_out_reg_14_inst : DFERPQ1 port map( D => N2902, CEB => n811, CK =>
                           clk, RB => resetn, Q => siso_data_out(14));
   siso_data_out_reg_13_inst : DFERPQ1 port map( D => N2901, CEB => n811, CK =>
                           clk, RB => resetn, Q => siso_data_out(13));
   siso_data_out_reg_12_inst : DFERPQ1 port map( D => N2900, CEB => n811, CK =>
                           clk, RB => resetn, Q => siso_data_out(12));
   siso_data_out_reg_11_inst : DFERPQ1 port map( D => N2899, CEB => n811, CK =>
                           clk, RB => resetn, Q => siso_data_out(11));
   siso_data_out_reg_10_inst : DFERPQ1 port map( D => N2898, CEB => n811, CK =>
                           clk, RB => resetn, Q => siso_data_out(10));
   siso_data_out_reg_9_inst : DFERPQ1 port map( D => N2897, CEB => n811, CK => 
                           clk, RB => resetn, Q => siso_data_out(9));
   siso_data_out_reg_8_inst : DFERPQ1 port map( D => N2896, CEB => n811, CK => 
                           clk, RB => resetn, Q => siso_data_out(8));
   siso_data_out_reg_7_inst : DFERPQ1 port map( D => N2895, CEB => n811, CK => 
                           clk, RB => resetn, Q => siso_data_out(7));
   siso_data_out_reg_6_inst : DFERPQ1 port map( D => N2894, CEB => n811, CK => 
                           clk, RB => resetn, Q => siso_data_out(6));
   siso_data_out_reg_5_inst : DFERPQ1 port map( D => N2893, CEB => n811, CK => 
                           clk, RB => resetn, Q => siso_data_out(5));
   siso_data_out_reg_4_inst : DFERPQ1 port map( D => N2892, CEB => n811, CK => 
                           clk, RB => resetn, Q => siso_data_out(4));
   siso_data_out_reg_3_inst : DFERPQ1 port map( D => N2891, CEB => n811, CK => 
                           clk, RB => resetn, Q => siso_data_out(3));
   siso_data_out_reg_2_inst : DFERPQ1 port map( D => N2890, CEB => n811, CK => 
                           clk, RB => resetn, Q => siso_data_out(2));
   siso_data_out_reg_1_inst : DFERPQ1 port map( D => N2889, CEB => n811, CK => 
                           clk, RB => resetn, Q => siso_data_out(1));
   siso_ready_reg : DFFRPQ1 port map( D => out_busy, CK => clk, RB => resetn, Q
                           => siso_ready);
   U642 : NAN3D1 port map( A1 => n309, A2 => avs_addr(0), A3 => n254, Z => n242
                           );
   U643 : AND2D1 port map( A1 => n313, A2 => avs_addr(0), Z => n243);
   U644 : AND2D1 port map( A1 => n561, A2 => N62, Z => n244);
   U645 : AND2D1 port map( A1 => n563, A2 => N62, Z => n245);
   U646 : NAN3D1 port map( A1 => n309, A2 => avs_addr(0), A3 => n110, Z => n246
                           );
   U647 : NAN2D1 port map( A1 => n110, A2 => n276, Z => n247);
   U648 : NAN2D1 port map( A1 => n110, A2 => n275, Z => n248);
   U649 : NAN2D1 port map( A1 => n110, A2 => n308, Z => n249);
   U650 : NAN2D1 port map( A1 => n110, A2 => n304, Z => n250);
   U651 : NAN2D1 port map( A1 => n110, A2 => n277, Z => n251);
   U652 : NAN2D1 port map( A1 => n110, A2 => n307, Z => n252);
   U653 : NAN2D1 port map( A1 => n110, A2 => n306, Z => n253);
   U654 : AND3D1 port map( A1 => operand_load, A2 => n104, A3 => n729, Z => 
                           n254);
   U655 : NAN2D1 port map( A1 => n275, A2 => n254, Z => n255);
   U656 : NAN2D1 port map( A1 => n277, A2 => n254, Z => n256);
   U657 : NAN2D1 port map( A1 => n276, A2 => n254, Z => n257);
   U658 : NAN2D1 port map( A1 => n307, A2 => n254, Z => n258);
   U659 : NAN2D1 port map( A1 => n308, A2 => n254, Z => n259);
   U660 : NAN2D1 port map( A1 => n304, A2 => n254, Z => n260);
   U661 : NAN2D1 port map( A1 => n306, A2 => n254, Z => n261);
   U662 : AND2D1 port map( A1 => n314, A2 => avs_addr(0), Z => n262);
   U663 : NAN2D1 port map( A1 => n306, A2 => n301, Z => n263);
   U664 : NAN2D1 port map( A1 => n307, A2 => n301, Z => n264);
   U665 : NAN2D1 port map( A1 => n276, A2 => n301, Z => n265);
   U666 : NAN2D1 port map( A1 => n308, A2 => n301, Z => n266);
   U667 : NAN2D1 port map( A1 => n275, A2 => n301, Z => n267);
   U668 : AND3D1 port map( A1 => N66, A2 => n300, A3 => read_comp_res, Z => 
                           n268);
   U669 : AND2D1 port map( A1 => n560, A2 => N62, Z => n269);
   U670 : AND2D1 port map( A1 => n562, A2 => N62, Z => n270);
   U671 : MUX2D1 port map( A0 => operand_regs_12_port, A1 => 
                           operand_regs_204_port, SL => n720, Z => n271);
   U672 : MUX2DL port map( A0 => operand_regs_13_port, A1 => 
                           operand_regs_205_port, SL => n719, Z => n272);
   U673 : MUX2DL port map( A0 => operand_regs_14_port, A1 => 
                           operand_regs_206_port, SL => n720, Z => n273);
   U674 : MUX2D1 port map( A0 => operand_regs_11_port, A1 => 
                           operand_regs_203_port, SL => n719, Z => n274);
   U675 : INVD1 port map( A => n724, Z => n710);
   U676 : INVD1 port map( A => n724, Z => n712);
   U677 : INVD1 port map( A => n724, Z => n711);
   U678 : INVD1 port map( A => n725, Z => n709);
   U679 : INVD1 port map( A => n725, Z => n707);
   U680 : INVD1 port map( A => n725, Z => n708);
   U681 : INVD1 port map( A => n726, Z => n706);
   U682 : INVD1 port map( A => n96, Z => n798);
   U683 : INVD1 port map( A => n702, Z => n724);
   U684 : INVD1 port map( A => n722, Z => n716);
   U685 : INVD1 port map( A => n723, Z => n714);
   U686 : INVD1 port map( A => n722, Z => n718);
   U687 : INVD1 port map( A => n723, Z => n715);
   U688 : INVD1 port map( A => n722, Z => n717);
   U689 : INVD1 port map( A => n702, Z => n725);
   U690 : INVD1 port map( A => n721, Z => n720);
   U691 : INVD1 port map( A => n721, Z => n719);
   U692 : INVD1 port map( A => n723, Z => n713);
   U693 : INVD1 port map( A => n702, Z => n726);
   U694 : INVD1 port map( A => n703, Z => n727);
   U695 : INVD1 port map( A => n703, Z => n728);
   U696 : INVD1 port map( A => n553, Z => n554);
   U697 : INVD1 port map( A => n558, Z => n559);
   U698 : INVD1 port map( A => n555, Z => n557);
   U699 : INVD1 port map( A => n555, Z => n556);
   U700 : INVD1 port map( A => n548, Z => n549);
   U701 : INVD1 port map( A => n548, Z => n550);
   U702 : INVD1 port map( A => n551, Z => n552);
   U703 : NAN2D1 port map( A1 => n275, A2 => n795, Z => n96);
   U704 : INVD1 port map( A => n74, Z => n797);
   U705 : NAN2D1 port map( A1 => n118, A2 => n807, Z => n176);
   U706 : NAN2D1 port map( A1 => n805, A2 => n118, Z => n174);
   U707 : INVD1 port map( A => n704, Z => n702);
   U708 : INVD1 port map( A => n701, Z => n722);
   U709 : INVD1 port map( A => n701, Z => n723);
   U710 : INVD1 port map( A => n701, Z => n721);
   U711 : INVD1 port map( A => n704, Z => n703);
   U712 : INVD1 port map( A => n300, Z => n700);
   U713 : INVD1 port map( A => n541, Z => n553);
   U714 : INVD1 port map( A => n543, Z => n558);
   U715 : INVD1 port map( A => n542, Z => n555);
   U716 : INVD1 port map( A => n699, Z => n698);
   U717 : INVD1 port map( A => n538, Z => n548);
   U718 : INVD1 port map( A => n539, Z => n551);
   U719 : OAI211D1 port map( A1 => n6300, A2 => n6400, B => n300, C => n65, Z 
                           => n14);
   U720 : NOR2D1 port map( A1 => n306, A2 => n307, Z => n6300);
   U721 : NOR3D1 port map( A1 => n797, A2 => N66, A3 => n798, Z => n65);
   U722 : INVD1 port map( A => n6400, Z => n795);
   U723 : NAN2D1 port map( A1 => n308, A2 => n795, Z => n74);
   U724 : AND3D1 port map( A1 => n796, A2 => n547, A3 => n762, Z => n275);
   U725 : AND2D1 port map( A1 => n111, A2 => n762, Z => n276);
   U726 : AND2D1 port map( A1 => n309, A2 => n762, Z => n277);
   U727 : NOR3D1 port map( A1 => n813, A2 => n810, A3 => n696, Z => n78);
   U728 : INVD1 port map( A => n81, Z => n801);
   U729 : INVD1 port map( A => n697, Z => n812);
   U730 : NOR2D1 port map( A1 => n809, A2 => n803, Z => n118);
   U731 : INVD1 port map( A => n88, Z => n807);
   U732 : NOR2D1 port map( A1 => n800, A2 => n91, Z => n89);
   U733 : INVD1 port map( A => n84, Z => n800);
   U734 : INVD1 port map( A => n155, Z => n804);
   U735 : NAN2D1 port map( A1 => n119, A2 => n115, Z => n171);
   U736 : NAN2D1 port map( A1 => n119, A2 => n101, Z => n162);
   U737 : NAN2D1 port map( A1 => n119, A2 => n118, Z => n170);
   U738 : NAN2D1 port map( A1 => n120, A2 => n119, Z => n163);
   U739 : NAN2D1 port map( A1 => n87, A2 => n84, Z => n86);
   U740 : NAN2D1 port map( A1 => n805, A2 => n101, Z => n166);
   U741 : INVD1 port map( A => n85, Z => n805);
   U742 : NAN2D1 port map( A1 => n120, A2 => n805, Z => n167);
   U743 : NAN2D1 port map( A1 => n805, A2 => n115, Z => n175);
   U744 : NAN2D1 port map( A1 => n87, A2 => n101, Z => n164);
   U745 : NAN2D1 port map( A1 => n115, A2 => n87, Z => n173);
   U746 : NAN2D1 port map( A1 => n120, A2 => n87, Z => n165);
   U747 : NAN2D1 port map( A1 => n118, A2 => n87, Z => n172);
   U748 : NAN2D1 port map( A1 => n807, A2 => n101, Z => n168);
   U749 : NAN2D1 port map( A1 => n115, A2 => n807, Z => n177);
   U750 : NAN2D1 port map( A1 => n120, A2 => n807, Z => n169);
   U751 : MUX2DL port map( A0 => operand_regs_33_port, A1 => 
                           coeff_memory_3_1_port, SL => n712, Z => N3010);
   U752 : MUX2DL port map( A0 => operand_regs_97_port, A1 => 
                           coeff_memory_2_1_port, SL => n710, Z => N2978);
   U753 : INVD1 port map( A => filt_mult_inputs, Z => n704);
   U754 : MUX2DL port map( A0 => operand_regs_1_port, A1 => 
                           coeff_memory_4_1_port, SL => n714, Z => N3042);
   U755 : MUX2DL port map( A0 => operand_regs_161_port, A1 => 
                           coeff_memory_1_1_port, SL => n718, Z => N2946);
   U756 : MUX2DL port map( A0 => operand_regs_225_port, A1 => 
                           coeff_memory_0_1_port, SL => n716, Z => N2914);
   U757 : INVD1 port map( A => n705, Z => n701);
   U758 : INVD1 port map( A => filt_mult_inputs, Z => n705);
   U759 : MUX2DL port map( A0 => operand_regs_37_port, A1 => 
                           coeff_memory_3_5_port, SL => n712, Z => N3014);
   U760 : MUX2DL port map( A0 => operand_regs_101_port, A1 => 
                           coeff_memory_2_5_port, SL => n711, Z => N2982);
   U761 : MUX2DL port map( A0 => operand_regs_5_port, A1 => 
                           coeff_memory_4_5_port, SL => n714, Z => N3046);
   U762 : MUX2DL port map( A0 => operand_regs_165_port, A1 => 
                           coeff_memory_1_5_port, SL => n718, Z => N2950);
   U763 : MUX2DL port map( A0 => operand_regs_229_port, A1 => 
                           coeff_memory_0_5_port, SL => n715, Z => N2918);
   U764 : MUX2DL port map( A0 => operand_regs_34_port, A1 => 
                           coeff_memory_3_2_port, SL => n712, Z => N3011);
   U765 : MUX2DL port map( A0 => operand_regs_98_port, A1 => 
                           coeff_memory_2_2_port, SL => n710, Z => N2979);
   U766 : MUX2DL port map( A0 => operand_regs_35_port, A1 => 
                           coeff_memory_3_3_port, SL => n712, Z => N3012);
   U767 : MUX2DL port map( A0 => operand_regs_99_port, A1 => 
                           coeff_memory_2_3_port, SL => n710, Z => N2980);
   U768 : MUX2DL port map( A0 => operand_regs_2_port, A1 => 
                           coeff_memory_4_2_port, SL => n714, Z => N3043);
   U769 : MUX2DL port map( A0 => operand_regs_162_port, A1 => 
                           coeff_memory_1_2_port, SL => n717, Z => N2947);
   U770 : MUX2DL port map( A0 => operand_regs_226_port, A1 => 
                           coeff_memory_0_2_port, SL => n716, Z => N2915);
   U771 : MUX2DL port map( A0 => operand_regs_39_port, A1 => 
                           coeff_memory_3_7_port, SL => n712, Z => N3016);
   U772 : MUX2DL port map( A0 => operand_regs_103_port, A1 => 
                           coeff_memory_2_7_port, SL => n711, Z => N2984);
   U773 : MUX2DL port map( A0 => operand_regs_3_port, A1 => 
                           coeff_memory_4_3_port, SL => n714, Z => N3044);
   U774 : MUX2DL port map( A0 => operand_regs_163_port, A1 => 
                           coeff_memory_1_3_port, SL => n718, Z => N2948);
   U775 : MUX2DL port map( A0 => operand_regs_227_port, A1 => 
                           coeff_memory_0_3_port, SL => n716, Z => N2916);
   U776 : MUX2DL port map( A0 => operand_regs_7_port, A1 => 
                           coeff_memory_4_7_port, SL => n714, Z => N3048);
   U777 : MUX2DL port map( A0 => operand_regs_167_port, A1 => 
                           coeff_memory_1_7_port, SL => n718, Z => N2952);
   U778 : MUX2DL port map( A0 => operand_regs_231_port, A1 => 
                           coeff_memory_0_7_port, SL => n715, Z => N2920);
   U779 : MUX2DL port map( A0 => operand_regs_38_port, A1 => 
                           coeff_memory_3_6_port, SL => n712, Z => N3015);
   U780 : MUX2DL port map( A0 => operand_regs_102_port, A1 => 
                           coeff_memory_2_6_port, SL => n711, Z => N2983);
   U781 : MUX2DL port map( A0 => operand_regs_6_port, A1 => 
                           coeff_memory_4_6_port, SL => n714, Z => N3047);
   U782 : MUX2DL port map( A0 => operand_regs_166_port, A1 => 
                           coeff_memory_1_6_port, SL => n717, Z => N2951);
   U783 : MUX2DL port map( A0 => operand_regs_230_port, A1 => 
                           coeff_memory_0_6_port, SL => n715, Z => N2919);
   U784 : MUX2DL port map( A0 => operand_regs_36_port, A1 => 
                           coeff_memory_3_4_port, SL => n712, Z => N3013);
   U785 : MUX2DL port map( A0 => operand_regs_100_port, A1 => 
                           coeff_memory_2_4_port, SL => n711, Z => N2981);
   U786 : MUX2DL port map( A0 => operand_regs_104_port, A1 => 
                           coeff_memory_2_8_port, SL => n711, Z => N2985);
   U787 : MUX2DL port map( A0 => operand_regs_40_port, A1 => 
                           coeff_memory_3_8_port, SL => n709, Z => N3017);
   U788 : MUX2DL port map( A0 => operand_regs_4_port, A1 => 
                           coeff_memory_4_4_port, SL => n714, Z => N3045);
   U789 : MUX2DL port map( A0 => operand_regs_164_port, A1 => 
                           coeff_memory_1_4_port, SL => n717, Z => N2949);
   U790 : MUX2DL port map( A0 => operand_regs_228_port, A1 => 
                           coeff_memory_0_4_port, SL => n716, Z => N2917);
   U791 : MUX2DL port map( A0 => operand_regs_8_port, A1 => 
                           coeff_memory_4_8_port, SL => n714, Z => N3049);
   U792 : MUX2DL port map( A0 => operand_regs_168_port, A1 => 
                           coeff_memory_1_8_port, SL => n717, Z => N2953);
   U793 : MUX2DL port map( A0 => operand_regs_232_port, A1 => 
                           coeff_memory_0_8_port, SL => n715, Z => N2921);
   U794 : MUX2DL port map( A0 => operand_regs_6_port, A1 => 
                           operand_regs_198_port, SL => n720, Z => n278);
   U795 : MUX2DL port map( A0 => operand_regs_7_port, A1 => 
                           operand_regs_199_port, SL => n719, Z => n279);
   U796 : MUX2DL port map( A0 => operand_regs_43_port, A1 => 
                           coeff_memory_3_11_port, SL => n711, Z => N3020);
   U797 : MUX2DL port map( A0 => operand_regs_107_port, A1 => 
                           coeff_memory_2_11_port, SL => n711, Z => N2988);
   U798 : MUX2DL port map( A0 => operand_regs_8_port, A1 => 
                           operand_regs_200_port, SL => n720, Z => n280);
   U799 : MUX2DL port map( A0 => operand_regs_11_port, A1 => 
                           coeff_memory_4_11_port, SL => n713, Z => N3052);
   U800 : MUX2DL port map( A0 => operand_regs_171_port, A1 => 
                           coeff_memory_1_11_port, SL => n718, Z => N2956);
   U801 : MUX2DL port map( A0 => operand_regs_235_port, A1 => 
                           coeff_memory_0_11_port, SL => n715, Z => N2924);
   U802 : MUX2DL port map( A0 => operand_regs_9_port, A1 => 
                           operand_regs_201_port, SL => n719, Z => n281);
   U803 : MUX2DL port map( A0 => operand_regs_5_port, A1 => 
                           operand_regs_197_port, SL => n719, Z => n282);
   U804 : MUX2DL port map( A0 => operand_regs_1_port, A1 => 
                           operand_regs_193_port, SL => n720, Z => n283);
   U805 : MUX2DL port map( A0 => operand_regs_2_port, A1 => 
                           operand_regs_194_port, SL => n720, Z => n284);
   U806 : MUX2DL port map( A0 => operand_regs_44_port, A1 => 
                           coeff_memory_3_12_port, SL => n711, Z => N3021);
   U807 : MUX2DL port map( A0 => operand_regs_108_port, A1 => 
                           coeff_memory_2_12_port, SL => n711, Z => N2989);
   U808 : MUX2DL port map( A0 => operand_regs_10_port, A1 => 
                           operand_regs_202_port, SL => n720, Z => n285);
   U809 : MUX2DL port map( A0 => operand_regs_41_port, A1 => 
                           coeff_memory_3_9_port, SL => n712, Z => N3018);
   U810 : MUX2DL port map( A0 => operand_regs_105_port, A1 => 
                           coeff_memory_2_9_port, SL => n711, Z => N2986);
   U811 : MUX2DL port map( A0 => operand_regs_12_port, A1 => 
                           coeff_memory_4_12_port, SL => n713, Z => N3053);
   U812 : MUX2DL port map( A0 => operand_regs_172_port, A1 => 
                           coeff_memory_1_12_port, SL => n717, Z => N2957);
   U813 : MUX2DL port map( A0 => operand_regs_236_port, A1 => 
                           coeff_memory_0_12_port, SL => n715, Z => N2925);
   U814 : MUX2DL port map( A0 => operand_regs_9_port, A1 => 
                           coeff_memory_4_9_port, SL => n713, Z => N3050);
   U815 : MUX2DL port map( A0 => operand_regs_169_port, A1 => 
                           coeff_memory_1_9_port, SL => n718, Z => N2954);
   U816 : MUX2DL port map( A0 => operand_regs_233_port, A1 => 
                           coeff_memory_0_9_port, SL => n715, Z => N2922);
   U817 : MUX2DL port map( A0 => operand_regs_3_port, A1 => 
                           operand_regs_195_port, SL => n720, Z => n286);
   U818 : MUX2DL port map( A0 => operand_regs_45_port, A1 => 
                           coeff_memory_3_13_port, SL => n711, Z => N3022);
   U819 : MUX2DL port map( A0 => operand_regs_109_port, A1 => 
                           coeff_memory_2_13_port, SL => n711, Z => N2990);
   U820 : MUX2DL port map( A0 => operand_regs_47_port, A1 => 
                           coeff_memory_3_15_port, SL => n711, Z => N3024);
   U821 : MUX2DL port map( A0 => operand_regs_111_port, A1 => 
                           coeff_memory_2_15_port, SL => n712, Z => N2992);
   U822 : MUX2DL port map( A0 => operand_regs_4_port, A1 => 
                           operand_regs_196_port, SL => n720, Z => n287);
   U823 : MUX2DL port map( A0 => operand_regs_13_port, A1 => 
                           coeff_memory_4_13_port, SL => n713, Z => N3054);
   U824 : MUX2DL port map( A0 => operand_regs_173_port, A1 => 
                           coeff_memory_1_13_port, SL => n718, Z => N2958);
   U825 : MUX2DL port map( A0 => operand_regs_237_port, A1 => 
                           coeff_memory_0_13_port, SL => n715, Z => N2926);
   U826 : MUX2DL port map( A0 => operand_regs_15_port, A1 => 
                           coeff_memory_4_15_port, SL => n713, Z => N3056);
   U827 : MUX2DL port map( A0 => operand_regs_175_port, A1 => 
                           coeff_memory_1_15_port, SL => n718, Z => N2960);
   U828 : MUX2DL port map( A0 => operand_regs_239_port, A1 => 
                           coeff_memory_0_15_port, SL => n715, Z => N2928);
   U829 : MUX2DL port map( A0 => operand_regs_192_port, A1 => 
                           operand_regs_0_port, SL => n721, Z => n288);
   U830 : INVD1 port map( A => operand_regs_198_port, Z => n755);
   U831 : INVD1 port map( A => operand_regs_199_port, Z => n754);
   U832 : MUX2DL port map( A0 => operand_regs_46_port, A1 => 
                           coeff_memory_3_14_port, SL => n711, Z => N3023);
   U833 : MUX2DL port map( A0 => operand_regs_110_port, A1 => 
                           coeff_memory_2_14_port, SL => n711, Z => N2991);
   U834 : INVD1 port map( A => operand_regs_200_port, Z => n753);
   U835 : MUX2DL port map( A0 => operand_regs_14_port, A1 => 
                           coeff_memory_4_14_port, SL => n713, Z => N3055);
   U836 : MUX2DL port map( A0 => operand_regs_174_port, A1 => 
                           coeff_memory_1_14_port, SL => n717, Z => N2959);
   U837 : MUX2DL port map( A0 => operand_regs_238_port, A1 => 
                           coeff_memory_0_14_port, SL => n715, Z => N2927);
   U838 : INVD1 port map( A => operand_regs_194_port, Z => n759);
   U839 : INVD1 port map( A => operand_regs_193_port, Z => n760);
   U840 : INVD1 port map( A => operand_regs_197_port, Z => n756);
   U841 : MUX2DL port map( A0 => operand_regs_48_port, A1 => 
                           coeff_memory_3_16_port, SL => n709, Z => N3025);
   U842 : MUX2DL port map( A0 => operand_regs_16_port, A1 => 
                           coeff_memory_4_16_port, SL => n713, Z => N3057);
   U843 : MUX2DL port map( A0 => operand_regs_112_port, A1 => 
                           coeff_memory_2_16_port, SL => n717, Z => N2993);
   U844 : MUX2DL port map( A0 => operand_regs_176_port, A1 => 
                           coeff_memory_1_16_port, SL => n717, Z => N2961);
   U845 : MUX2DL port map( A0 => operand_regs_240_port, A1 => 
                           coeff_memory_0_16_port, SL => n715, Z => N2929);
   U846 : MUX2DL port map( A0 => operand_regs_49_port, A1 => 
                           coeff_memory_3_17_port, SL => n709, Z => N3026);
   U847 : MUX2DL port map( A0 => operand_regs_17_port, A1 => 
                           coeff_memory_4_17_port, SL => n713, Z => N3058);
   U848 : MUX2DL port map( A0 => operand_regs_113_port, A1 => 
                           coeff_memory_2_17_port, SL => n719, Z => N2994);
   U849 : MUX2DL port map( A0 => operand_regs_177_port, A1 => 
                           coeff_memory_1_17_port, SL => n717, Z => N2962);
   U850 : MUX2DL port map( A0 => operand_regs_241_port, A1 => 
                           coeff_memory_0_17_port, SL => n715, Z => N2930);
   U851 : MUX2DL port map( A0 => operand_regs_42_port, A1 => 
                           coeff_memory_3_10_port, SL => n711, Z => N3019);
   U852 : MUX2DL port map( A0 => operand_regs_106_port, A1 => 
                           coeff_memory_2_10_port, SL => n711, Z => N2987);
   U853 : INVD1 port map( A => operand_regs_195_port, Z => n758);
   U854 : MUX2DL port map( A0 => operand_regs_10_port, A1 => 
                           coeff_memory_4_10_port, SL => n713, Z => N3051);
   U855 : MUX2DL port map( A0 => operand_regs_170_port, A1 => 
                           coeff_memory_1_10_port, SL => n717, Z => N2955);
   U856 : MUX2DL port map( A0 => operand_regs_234_port, A1 => 
                           coeff_memory_0_10_port, SL => n715, Z => N2923);
   U857 : INVD1 port map( A => operand_regs_192_port, Z => n761);
   U858 : INVD1 port map( A => operand_regs_196_port, Z => n757);
   U859 : MUX2DL port map( A0 => operand_regs_50_port, A1 => 
                           coeff_memory_3_18_port, SL => n709, Z => N3027);
   U860 : MUX2DL port map( A0 => operand_regs_18_port, A1 => 
                           coeff_memory_4_18_port, SL => n713, Z => N3059);
   U861 : MUX2DL port map( A0 => operand_regs_114_port, A1 => 
                           coeff_memory_2_18_port, SL => n718, Z => N2995);
   U862 : MUX2DL port map( A0 => operand_regs_178_port, A1 => 
                           coeff_memory_1_18_port, SL => n717, Z => N2963);
   U863 : MUX2DL port map( A0 => operand_regs_242_port, A1 => 
                           coeff_memory_0_18_port, SL => n715, Z => N2931);
   U864 : INVD1 port map( A => operand_regs_201_port, Z => n752);
   U865 : MUX2DL port map( A0 => operand_regs_96_port, A1 => 
                           coeff_memory_2_0_port, SL => n710, Z => N2977);
   U866 : MUX2DL port map( A0 => operand_regs_51_port, A1 => 
                           coeff_memory_3_19_port, SL => n710, Z => N3028);
   U867 : MUX2DL port map( A0 => operand_regs_32_port, A1 => 
                           coeff_memory_3_0_port, SL => n712, Z => N3009);
   U868 : MUX2DL port map( A0 => operand_regs_160_port, A1 => 
                           coeff_memory_1_0_port, SL => n717, Z => N2945);
   U869 : MUX2DL port map( A0 => operand_regs_19_port, A1 => 
                           coeff_memory_4_19_port, SL => n713, Z => N3060);
   U870 : MUX2DL port map( A0 => operand_regs_115_port, A1 => 
                           coeff_memory_2_19_port, SL => n719, Z => N2996);
   U871 : MUX2DL port map( A0 => operand_regs_179_port, A1 => 
                           coeff_memory_1_19_port, SL => n717, Z => N2964);
   U872 : MUX2DL port map( A0 => operand_regs_243_port, A1 => 
                           coeff_memory_0_19_port, SL => n715, Z => N2932);
   U873 : MUX2DL port map( A0 => operand_regs_224_port, A1 => 
                           coeff_memory_0_0_port, SL => n716, Z => N2913);
   U874 : MUX2DL port map( A0 => operand_regs_0_port, A1 => 
                           coeff_memory_4_0_port, SL => n714, Z => N3041);
   U875 : INVD1 port map( A => operand_regs_202_port, Z => n751);
   U876 : MUX2DL port map( A0 => operand_regs_17_port, A1 => 
                           operand_regs_209_port, SL => n719, Z => n289);
   U877 : MUX2DL port map( A0 => operand_regs_18_port, A1 => 
                           operand_regs_210_port, SL => n720, Z => n290);
   U878 : INVD1 port map( A => operand_regs_204_port, Z => n749);
   U879 : MUX2DL port map( A0 => operand_regs_15_port, A1 => 
                           operand_regs_207_port, SL => n719, Z => n291);
   U880 : INVD1 port map( A => operand_regs_203_port, Z => n750);
   U881 : MUX2DL port map( A0 => operand_regs_16_port, A1 => 
                           operand_regs_208_port, SL => n720, Z => n292);
   U882 : MUX2DL port map( A0 => operand_regs_52_port, A1 => 
                           coeff_memory_3_20_port, SL => n710, Z => N3029);
   U883 : INVD1 port map( A => operand_regs_205_port, Z => n748);
   U884 : MUX2DL port map( A0 => operand_regs_20_port, A1 => 
                           coeff_memory_4_20_port, SL => n713, Z => N3061);
   U885 : MUX2DL port map( A0 => operand_regs_116_port, A1 => 
                           coeff_memory_2_20_port, SL => n718, Z => N2997);
   U886 : MUX2DL port map( A0 => operand_regs_180_port, A1 => 
                           coeff_memory_1_20_port, SL => n717, Z => N2965);
   U887 : MUX2DL port map( A0 => operand_regs_244_port, A1 => 
                           coeff_memory_0_20_port, SL => n715, Z => N2933);
   U888 : INVD1 port map( A => operand_regs_206_port, Z => n747);
   U889 : INVD1 port map( A => operand_regs_209_port, Z => n744);
   U890 : MUX2DL port map( A0 => operand_regs_19_port, A1 => 
                           operand_regs_211_port, SL => n719, Z => n293);
   U891 : INVD1 port map( A => operand_regs_207_port, Z => n746);
   U892 : MUX2DL port map( A0 => operand_regs_20_port, A1 => 
                           operand_regs_212_port, SL => n720, Z => n294);
   U893 : INVD1 port map( A => operand_regs_210_port, Z => n743);
   U894 : INVD1 port map( A => operand_regs_208_port, Z => n745);
   U895 : INVD1 port map( A => operand_regs_211_port, Z => n742);
   U896 : INVD1 port map( A => operand_regs_212_port, Z => n741);
   U897 : MUX2DL port map( A0 => operand_regs_53_port, A1 => 
                           coeff_memory_3_21_port, SL => n710, Z => N3030);
   U898 : MUX2DL port map( A0 => operand_regs_21_port, A1 => 
                           coeff_memory_4_21_port, SL => n713, Z => N3062);
   U899 : MUX2DL port map( A0 => operand_regs_117_port, A1 => 
                           coeff_memory_2_21_port, SL => n719, Z => N2998);
   U900 : MUX2DL port map( A0 => operand_regs_181_port, A1 => 
                           coeff_memory_1_21_port, SL => n716, Z => N2966);
   U901 : MUX2DL port map( A0 => operand_regs_245_port, A1 => 
                           coeff_memory_0_21_port, SL => n715, Z => N2934);
   U902 : MUX2DL port map( A0 => operand_regs_21_port, A1 => 
                           operand_regs_213_port, SL => n719, Z => n295);
   U903 : MUX2DL port map( A0 => operand_regs_54_port, A1 => 
                           coeff_memory_3_22_port, SL => n710, Z => N3031);
   U904 : MUX2DL port map( A0 => operand_regs_22_port, A1 => 
                           coeff_memory_4_22_port, SL => n713, Z => N3063);
   U905 : MUX2DL port map( A0 => operand_regs_118_port, A1 => 
                           coeff_memory_2_22_port, SL => n717, Z => N2999);
   U906 : MUX2DL port map( A0 => operand_regs_182_port, A1 => 
                           coeff_memory_1_22_port, SL => n716, Z => N2967);
   U907 : MUX2DL port map( A0 => operand_regs_246_port, A1 => 
                           coeff_memory_0_22_port, SL => n714, Z => N2935);
   U908 : MUX2DL port map( A0 => operand_regs_22_port, A1 => 
                           operand_regs_214_port, SL => n720, Z => n296);
   U909 : INVD1 port map( A => operand_regs_213_port, Z => n740);
   U910 : INVD1 port map( A => operand_regs_214_port, Z => n739);
   U911 : MUX2DL port map( A0 => operand_regs_55_port, A1 => 
                           coeff_memory_3_23_port, SL => n710, Z => N3032);
   U912 : MUX2DL port map( A0 => operand_regs_23_port, A1 => 
                           coeff_memory_4_23_port, SL => n713, Z => N3064);
   U913 : MUX2DL port map( A0 => operand_regs_119_port, A1 => 
                           coeff_memory_2_23_port, SL => n718, Z => N3000);
   U914 : MUX2DL port map( A0 => operand_regs_183_port, A1 => 
                           coeff_memory_1_23_port, SL => n716, Z => N2968);
   U915 : MUX2DL port map( A0 => operand_regs_247_port, A1 => 
                           coeff_memory_0_23_port, SL => n714, Z => N2936);
   U916 : MUX2DL port map( A0 => operand_regs_56_port, A1 => 
                           coeff_memory_3_24_port, SL => n710, Z => N3033);
   U917 : MUX2DL port map( A0 => operand_regs_24_port, A1 => 
                           coeff_memory_4_24_port, SL => n713, Z => N3065);
   U918 : MUX2DL port map( A0 => operand_regs_120_port, A1 => 
                           coeff_memory_2_24_port, SL => n718, Z => N3001);
   U919 : MUX2DL port map( A0 => operand_regs_184_port, A1 => 
                           coeff_memory_1_24_port, SL => n716, Z => N2969);
   U920 : MUX2DL port map( A0 => operand_regs_248_port, A1 => 
                           coeff_memory_0_24_port, SL => n714, Z => N2937);
   U921 : MUX2DL port map( A0 => operand_regs_23_port, A1 => 
                           operand_regs_215_port, SL => n719, Z => n297);
   U922 : INVD1 port map( A => operand_regs_215_port, Z => n738);
   U923 : MUX2DL port map( A0 => operand_regs_57_port, A1 => 
                           coeff_memory_3_25_port, SL => n710, Z => N3034);
   U924 : MUX2DL port map( A0 => operand_regs_25_port, A1 => 
                           coeff_memory_4_25_port, SL => n713, Z => N3066);
   U925 : MUX2DL port map( A0 => operand_regs_121_port, A1 => 
                           coeff_memory_2_25_port, SL => n718, Z => N3002);
   U926 : MUX2DL port map( A0 => operand_regs_185_port, A1 => 
                           coeff_memory_1_25_port, SL => n716, Z => N2970);
   U927 : MUX2DL port map( A0 => operand_regs_249_port, A1 => 
                           coeff_memory_0_25_port, SL => n714, Z => N2938);
   U928 : NOR3M1D1 port map( A1 => n104, A2 => coeff_load, A3 => operand_load, 
                           Z => n110);
   U929 : AND2D1 port map( A1 => N66, A2 => avs_write, Z => n104);
   U930 : MUX2DL port map( A0 => operand_regs_24_port, A1 => 
                           operand_regs_216_port, SL => n720, Z => n298);
   U931 : INVD1 port map( A => operand_regs_216_port, Z => n737);
   U932 : MUX2DL port map( A0 => operand_regs_25_port, A1 => 
                           operand_regs_217_port, SL => n719, Z => n299);
   U933 : MUX2DL port map( A0 => operand_regs_26_port, A1 => 
                           coeff_memory_4_26_port, SL => n712, Z => N3067);
   U934 : MUX2DL port map( A0 => operand_regs_58_port, A1 => 
                           coeff_memory_3_26_port, SL => n710, Z => N3035);
   U935 : MUX2DL port map( A0 => operand_regs_122_port, A1 => 
                           coeff_memory_2_26_port, SL => n718, Z => N3003);
   U936 : MUX2DL port map( A0 => operand_regs_186_port, A1 => 
                           coeff_memory_1_26_port, SL => n716, Z => N2971);
   U937 : MUX2DL port map( A0 => operand_regs_250_port, A1 => 
                           coeff_memory_0_26_port, SL => n714, Z => N2939);
   U938 : INVD1 port map( A => coeff_load, Z => n729);
   U939 : INVD1 port map( A => operand_regs_217_port, Z => n736);
   U940 : NAN4D1 port map( A1 => n5900, A2 => n14, A3 => n6000, A4 => n6100, Z 
                           => n233);
   U941 : NAN2M1D1 port map( A1 => n70, A2 => n300, Z => n5900);
   U942 : NAN2D1 port map( A1 => N2009, A2 => n268, Z => n6000);
   U943 : INVD1 port map( A => avs_write, Z => n799);
   U944 : AND2D1 port map( A1 => avs_read, A2 => n799, Z => n300);
   U945 : INVD1 port map( A => n12, Z => n699);
   U946 : NOR3M1D1 port map( A1 => N66, A2 => n700, A3 => read_comp_res, Z => 
                           n12);
   U947 : NAN3D1 port map( A1 => n56, A2 => n14, A3 => n57, Z => n231);
   U948 : NAN2D1 port map( A1 => N2007, A2 => n268, Z => n56);
   U949 : NAN3D1 port map( A1 => n452, A2 => n451, A3 => n453, Z => N2007);
   U950 : NAN3D1 port map( A1 => n53, A2 => n14, A3 => n54, Z => n229);
   U951 : NAN2D1 port map( A1 => N2005, A2 => n268, Z => n53);
   U952 : NAN3D1 port map( A1 => n458, A2 => n457, A3 => n459, Z => N2005);
   U953 : NAN3D1 port map( A1 => n50, A2 => n14, A3 => n51, Z => n227);
   U954 : NAN2D1 port map( A1 => N2003, A2 => n268, Z => n50);
   U955 : NAN3D1 port map( A1 => n464, A2 => n463, A3 => n465, Z => N2003);
   U956 : NAN3D1 port map( A1 => n47, A2 => n14, A3 => n48, Z => n225);
   U957 : NAN2D1 port map( A1 => N2001, A2 => n268, Z => n47);
   U958 : NAN3D1 port map( A1 => n470, A2 => n469, A3 => n471, Z => N2001);
   U959 : NAN3D1 port map( A1 => n44, A2 => n14, A3 => n45, Z => n223);
   U960 : NAN2D1 port map( A1 => N1999, A2 => n268, Z => n44);
   U961 : NAN3D1 port map( A1 => n476, A2 => n475, A3 => n477, Z => N1999);
   U962 : NAN3D1 port map( A1 => n41, A2 => n14, A3 => n42, Z => n221);
   U963 : NAN2D1 port map( A1 => N1997, A2 => n268, Z => n41);
   U964 : NAN3D1 port map( A1 => n482, A2 => n481, A3 => n483, Z => N1997);
   U965 : NAN3D1 port map( A1 => n38, A2 => n14, A3 => n39, Z => n219);
   U966 : NAN2D1 port map( A1 => N1995, A2 => n268, Z => n38);
   U967 : NAN3D1 port map( A1 => n488, A2 => n487, A3 => n489, Z => N1995);
   U968 : NAN3D1 port map( A1 => n35, A2 => n14, A3 => n36, Z => n217);
   U969 : NAN2D1 port map( A1 => N1993, A2 => n268, Z => n35);
   U970 : NAN3D1 port map( A1 => n494, A2 => n493, A3 => n495, Z => N1993);
   U971 : NAN3D1 port map( A1 => n13, A2 => n14, A3 => n15, Z => n203);
   U972 : NAN2D1 port map( A1 => N1979, A2 => n268, Z => n13);
   U973 : NAN3D1 port map( A1 => n536, A2 => n535, A3 => n537, Z => N1979);
   U974 : INVD1 port map( A => avs_addr(2), Z => n547);
   U975 : NAN3D1 port map( A1 => n32, A2 => n14, A3 => n33, Z => n215);
   U976 : NAN2D1 port map( A1 => N1991, A2 => n268, Z => n32);
   U977 : NAN3D1 port map( A1 => n500, A2 => n499, A3 => n501, Z => N1991);
   U978 : NAN3D1 port map( A1 => n29, A2 => n14, A3 => n30, Z => n213);
   U979 : NAN2D1 port map( A1 => N1989, A2 => n268, Z => n29);
   U980 : NAN3D1 port map( A1 => n506, A2 => n505, A3 => n507, Z => N1989);
   U981 : NAN3D1 port map( A1 => n26, A2 => n14, A3 => n27, Z => n211);
   U982 : NAN2D1 port map( A1 => N1987, A2 => n268, Z => n26);
   U983 : NAN3D1 port map( A1 => n512, A2 => n511, A3 => n513, Z => N1987);
   U984 : NAN3D1 port map( A1 => n23, A2 => n14, A3 => n24, Z => n209);
   U985 : NAN2D1 port map( A1 => N1985, A2 => n268, Z => n23);
   U986 : NAN3D1 port map( A1 => n518, A2 => n517, A3 => n519, Z => N1985);
   U987 : NAN3D1 port map( A1 => n20, A2 => n14, A3 => n21, Z => n207);
   U988 : NAN2D1 port map( A1 => N1983, A2 => n268, Z => n20);
   U989 : NAN3D1 port map( A1 => n524, A2 => n523, A3 => n525, Z => N1983);
   U990 : NAN3D1 port map( A1 => n17, A2 => n14, A3 => n18, Z => n205);
   U991 : NAN2D1 port map( A1 => N1981, A2 => n268, Z => n17);
   U992 : NAN3D1 port map( A1 => n530, A2 => n529, A3 => n531, Z => N1981);
   U993 : OAI21M20D1 port map( A1 => avs_readdata_1_port, A2 => n700, B => n58,
                           Z => n232);
   U994 : NAN3D1 port map( A1 => n449, A2 => n448, A3 => n450, Z => N2008);
   U995 : OAI21M20D1 port map( A1 => avs_readdata_3_port, A2 => n700, B => n55,
                           Z => n230);
   U996 : NAN3D1 port map( A1 => n455, A2 => n454, A3 => n456, Z => N2006);
   U997 : OAI21M20D1 port map( A1 => avs_readdata_5_port, A2 => n700, B => n52,
                           Z => n228);
   U998 : NAN3D1 port map( A1 => n461, A2 => n460, A3 => n462, Z => N2004);
   U999 : OAI21M20D1 port map( A1 => avs_readdata_7_port, A2 => n700, B => n49,
                           Z => n226);
   U1000 : NAN3D1 port map( A1 => n467, A2 => n466, A3 => n468, Z => N2002);
   U1001 : OAI21M20D1 port map( A1 => avs_readdata_15_port, A2 => n700, B => 
                           n37, Z => n218);
   U1002 : NAN3D1 port map( A1 => n491, A2 => n490, A3 => n492, Z => N1994);
   U1003 : OAI21M20D1 port map( A1 => avs_readdata_17_port, A2 => n700, B => 
                           n34, Z => n216);
   U1004 : NAN3D1 port map( A1 => n497, A2 => n496, A3 => n498, Z => N1992);
   U1005 : OAI21M20D1 port map( A1 => avs_readdata_19_port, A2 => n700, B => 
                           n31, Z => n214);
   U1006 : NAN3D1 port map( A1 => n503, A2 => n502, A3 => n504, Z => N1990);
   U1007 : OAI21M20D1 port map( A1 => avs_readdata_21_port, A2 => n700, B => 
                           n28, Z => n212);
   U1008 : NAN3D1 port map( A1 => n509, A2 => n508, A3 => n510, Z => N1988);
   U1009 : OAI21M20D1 port map( A1 => avs_readdata_23_port, A2 => n700, B => 
                           n25, Z => n210);
   U1010 : NAN3D1 port map( A1 => n515, A2 => n514, A3 => n516, Z => N1986);
   U1011 : OAI21M20D1 port map( A1 => avs_readdata_25_port, A2 => n700, B => 
                           n22, Z => n208);
   U1012 : NAN3D1 port map( A1 => n521, A2 => n520, A3 => n522, Z => N1984);
   U1013 : OAI21M20D1 port map( A1 => avs_readdata_27_port, A2 => n700, B => 
                           n19, Z => n206);
   U1014 : NAN3D1 port map( A1 => n527, A2 => n526, A3 => n528, Z => N1982);
   U1015 : OAI21M20D1 port map( A1 => avs_readdata_29_port, A2 => n700, B => 
                           n16, Z => n204);
   U1016 : NAN3D1 port map( A1 => n533, A2 => n532, A3 => n534, Z => N1980);
   U1017 : OAI21M20D1 port map( A1 => avs_readdata_31_port, A2 => n700, B => 
                           n10, Z => n202);
   U1018 : OAI21M20D1 port map( A1 => avs_readdata_9_port, A2 => n700, B => n46
                           , Z => n224);
   U1019 : NAN3D1 port map( A1 => n473, A2 => n472, A3 => n474, Z => N2000);
   U1020 : OAI21M20D1 port map( A1 => avs_readdata_11_port, A2 => n700, B => 
                           n43, Z => n222);
   U1021 : NAN3D1 port map( A1 => n479, A2 => n478, A3 => n480, Z => N1998);
   U1022 : OAI21M20D1 port map( A1 => avs_readdata_13_port, A2 => n700, B => 
                           n40, Z => n220);
   U1023 : NAN3D1 port map( A1 => n485, A2 => n484, A3 => n486, Z => N1996);
   U1024 : AND2D1 port map( A1 => coeff_load, A2 => n104, Z => n301);
   U1025 : MUX2DL port map( A0 => operand_regs_27_port, A1 => 
                           coeff_memory_4_27_port, SL => n712, Z => N3068);
   U1026 : MUX2DL port map( A0 => operand_regs_59_port, A1 => 
                           coeff_memory_3_27_port, SL => n710, Z => N3036);
   U1027 : MUX2DL port map( A0 => operand_regs_123_port, A1 => 
                           coeff_memory_2_27_port, SL => n718, Z => N3004);
   U1028 : MUX2DL port map( A0 => operand_regs_187_port, A1 => 
                           coeff_memory_1_27_port, SL => n716, Z => N2972);
   U1029 : MUX2DL port map( A0 => operand_regs_251_port, A1 => 
                           coeff_memory_0_27_port, SL => n714, Z => N2940);
   U1030 : NAN3D1 port map( A1 => n545, A2 => n544, A3 => n546, Z => N1978);
   U1031 : NAN2D1 port map( A1 => comp_res_31_port, A2 => n554, Z => n545);
   U1032 : AOI22M10D1 port map( B1 => in_buf_63_port, B2 => n540, A1 => n553, 
                           A2 => in_buf_127_port, Z => n442);
   U1033 : NAN3D1 port map( A1 => n446, A2 => n445, A3 => n447, Z => N2009);
   U1034 : NAN2D1 port map( A1 => comp_res_0_port, A2 => n554, Z => n446);
   U1035 : MUX2DL port map( A0 => operand_regs_26_port, A1 => 
                           operand_regs_218_port, SL => n720, Z => n302);
   U1036 : NAN2D1 port map( A1 => comp_res_25_port, A2 => n554, Z => n521);
   U1037 : NAN2D1 port map( A1 => comp_res_27_port, A2 => n554, Z => n527);
   U1038 : NAN2D1 port map( A1 => comp_res_29_port, A2 => n554, Z => n533);
   U1039 : NAN2D1 port map( A1 => comp_res_1_port, A2 => n554, Z => n449);
   U1040 : NAN2D1 port map( A1 => comp_res_3_port, A2 => n541, Z => n455);
   U1041 : NAN2D1 port map( A1 => comp_res_5_port, A2 => n541, Z => n461);
   U1042 : NAN2D1 port map( A1 => comp_res_7_port, A2 => n554, Z => n467);
   U1043 : NAN2D1 port map( A1 => comp_res_9_port, A2 => n541, Z => n473);
   U1044 : NAN2D1 port map( A1 => comp_res_11_port, A2 => n554, Z => n479);
   U1045 : NAN2D1 port map( A1 => comp_res_13_port, A2 => n554, Z => n485);
   U1046 : NAN2D1 port map( A1 => comp_res_15_port, A2 => n554, Z => n491);
   U1047 : NAN2D1 port map( A1 => comp_res_17_port, A2 => n554, Z => n497);
   U1048 : NAN2D1 port map( A1 => comp_res_19_port, A2 => n554, Z => n503);
   U1049 : NAN2D1 port map( A1 => comp_res_21_port, A2 => n554, Z => n509);
   U1050 : NAN2D1 port map( A1 => comp_res_23_port, A2 => n554, Z => n515);
   U1051 : NAN2D1 port map( A1 => comp_res_24_port, A2 => n554, Z => n518);
   U1052 : NAN2D1 port map( A1 => comp_res_26_port, A2 => n554, Z => n524);
   U1053 : NAN2D1 port map( A1 => comp_res_28_port, A2 => n554, Z => n530);
   U1054 : NAN2D1 port map( A1 => comp_res_30_port, A2 => n554, Z => n536);
   U1055 : NAN2D1 port map( A1 => comp_res_2_port, A2 => n541, Z => n452);
   U1056 : NAN2D1 port map( A1 => comp_res_4_port, A2 => n541, Z => n458);
   U1057 : NAN2D1 port map( A1 => comp_res_6_port, A2 => n541, Z => n464);
   U1058 : NAN2D1 port map( A1 => comp_res_8_port, A2 => n541, Z => n470);
   U1059 : NAN2D1 port map( A1 => comp_res_10_port, A2 => n541, Z => n476);
   U1060 : NAN2D1 port map( A1 => comp_res_12_port, A2 => n541, Z => n482);
   U1061 : NAN2D1 port map( A1 => comp_res_14_port, A2 => n541, Z => n488);
   U1062 : NAN2D1 port map( A1 => comp_res_16_port, A2 => n541, Z => n494);
   U1063 : NAN2D1 port map( A1 => comp_res_18_port, A2 => n541, Z => n500);
   U1064 : NAN2D1 port map( A1 => comp_res_20_port, A2 => n541, Z => n506);
   U1065 : NAN2D1 port map( A1 => comp_res_22_port, A2 => n541, Z => n512);
   U1066 : INVD1 port map( A => operand_regs_218_port, Z => n735);
   U1067 : MUX2DL port map( A0 => operand_regs_27_port, A1 => 
                           operand_regs_219_port, SL => n719, Z => n303);
   U1068 : MUX2DL port map( A0 => operand_regs_28_port, A1 => 
                           coeff_memory_4_28_port, SL => n712, Z => N3069);
   U1069 : MUX2DL port map( A0 => operand_regs_60_port, A1 => 
                           coeff_memory_3_28_port, SL => n710, Z => N3037);
   U1070 : MUX2DL port map( A0 => operand_regs_124_port, A1 => 
                           coeff_memory_2_28_port, SL => n717, Z => N3005);
   U1071 : MUX2DL port map( A0 => operand_regs_188_port, A1 => 
                           coeff_memory_1_28_port, SL => n716, Z => N2973);
   U1072 : MUX2DL port map( A0 => operand_regs_252_port, A1 => 
                           coeff_memory_0_28_port, SL => n714, Z => N2941);
   U1073 : NOR2D1 port map( A1 => avs_addr(5), A2 => avs_addr(4), Z => n114);
   U1074 : INVD1 port map( A => operand_regs_219_port, Z => n734);
   U1075 : INVD1 port map( A => avs_addr(0), Z => n762);
   U1076 : AND2D1 port map( A1 => avs_addr(2), A2 => n796, Z => n111);
   U1077 : INVD1 port map( A => avs_addr(1), Z => n796);
   U1078 : AND2D1 port map( A1 => n111, A2 => avs_addr(0), Z => n304);
   U1079 : MUX2DL port map( A0 => operand_regs_28_port, A1 => 
                           operand_regs_220_port, SL => n720, Z => n305);
   U1080 : AND3D1 port map( A1 => avs_addr(0), A2 => avs_addr(1), A3 => n547, Z
                           => n306);
   U1081 : AND3D1 port map( A1 => avs_addr(1), A2 => n547, A3 => n762, Z => 
                           n307);
   U1082 : AND3D1 port map( A1 => avs_addr(0), A2 => n796, A3 => n547, Z => 
                           n308);
   U1083 : AND2D1 port map( A1 => avs_addr(2), A2 => avs_addr(1), Z => n309);
   U1084 : MUX2DL port map( A0 => operand_regs_29_port, A1 => 
                           coeff_memory_4_29_port, SL => n712, Z => N3070);
   U1085 : MUX2DL port map( A0 => operand_regs_61_port, A1 => 
                           coeff_memory_3_29_port, SL => n710, Z => N3038);
   U1086 : MUX2DL port map( A0 => operand_regs_125_port, A1 => 
                           coeff_memory_2_29_port, SL => n718, Z => N3006);
   U1087 : MUX2DL port map( A0 => operand_regs_189_port, A1 => 
                           coeff_memory_1_29_port, SL => n716, Z => N2974);
   U1088 : MUX2DL port map( A0 => operand_regs_253_port, A1 => 
                           coeff_memory_0_29_port, SL => n714, Z => N2942);
   U1089 : INVD1 port map( A => operand_regs_220_port, Z => n733);
   U1090 : NOR2D1 port map( A1 => n92, A2 => n799, Z => n240);
   U1091 : NOR2D1 port map( A1 => n95, A2 => n799, Z => n241);
   U1092 : NAN3D1 port map( A1 => avs_write, A2 => n795, A3 => n304, Z => n179)
                           ;
   U1093 : MUX2DL port map( A0 => operand_regs_29_port, A1 => 
                           operand_regs_221_port, SL => n719, Z => n310);
   U1094 : AO31D1 port map( A1 => avs_write, A2 => n795, A3 => n276, B => 
                           stop_sim_port, Z => n157);
   U1095 : MUX2DL port map( A0 => operand_regs_30_port, A1 => 
                           coeff_memory_4_30_port, SL => n712, Z => N3071);
   U1096 : MUX2DL port map( A0 => operand_regs_62_port, A1 => 
                           coeff_memory_3_30_port, SL => n710, Z => N3039);
   U1097 : MUX2DL port map( A0 => operand_regs_126_port, A1 => 
                           coeff_memory_2_30_port, SL => n717, Z => N3007);
   U1098 : MUX2DL port map( A0 => operand_regs_190_port, A1 => 
                           coeff_memory_1_30_port, SL => n716, Z => N2975);
   U1099 : MUX2DL port map( A0 => operand_regs_254_port, A1 => 
                           coeff_memory_0_30_port, SL => n716, Z => N2943);
   U1100 : MUX2DL port map( A0 => operand_regs_30_port, A1 => 
                           operand_regs_222_port, SL => n720, Z => n311);
   U1101 : INVD1 port map( A => operand_regs_223_port, Z => n730);
   U1102 : INVD1 port map( A => operand_regs_221_port, Z => n732);
   U1103 : INVD1 port map( A => operand_regs_222_port, Z => n731);
   U1104 : MUX2DL port map( A0 => operand_regs_31_port, A1 => 
                           coeff_memory_4_31_port, SL => n712, Z => N3072);
   U1105 : MUX2DL port map( A0 => operand_regs_63_port, A1 => 
                           coeff_memory_3_31_port, SL => n710, Z => N3040);
   U1106 : MUX2DL port map( A0 => operand_regs_255_port, A1 => 
                           coeff_memory_0_31_port, SL => n712, Z => N2944);
   U1107 : MUX2DL port map( A0 => operand_regs_127_port, A1 => 
                           coeff_memory_2_31_port, SL => n718, Z => N3008);
   U1108 : MUX2DL port map( A0 => operand_regs_191_port, A1 => 
                           coeff_memory_1_31_port, SL => n716, Z => N2976);
   U1109 : MUX2DL port map( A0 => operand_regs_31_port, A1 => 
                           operand_regs_223_port, SL => n719, Z => n312);
   U1110 : AO22D1 port map( A1 => N2876, A2 => n697, B1 => N2859, B2 => n812, Z
                           => N2894);
   U1111 : AO22D1 port map( A1 => N2875, A2 => n697, B1 => N2858, B2 => n812, Z
                           => N2895);
   U1112 : AO22D1 port map( A1 => N2874, A2 => n697, B1 => N2857, B2 => n812, Z
                           => N2896);
   U1113 : AO22D1 port map( A1 => N2873, A2 => n697, B1 => N2856, B2 => n812, Z
                           => N2897);
   U1114 : AO22D1 port map( A1 => N2872, A2 => n697, B1 => N2855, B2 => n812, Z
                           => N2898);
   U1115 : AO22D1 port map( A1 => N2871, A2 => n697, B1 => N2854, B2 => n812, Z
                           => N2899);
   U1116 : AO22D1 port map( A1 => N2870, A2 => n697, B1 => N2853, B2 => n812, Z
                           => N2900);
   U1117 : AO22D1 port map( A1 => N2869, A2 => n697, B1 => N2852, B2 => n812, Z
                           => N2901);
   U1118 : AO22D1 port map( A1 => N2868, A2 => n697, B1 => N2851, B2 => n812, Z
                           => N2902);
   U1119 : AO22D1 port map( A1 => N2867, A2 => n697, B1 => N2850, B2 => n812, Z
                           => N2903);
   U1120 : AO22D1 port map( A1 => N2881, A2 => n697, B1 => N2864, B2 => n812, Z
                           => N2889);
   U1121 : AO22D1 port map( A1 => N2880, A2 => n697, B1 => N2863, B2 => n812, Z
                           => N2890);
   U1122 : AO22D1 port map( A1 => N2879, A2 => n697, B1 => N2862, B2 => n812, Z
                           => N2891);
   U1123 : AO22D1 port map( A1 => N2878, A2 => n697, B1 => N2861, B2 => n812, Z
                           => N2892);
   U1124 : AO22D1 port map( A1 => N2877, A2 => n697, B1 => N2860, B2 => n812, Z
                           => N2893);
   U1125 : AO22D1 port map( A1 => N2882, A2 => n697, B1 => N2865, B2 => n812, Z
                           => N2888);
   U1126 : INVD1 port map( A => N64, Z => n696);
   U1127 : NOR2D1 port map( A1 => n801, A2 => out_busy, Z => n79);
   U1128 : NAN3D1 port map( A1 => n81, A2 => out_busy, A3 => N62, Z => n4);
   U1129 : INVD1 port map( A => N62, Z => n810);
   U1130 : BUFD1 port map( A => odd1, Z => n697);
   U1131 : INVD1 port map( A => out_busy, Z => n811);
   U1132 : INVD1 port map( A => odd, Z => n803);
   U1133 : NAN3D1 port map( A1 => in_counter_1_port, A2 => in_busy, A3 => 
                           in_counter_0_port, Z => n88);
   U1134 : NOR2D1 port map( A1 => n806, A2 => in_counter_0_port, Z => n155);
   U1135 : OAI21M20D1 port map( A1 => n806, A2 => in_trigger, B => n100, Z => 
                           n84);
   U1136 : INVD1 port map( A => in_busy, Z => n806);
   U1137 : INVD1 port map( A => in_counter_2_port, Z => n809);
   U1138 : INVD1 port map( A => N63, Z => n813);
   U1139 : NOR2D1 port map( A1 => n804, A2 => in_counter_1_port, Z => n119);
   U1140 : NAN2D1 port map( A1 => in_counter_1_port, A2 => n155, Z => n85);
   U1141 : AND3D1 port map( A1 => in_counter_0_port, A2 => in_busy, A3 => n808,
                           Z => n87);
   U1142 : INVD1 port map( A => in_counter_1_port, Z => n808);
   U1143 : NAN2D1 port map( A1 => n78, A2 => n697, Z => n77);
   U1144 : NOR2D1 port map( A1 => n803, A2 => in_counter_2_port, Z => n101);
   U1145 : NOR2D1 port map( A1 => n809, A2 => odd, Z => n115);
   U1146 : NOR2D1 port map( A1 => odd, A2 => in_counter_2_port, Z => n120);
   U1147 : INVD1 port map( A => out_trigger, Z => n802);
   U1148 : NOR2D1 port map( A1 => n547, A2 => avs_addr(1), Z => n313);
   U1149 : NOR2D1 port map( A1 => n547, A2 => n796, Z => n314);
   U1150 : AOI22D1 port map( A1 => in_buf_64_port, A2 => n243, B1 => 
                           in_buf_0_port, B2 => n262, Z => n320);
   U1151 : NOR2D1 port map( A1 => avs_addr(1), A2 => avs_addr(2), Z => n315);
   U1152 : AND2D1 port map( A1 => n315, A2 => avs_addr(0), Z => n539);
   U1153 : NOR2D1 port map( A1 => n796, A2 => avs_addr(2), Z => n316);
   U1154 : AND2D1 port map( A1 => n316, A2 => avs_addr(0), Z => n538);
   U1155 : AOI22D1 port map( A1 => in_buf_192_port, A2 => n552, B1 => 
                           in_buf_128_port, B2 => n550, Z => n319);
   U1156 : NOR2M1D1 port map( A1 => n313, A2 => avs_addr(0), Z => n541);
   U1157 : NOR2M1D1 port map( A1 => n314, A2 => avs_addr(0), Z => n540);
   U1158 : AOI22D1 port map( A1 => in_buf_96_port, A2 => n554, B1 => 
                           in_buf_32_port, B2 => n540, Z => n318);
   U1159 : NOR2M1D1 port map( A1 => n315, A2 => avs_addr(0), Z => n543);
   U1160 : NOR2M1D1 port map( A1 => n316, A2 => avs_addr(0), Z => n542);
   U1161 : AOI22D1 port map( A1 => in_buf_224_port, A2 => n559, B1 => 
                           in_buf_160_port, B2 => n557, Z => n317);
   U1162 : NAN4D1 port map( A1 => n320, A2 => n319, A3 => n318, A4 => n317, Z 
                           => N2041);
   U1163 : AOI22D1 port map( A1 => in_buf_65_port, A2 => n243, B1 => 
                           in_buf_1_port, B2 => n262, Z => n324);
   U1164 : AOI22D1 port map( A1 => in_buf_193_port, A2 => n539, B1 => 
                           in_buf_129_port, B2 => n538, Z => n323);
   U1165 : AOI22D1 port map( A1 => in_buf_97_port, A2 => n554, B1 => 
                           in_buf_33_port, B2 => n540, Z => n322);
   U1166 : AOI22D1 port map( A1 => in_buf_225_port, A2 => n543, B1 => 
                           in_buf_161_port, B2 => n542, Z => n321);
   U1167 : NAN4D1 port map( A1 => n324, A2 => n323, A3 => n322, A4 => n321, Z 
                           => N2040);
   U1168 : AOI22D1 port map( A1 => in_buf_66_port, A2 => n243, B1 => 
                           in_buf_2_port, B2 => n262, Z => n328);
   U1169 : AOI22D1 port map( A1 => in_buf_194_port, A2 => n539, B1 => 
                           in_buf_130_port, B2 => n538, Z => n327);
   U1170 : AOI22D1 port map( A1 => in_buf_98_port, A2 => n554, B1 => 
                           in_buf_34_port, B2 => n540, Z => n326);
   U1171 : AOI22D1 port map( A1 => in_buf_226_port, A2 => n543, B1 => 
                           in_buf_162_port, B2 => n542, Z => n325);
   U1172 : NAN4D1 port map( A1 => n328, A2 => n327, A3 => n326, A4 => n325, Z 
                           => N2039);
   U1173 : AOI22D1 port map( A1 => in_buf_67_port, A2 => n243, B1 => 
                           in_buf_3_port, B2 => n262, Z => n332);
   U1174 : AOI22D1 port map( A1 => in_buf_195_port, A2 => n539, B1 => 
                           in_buf_131_port, B2 => n538, Z => n331);
   U1175 : AOI22D1 port map( A1 => in_buf_99_port, A2 => n554, B1 => 
                           in_buf_35_port, B2 => n540, Z => n330);
   U1176 : AOI22D1 port map( A1 => in_buf_227_port, A2 => n543, B1 => 
                           in_buf_163_port, B2 => n542, Z => n329);
   U1177 : NAN4D1 port map( A1 => n332, A2 => n331, A3 => n330, A4 => n329, Z 
                           => N2038);
   U1178 : AOI22D1 port map( A1 => in_buf_68_port, A2 => n243, B1 => 
                           in_buf_4_port, B2 => n262, Z => n336);
   U1179 : AOI22D1 port map( A1 => in_buf_196_port, A2 => n539, B1 => 
                           in_buf_132_port, B2 => n538, Z => n335);
   U1180 : AOI22D1 port map( A1 => in_buf_100_port, A2 => n554, B1 => 
                           in_buf_36_port, B2 => n540, Z => n334);
   U1181 : AOI22D1 port map( A1 => in_buf_228_port, A2 => n543, B1 => 
                           in_buf_164_port, B2 => n542, Z => n333);
   U1182 : NAN4D1 port map( A1 => n336, A2 => n335, A3 => n334, A4 => n333, Z 
                           => N2037);
   U1183 : AOI22D1 port map( A1 => in_buf_69_port, A2 => n243, B1 => 
                           in_buf_5_port, B2 => n262, Z => n340);
   U1184 : AOI22D1 port map( A1 => in_buf_197_port, A2 => n539, B1 => 
                           in_buf_133_port, B2 => n538, Z => n339);
   U1185 : AOI22D1 port map( A1 => in_buf_101_port, A2 => n554, B1 => 
                           in_buf_37_port, B2 => n540, Z => n338);
   U1186 : AOI22D1 port map( A1 => in_buf_229_port, A2 => n543, B1 => 
                           in_buf_165_port, B2 => n542, Z => n337);
   U1187 : NAN4D1 port map( A1 => n340, A2 => n339, A3 => n338, A4 => n337, Z 
                           => N2036);
   U1188 : AOI22D1 port map( A1 => in_buf_70_port, A2 => n243, B1 => 
                           in_buf_6_port, B2 => n262, Z => n344);
   U1189 : AOI22D1 port map( A1 => in_buf_198_port, A2 => n539, B1 => 
                           in_buf_134_port, B2 => n538, Z => n343);
   U1190 : AOI22D1 port map( A1 => in_buf_102_port, A2 => n554, B1 => 
                           in_buf_38_port, B2 => n540, Z => n342);
   U1191 : AOI22D1 port map( A1 => in_buf_230_port, A2 => n543, B1 => 
                           in_buf_166_port, B2 => n542, Z => n341);
   U1192 : NAN4D1 port map( A1 => n344, A2 => n343, A3 => n342, A4 => n341, Z 
                           => N2035);
   U1193 : AOI22D1 port map( A1 => in_buf_71_port, A2 => n243, B1 => 
                           in_buf_7_port, B2 => n262, Z => n348);
   U1194 : AOI22D1 port map( A1 => in_buf_199_port, A2 => n539, B1 => 
                           in_buf_135_port, B2 => n538, Z => n347);
   U1195 : AOI22D1 port map( A1 => in_buf_103_port, A2 => n554, B1 => 
                           in_buf_39_port, B2 => n540, Z => n346);
   U1196 : AOI22D1 port map( A1 => in_buf_231_port, A2 => n543, B1 => 
                           in_buf_167_port, B2 => n542, Z => n345);
   U1197 : NAN4D1 port map( A1 => n348, A2 => n347, A3 => n346, A4 => n345, Z 
                           => N2034);
   U1198 : AOI22D1 port map( A1 => in_buf_72_port, A2 => n243, B1 => 
                           in_buf_8_port, B2 => n262, Z => n352);
   U1199 : AOI22D1 port map( A1 => in_buf_200_port, A2 => n539, B1 => 
                           in_buf_136_port, B2 => n538, Z => n351);
   U1200 : AOI22D1 port map( A1 => in_buf_104_port, A2 => n541, B1 => 
                           in_buf_40_port, B2 => n540, Z => n350);
   U1201 : AOI22D1 port map( A1 => in_buf_232_port, A2 => n543, B1 => 
                           in_buf_168_port, B2 => n542, Z => n349);
   U1202 : NAN4D1 port map( A1 => n352, A2 => n351, A3 => n350, A4 => n349, Z 
                           => N2033);
   U1203 : AOI22D1 port map( A1 => in_buf_73_port, A2 => n243, B1 => 
                           in_buf_9_port, B2 => n262, Z => n356);
   U1204 : AOI22D1 port map( A1 => in_buf_201_port, A2 => n539, B1 => 
                           in_buf_137_port, B2 => n538, Z => n355);
   U1205 : AOI22D1 port map( A1 => in_buf_105_port, A2 => n541, B1 => 
                           in_buf_41_port, B2 => n540, Z => n354);
   U1206 : AOI22D1 port map( A1 => in_buf_233_port, A2 => n543, B1 => 
                           in_buf_169_port, B2 => n542, Z => n353);
   U1207 : NAN4D1 port map( A1 => n356, A2 => n355, A3 => n354, A4 => n353, Z 
                           => N2032);
   U1208 : AOI22D1 port map( A1 => in_buf_74_port, A2 => n243, B1 => 
                           in_buf_10_port, B2 => n262, Z => n360);
   U1209 : AOI22D1 port map( A1 => in_buf_202_port, A2 => n539, B1 => 
                           in_buf_138_port, B2 => n538, Z => n359);
   U1210 : AOI22D1 port map( A1 => in_buf_106_port, A2 => n541, B1 => 
                           in_buf_42_port, B2 => n540, Z => n358);
   U1211 : AOI22D1 port map( A1 => in_buf_234_port, A2 => n559, B1 => 
                           in_buf_170_port, B2 => n542, Z => n357);
   U1212 : NAN4D1 port map( A1 => n360, A2 => n359, A3 => n358, A4 => n357, Z 
                           => N2031);
   U1213 : AOI22D1 port map( A1 => in_buf_75_port, A2 => n243, B1 => 
                           in_buf_11_port, B2 => n262, Z => n364);
   U1214 : AOI22D1 port map( A1 => in_buf_203_port, A2 => n539, B1 => 
                           in_buf_139_port, B2 => n538, Z => n363);
   U1215 : AOI22D1 port map( A1 => in_buf_107_port, A2 => n541, B1 => 
                           in_buf_43_port, B2 => n540, Z => n362);
   U1216 : AOI22D1 port map( A1 => in_buf_235_port, A2 => n543, B1 => 
                           in_buf_171_port, B2 => n542, Z => n361);
   U1217 : NAN4D1 port map( A1 => n364, A2 => n363, A3 => n362, A4 => n361, Z 
                           => N2030);
   U1218 : AOI22D1 port map( A1 => in_buf_76_port, A2 => n243, B1 => 
                           in_buf_12_port, B2 => n262, Z => n368);
   U1219 : AOI22D1 port map( A1 => in_buf_204_port, A2 => n539, B1 => 
                           in_buf_140_port, B2 => n538, Z => n367);
   U1220 : AOI22D1 port map( A1 => in_buf_108_port, A2 => n554, B1 => 
                           in_buf_44_port, B2 => n540, Z => n366);
   U1221 : AOI22D1 port map( A1 => in_buf_236_port, A2 => n559, B1 => 
                           in_buf_172_port, B2 => n557, Z => n365);
   U1222 : NAN4D1 port map( A1 => n368, A2 => n367, A3 => n366, A4 => n365, Z 
                           => N2029);
   U1223 : AOI22D1 port map( A1 => in_buf_77_port, A2 => n243, B1 => 
                           in_buf_13_port, B2 => n262, Z => n372);
   U1224 : AOI22D1 port map( A1 => in_buf_205_port, A2 => n552, B1 => 
                           in_buf_141_port, B2 => n550, Z => n371);
   U1225 : AOI22D1 port map( A1 => in_buf_109_port, A2 => n541, B1 => 
                           in_buf_45_port, B2 => n540, Z => n370);
   U1226 : AOI22D1 port map( A1 => in_buf_237_port, A2 => n559, B1 => 
                           in_buf_173_port, B2 => n556, Z => n369);
   U1227 : NAN4D1 port map( A1 => n372, A2 => n371, A3 => n370, A4 => n369, Z 
                           => N2028);
   U1228 : AOI22D1 port map( A1 => in_buf_78_port, A2 => n243, B1 => 
                           in_buf_14_port, B2 => n262, Z => n376);
   U1229 : AOI22D1 port map( A1 => in_buf_206_port, A2 => n552, B1 => 
                           in_buf_142_port, B2 => n550, Z => n375);
   U1230 : AOI22D1 port map( A1 => in_buf_110_port, A2 => n541, B1 => 
                           in_buf_46_port, B2 => n540, Z => n374);
   U1231 : AOI22D1 port map( A1 => in_buf_238_port, A2 => n559, B1 => 
                           in_buf_174_port, B2 => n542, Z => n373);
   U1232 : NAN4D1 port map( A1 => n376, A2 => n375, A3 => n374, A4 => n373, Z 
                           => N2027);
   U1233 : AOI22D1 port map( A1 => in_buf_79_port, A2 => n243, B1 => 
                           in_buf_15_port, B2 => n262, Z => n380);
   U1234 : AOI22D1 port map( A1 => in_buf_207_port, A2 => n552, B1 => 
                           in_buf_143_port, B2 => n550, Z => n379);
   U1235 : AOI22D1 port map( A1 => in_buf_111_port, A2 => n541, B1 => 
                           in_buf_47_port, B2 => n540, Z => n378);
   U1236 : AOI22D1 port map( A1 => in_buf_239_port, A2 => n559, B1 => 
                           in_buf_175_port, B2 => n542, Z => n377);
   U1237 : NAN4D1 port map( A1 => n380, A2 => n379, A3 => n378, A4 => n377, Z 
                           => N2026);
   U1238 : AOI22D1 port map( A1 => in_buf_80_port, A2 => n243, B1 => 
                           in_buf_16_port, B2 => n262, Z => n384);
   U1239 : AOI22D1 port map( A1 => in_buf_208_port, A2 => n552, B1 => 
                           in_buf_144_port, B2 => n550, Z => n383);
   U1240 : AOI22D1 port map( A1 => in_buf_112_port, A2 => n541, B1 => 
                           in_buf_48_port, B2 => n540, Z => n382);
   U1241 : AOI22D1 port map( A1 => in_buf_240_port, A2 => n559, B1 => 
                           in_buf_176_port, B2 => n542, Z => n381);
   U1242 : NAN4D1 port map( A1 => n384, A2 => n383, A3 => n382, A4 => n381, Z 
                           => N2025);
   U1243 : AOI22D1 port map( A1 => in_buf_81_port, A2 => n243, B1 => 
                           in_buf_17_port, B2 => n262, Z => n388);
   U1244 : AOI22D1 port map( A1 => in_buf_209_port, A2 => n552, B1 => 
                           in_buf_145_port, B2 => n550, Z => n387);
   U1245 : AOI22D1 port map( A1 => in_buf_113_port, A2 => n541, B1 => 
                           in_buf_49_port, B2 => n540, Z => n386);
   U1246 : AOI22D1 port map( A1 => in_buf_241_port, A2 => n559, B1 => 
                           in_buf_177_port, B2 => n542, Z => n385);
   U1247 : NAN4D1 port map( A1 => n388, A2 => n387, A3 => n386, A4 => n385, Z 
                           => N2024);
   U1248 : AOI22D1 port map( A1 => in_buf_82_port, A2 => n243, B1 => 
                           in_buf_18_port, B2 => n262, Z => n392);
   U1249 : AOI22D1 port map( A1 => in_buf_210_port, A2 => n552, B1 => 
                           in_buf_146_port, B2 => n550, Z => n391);
   U1250 : AOI22D1 port map( A1 => in_buf_114_port, A2 => n541, B1 => 
                           in_buf_50_port, B2 => n540, Z => n390);
   U1251 : AOI22D1 port map( A1 => in_buf_242_port, A2 => n559, B1 => 
                           in_buf_178_port, B2 => n542, Z => n389);
   U1252 : NAN4D1 port map( A1 => n392, A2 => n391, A3 => n390, A4 => n389, Z 
                           => N2023);
   U1253 : AOI22D1 port map( A1 => in_buf_83_port, A2 => n243, B1 => 
                           in_buf_19_port, B2 => n262, Z => n396);
   U1254 : AOI22D1 port map( A1 => in_buf_211_port, A2 => n552, B1 => 
                           in_buf_147_port, B2 => n550, Z => n395);
   U1255 : AOI22D1 port map( A1 => in_buf_115_port, A2 => n541, B1 => 
                           in_buf_51_port, B2 => n540, Z => n394);
   U1256 : AOI22D1 port map( A1 => in_buf_243_port, A2 => n559, B1 => 
                           in_buf_179_port, B2 => n542, Z => n393);
   U1257 : NAN4D1 port map( A1 => n396, A2 => n395, A3 => n394, A4 => n393, Z 
                           => N2022);
   U1258 : AOI22D1 port map( A1 => in_buf_84_port, A2 => n243, B1 => 
                           in_buf_20_port, B2 => n262, Z => n400);
   U1259 : AOI22D1 port map( A1 => in_buf_212_port, A2 => n552, B1 => 
                           in_buf_148_port, B2 => n550, Z => n399);
   U1260 : AOI22D1 port map( A1 => in_buf_116_port, A2 => n541, B1 => 
                           in_buf_52_port, B2 => n540, Z => n398);
   U1261 : AOI22D1 port map( A1 => in_buf_244_port, A2 => n559, B1 => 
                           in_buf_180_port, B2 => n542, Z => n397);
   U1262 : NAN4D1 port map( A1 => n400, A2 => n399, A3 => n398, A4 => n397, Z 
                           => N2021);
   U1263 : AOI22D1 port map( A1 => in_buf_85_port, A2 => n243, B1 => 
                           in_buf_21_port, B2 => n262, Z => n404);
   U1264 : AOI22D1 port map( A1 => in_buf_213_port, A2 => n552, B1 => 
                           in_buf_149_port, B2 => n550, Z => n403);
   U1265 : AOI22D1 port map( A1 => in_buf_117_port, A2 => n541, B1 => 
                           in_buf_53_port, B2 => n540, Z => n402);
   U1266 : AOI22D1 port map( A1 => in_buf_245_port, A2 => n559, B1 => 
                           in_buf_181_port, B2 => n542, Z => n401);
   U1267 : NAN4D1 port map( A1 => n404, A2 => n403, A3 => n402, A4 => n401, Z 
                           => N2020);
   U1268 : AOI22D1 port map( A1 => in_buf_86_port, A2 => n243, B1 => 
                           in_buf_22_port, B2 => n262, Z => n408);
   U1269 : AOI22D1 port map( A1 => in_buf_214_port, A2 => n552, B1 => 
                           in_buf_150_port, B2 => n550, Z => n407);
   U1270 : AOI22D1 port map( A1 => in_buf_118_port, A2 => n541, B1 => 
                           in_buf_54_port, B2 => n540, Z => n406);
   U1271 : AOI22D1 port map( A1 => in_buf_246_port, A2 => n559, B1 => 
                           in_buf_182_port, B2 => n542, Z => n405);
   U1272 : NAN4D1 port map( A1 => n408, A2 => n407, A3 => n406, A4 => n405, Z 
                           => N2019);
   U1273 : AOI22D1 port map( A1 => in_buf_87_port, A2 => n243, B1 => 
                           in_buf_23_port, B2 => n262, Z => n412);
   U1274 : AOI22D1 port map( A1 => in_buf_215_port, A2 => n552, B1 => 
                           in_buf_151_port, B2 => n550, Z => n411);
   U1275 : AOI22D1 port map( A1 => in_buf_119_port, A2 => n541, B1 => 
                           in_buf_55_port, B2 => n540, Z => n410);
   U1276 : AOI22D1 port map( A1 => in_buf_247_port, A2 => n559, B1 => 
                           in_buf_183_port, B2 => n542, Z => n409);
   U1277 : NAN4D1 port map( A1 => n412, A2 => n411, A3 => n410, A4 => n409, Z 
                           => N2018);
   U1278 : AOI22D1 port map( A1 => in_buf_88_port, A2 => n243, B1 => 
                           in_buf_24_port, B2 => n262, Z => n416);
   U1279 : AOI22D1 port map( A1 => in_buf_216_port, A2 => n552, B1 => 
                           in_buf_152_port, B2 => n550, Z => n415);
   U1280 : AOI22D1 port map( A1 => in_buf_120_port, A2 => n541, B1 => 
                           in_buf_56_port, B2 => n540, Z => n414);
   U1281 : AOI22D1 port map( A1 => in_buf_248_port, A2 => n559, B1 => 
                           in_buf_184_port, B2 => n542, Z => n413);
   U1282 : NAN4D1 port map( A1 => n416, A2 => n415, A3 => n414, A4 => n413, Z 
                           => N2017);
   U1283 : AOI22D1 port map( A1 => in_buf_89_port, A2 => n243, B1 => 
                           in_buf_25_port, B2 => n262, Z => n420);
   U1284 : AOI22D1 port map( A1 => in_buf_217_port, A2 => n552, B1 => 
                           in_buf_153_port, B2 => n550, Z => n419);
   U1285 : AOI22D1 port map( A1 => in_buf_121_port, A2 => n541, B1 => 
                           in_buf_57_port, B2 => n540, Z => n418);
   U1286 : AOI22D1 port map( A1 => in_buf_249_port, A2 => n559, B1 => 
                           in_buf_185_port, B2 => n556, Z => n417);
   U1287 : NAN4D1 port map( A1 => n420, A2 => n419, A3 => n418, A4 => n417, Z 
                           => N2016);
   U1288 : AOI22D1 port map( A1 => in_buf_90_port, A2 => n243, B1 => 
                           in_buf_26_port, B2 => n262, Z => n424);
   U1289 : AOI22D1 port map( A1 => in_buf_218_port, A2 => n552, B1 => 
                           in_buf_154_port, B2 => n549, Z => n423);
   U1290 : AOI22D1 port map( A1 => in_buf_122_port, A2 => n541, B1 => 
                           in_buf_58_port, B2 => n540, Z => n422);
   U1291 : AOI22D1 port map( A1 => in_buf_250_port, A2 => n543, B1 => 
                           in_buf_186_port, B2 => n557, Z => n421);
   U1292 : NAN4D1 port map( A1 => n424, A2 => n423, A3 => n422, A4 => n421, Z 
                           => N2015);
   U1293 : AOI22D1 port map( A1 => in_buf_91_port, A2 => n243, B1 => 
                           in_buf_27_port, B2 => n262, Z => n428);
   U1294 : AOI22D1 port map( A1 => in_buf_219_port, A2 => n539, B1 => 
                           in_buf_155_port, B2 => n549, Z => n427);
   U1295 : AOI22D1 port map( A1 => in_buf_123_port, A2 => n541, B1 => 
                           in_buf_59_port, B2 => n540, Z => n426);
   U1296 : AOI22D1 port map( A1 => in_buf_251_port, A2 => n543, B1 => 
                           in_buf_187_port, B2 => n557, Z => n425);
   U1297 : NAN4D1 port map( A1 => n428, A2 => n427, A3 => n426, A4 => n425, Z 
                           => N2014);
   U1298 : AOI22D1 port map( A1 => in_buf_92_port, A2 => n243, B1 => 
                           in_buf_28_port, B2 => n262, Z => n432);
   U1299 : AOI22D1 port map( A1 => in_buf_220_port, A2 => n539, B1 => 
                           in_buf_156_port, B2 => n549, Z => n431);
   U1300 : AOI22D1 port map( A1 => in_buf_124_port, A2 => n541, B1 => 
                           in_buf_60_port, B2 => n540, Z => n430);
   U1301 : AOI22D1 port map( A1 => in_buf_252_port, A2 => n543, B1 => 
                           in_buf_188_port, B2 => n557, Z => n429);
   U1302 : NAN4D1 port map( A1 => n432, A2 => n431, A3 => n430, A4 => n429, Z 
                           => N2013);
   U1303 : AOI22D1 port map( A1 => in_buf_93_port, A2 => n243, B1 => 
                           in_buf_29_port, B2 => n262, Z => n436);
   U1304 : AOI22D1 port map( A1 => in_buf_221_port, A2 => n539, B1 => 
                           in_buf_157_port, B2 => n549, Z => n435);
   U1305 : AOI22D1 port map( A1 => in_buf_125_port, A2 => n541, B1 => 
                           in_buf_61_port, B2 => n540, Z => n434);
   U1306 : AOI22D1 port map( A1 => in_buf_253_port, A2 => n543, B1 => 
                           in_buf_189_port, B2 => n557, Z => n433);
   U1307 : NAN4D1 port map( A1 => n436, A2 => n435, A3 => n434, A4 => n433, Z 
                           => N2012);
   U1308 : AOI22D1 port map( A1 => in_buf_94_port, A2 => n243, B1 => 
                           in_buf_30_port, B2 => n262, Z => n440);
   U1309 : AOI22D1 port map( A1 => in_buf_222_port, A2 => n552, B1 => 
                           in_buf_158_port, B2 => n549, Z => n439);
   U1310 : AOI22D1 port map( A1 => in_buf_126_port, A2 => n541, B1 => 
                           in_buf_62_port, B2 => n540, Z => n438);
   U1311 : AOI22D1 port map( A1 => in_buf_254_port, A2 => n559, B1 => 
                           in_buf_190_port, B2 => n557, Z => n437);
   U1312 : NAN4D1 port map( A1 => n440, A2 => n439, A3 => n438, A4 => n437, Z 
                           => N2011);
   U1313 : AOI22D1 port map( A1 => in_buf_95_port, A2 => n243, B1 => 
                           in_buf_31_port, B2 => n262, Z => n444);
   U1314 : AOI22D1 port map( A1 => in_buf_223_port, A2 => n539, B1 => 
                           in_buf_159_port, B2 => n549, Z => n443);
   U1315 : AOI22D1 port map( A1 => in_buf_255_port, A2 => n543, B1 => 
                           in_buf_191_port, B2 => n557, Z => n441);
   U1316 : NAN4D1 port map( A1 => n444, A2 => n443, A3 => n442, A4 => n441, Z 
                           => N2010);
   U1317 : AOI22D1 port map( A1 => comp_res_96_port, A2 => n539, B1 => 
                           comp_res_32_port, B2 => n549, Z => n447);
   U1318 : AOI22D1 port map( A1 => comp_res_128_port, A2 => n543, B1 => 
                           comp_res_64_port, B2 => n557, Z => n445);
   U1319 : AOI22D1 port map( A1 => comp_res_97_port, A2 => n539, B1 => 
                           comp_res_33_port, B2 => n549, Z => n450);
   U1320 : AOI22D1 port map( A1 => comp_res_129_port, A2 => n543, B1 => 
                           comp_res_65_port, B2 => n557, Z => n448);
   U1321 : AOI22D1 port map( A1 => comp_res_98_port, A2 => n539, B1 => 
                           comp_res_34_port, B2 => n549, Z => n453);
   U1322 : AOI22D1 port map( A1 => comp_res_130_port, A2 => n543, B1 => 
                           comp_res_66_port, B2 => n557, Z => n451);
   U1323 : AOI22D1 port map( A1 => comp_res_99_port, A2 => n539, B1 => 
                           comp_res_35_port, B2 => n549, Z => n456);
   U1324 : AOI22D1 port map( A1 => comp_res_131_port, A2 => n543, B1 => 
                           comp_res_67_port, B2 => n557, Z => n454);
   U1325 : AOI22D1 port map( A1 => comp_res_100_port, A2 => n539, B1 => 
                           comp_res_36_port, B2 => n549, Z => n459);
   U1326 : AOI22D1 port map( A1 => comp_res_132_port, A2 => n543, B1 => 
                           comp_res_68_port, B2 => n557, Z => n457);
   U1327 : AOI22D1 port map( A1 => comp_res_101_port, A2 => n539, B1 => 
                           comp_res_37_port, B2 => n549, Z => n462);
   U1328 : AOI22D1 port map( A1 => comp_res_133_port, A2 => n543, B1 => 
                           comp_res_69_port, B2 => n557, Z => n460);
   U1329 : AOI22D1 port map( A1 => comp_res_102_port, A2 => n539, B1 => 
                           comp_res_38_port, B2 => n549, Z => n465);
   U1330 : AOI22D1 port map( A1 => comp_res_134_port, A2 => n543, B1 => 
                           comp_res_70_port, B2 => n557, Z => n463);
   U1331 : AOI22D1 port map( A1 => comp_res_103_port, A2 => n539, B1 => 
                           comp_res_39_port, B2 => n550, Z => n468);
   U1332 : AOI22D1 port map( A1 => comp_res_135_port, A2 => n543, B1 => 
                           comp_res_71_port, B2 => n556, Z => n466);
   U1333 : AOI22D1 port map( A1 => comp_res_104_port, A2 => n539, B1 => 
                           comp_res_40_port, B2 => n538, Z => n471);
   U1334 : AOI22D1 port map( A1 => comp_res_136_port, A2 => n559, B1 => 
                           comp_res_72_port, B2 => n542, Z => n469);
   U1335 : AOI22D1 port map( A1 => comp_res_105_port, A2 => n539, B1 => 
                           comp_res_41_port, B2 => n550, Z => n474);
   U1336 : AOI22D1 port map( A1 => comp_res_137_port, A2 => n543, B1 => 
                           comp_res_73_port, B2 => n542, Z => n472);
   U1337 : AOI22D1 port map( A1 => comp_res_106_port, A2 => n539, B1 => 
                           comp_res_42_port, B2 => n549, Z => n477);
   U1338 : AOI22D1 port map( A1 => comp_res_138_port, A2 => n559, B1 => 
                           comp_res_74_port, B2 => n542, Z => n475);
   U1339 : AOI22D1 port map( A1 => comp_res_107_port, A2 => n552, B1 => 
                           comp_res_43_port, B2 => n538, Z => n480);
   U1340 : AOI22D1 port map( A1 => comp_res_139_port, A2 => n543, B1 => 
                           comp_res_75_port, B2 => n557, Z => n478);
   U1341 : AOI22D1 port map( A1 => comp_res_108_port, A2 => n539, B1 => 
                           comp_res_44_port, B2 => n550, Z => n483);
   U1342 : AOI22D1 port map( A1 => comp_res_140_port, A2 => n559, B1 => 
                           comp_res_76_port, B2 => n542, Z => n481);
   U1343 : AOI22D1 port map( A1 => comp_res_109_port, A2 => n539, B1 => 
                           comp_res_45_port, B2 => n549, Z => n486);
   U1344 : AOI22D1 port map( A1 => comp_res_141_port, A2 => n543, B1 => 
                           comp_res_77_port, B2 => n542, Z => n484);
   U1345 : AOI22D1 port map( A1 => comp_res_110_port, A2 => n539, B1 => 
                           comp_res_46_port, B2 => n538, Z => n489);
   U1346 : AOI22D1 port map( A1 => comp_res_142_port, A2 => n559, B1 => 
                           comp_res_78_port, B2 => n557, Z => n487);
   U1347 : AOI22D1 port map( A1 => comp_res_111_port, A2 => n539, B1 => 
                           comp_res_47_port, B2 => n549, Z => n492);
   U1348 : AOI22D1 port map( A1 => comp_res_143_port, A2 => n543, B1 => 
                           comp_res_79_port, B2 => n556, Z => n490);
   U1349 : AOI22D1 port map( A1 => comp_res_112_port, A2 => n539, B1 => 
                           comp_res_48_port, B2 => n538, Z => n495);
   U1350 : AOI22D1 port map( A1 => comp_res_144_port, A2 => n543, B1 => 
                           comp_res_80_port, B2 => n542, Z => n493);
   U1351 : AOI22D1 port map( A1 => comp_res_113_port, A2 => n539, B1 => 
                           comp_res_49_port, B2 => n538, Z => n498);
   U1352 : AOI22D1 port map( A1 => comp_res_145_port, A2 => n543, B1 => 
                           comp_res_81_port, B2 => n556, Z => n496);
   U1353 : AOI22D1 port map( A1 => comp_res_114_port, A2 => n539, B1 => 
                           comp_res_50_port, B2 => n549, Z => n501);
   U1354 : AOI22D1 port map( A1 => comp_res_146_port, A2 => n559, B1 => 
                           comp_res_82_port, B2 => n556, Z => n499);
   U1355 : AOI22D1 port map( A1 => comp_res_115_port, A2 => n539, B1 => 
                           comp_res_51_port, B2 => n549, Z => n504);
   U1356 : AOI22D1 port map( A1 => comp_res_147_port, A2 => n543, B1 => 
                           comp_res_83_port, B2 => n556, Z => n502);
   U1357 : AOI22D1 port map( A1 => comp_res_116_port, A2 => n539, B1 => 
                           comp_res_52_port, B2 => n538, Z => n507);
   U1358 : AOI22D1 port map( A1 => comp_res_148_port, A2 => n543, B1 => 
                           comp_res_84_port, B2 => n556, Z => n505);
   U1359 : AOI22D1 port map( A1 => comp_res_117_port, A2 => n539, B1 => 
                           comp_res_53_port, B2 => n538, Z => n510);
   U1360 : AOI22D1 port map( A1 => comp_res_149_port, A2 => n543, B1 => 
                           comp_res_85_port, B2 => n556, Z => n508);
   U1361 : AOI22D1 port map( A1 => comp_res_118_port, A2 => n539, B1 => 
                           comp_res_54_port, B2 => n538, Z => n513);
   U1362 : AOI22D1 port map( A1 => comp_res_150_port, A2 => n543, B1 => 
                           comp_res_86_port, B2 => n556, Z => n511);
   U1363 : AOI22D1 port map( A1 => comp_res_119_port, A2 => n539, B1 => 
                           comp_res_55_port, B2 => n538, Z => n516);
   U1364 : AOI22D1 port map( A1 => comp_res_151_port, A2 => n543, B1 => 
                           comp_res_87_port, B2 => n556, Z => n514);
   U1365 : AOI22D1 port map( A1 => comp_res_120_port, A2 => n539, B1 => 
                           comp_res_56_port, B2 => n538, Z => n519);
   U1366 : AOI22D1 port map( A1 => comp_res_152_port, A2 => n543, B1 => 
                           comp_res_88_port, B2 => n556, Z => n517);
   U1367 : AOI22D1 port map( A1 => comp_res_121_port, A2 => n539, B1 => 
                           comp_res_57_port, B2 => n538, Z => n522);
   U1368 : AOI22D1 port map( A1 => comp_res_153_port, A2 => n559, B1 => 
                           comp_res_89_port, B2 => n556, Z => n520);
   U1369 : AOI22D1 port map( A1 => comp_res_122_port, A2 => n539, B1 => 
                           comp_res_58_port, B2 => n538, Z => n525);
   U1370 : AOI22D1 port map( A1 => comp_res_154_port, A2 => n543, B1 => 
                           comp_res_90_port, B2 => n556, Z => n523);
   U1371 : AOI22D1 port map( A1 => comp_res_123_port, A2 => n552, B1 => 
                           comp_res_59_port, B2 => n538, Z => n528);
   U1372 : AOI22D1 port map( A1 => comp_res_155_port, A2 => n543, B1 => 
                           comp_res_91_port, B2 => n556, Z => n526);
   U1373 : AOI22D1 port map( A1 => comp_res_124_port, A2 => n539, B1 => 
                           comp_res_60_port, B2 => n538, Z => n531);
   U1374 : AOI22D1 port map( A1 => comp_res_156_port, A2 => n559, B1 => 
                           comp_res_92_port, B2 => n556, Z => n529);
   U1375 : AOI22D1 port map( A1 => comp_res_125_port, A2 => n539, B1 => 
                           comp_res_61_port, B2 => n538, Z => n534);
   U1376 : AOI22D1 port map( A1 => comp_res_157_port, A2 => n543, B1 => 
                           comp_res_93_port, B2 => n556, Z => n532);
   U1377 : AOI22D1 port map( A1 => comp_res_126_port, A2 => n539, B1 => 
                           comp_res_62_port, B2 => n538, Z => n537);
   U1378 : AOI22D1 port map( A1 => comp_res_158_port, A2 => n559, B1 => 
                           comp_res_94_port, B2 => n556, Z => n535);
   U1379 : AOI22D1 port map( A1 => comp_res_127_port, A2 => n539, B1 => 
                           comp_res_63_port, B2 => n550, Z => n546);
   U1380 : AOI22D1 port map( A1 => comp_res_159_port, A2 => n543, B1 => 
                           comp_res_95_port, B2 => n556, Z => n544);
   U1381 : NOR2D1 port map( A1 => n696, A2 => N63, Z => n560);
   U1382 : NOR2D1 port map( A1 => n696, A2 => n813, Z => n561);
   U1383 : AOI22D1 port map( A1 => out_buf_80_port, A2 => n269, B1 => 
                           out_buf_16_port, B2 => n244, Z => n567);
   U1384 : NOR2D1 port map( A1 => N63, A2 => N64, Z => n562);
   U1385 : NOR2D1 port map( A1 => n813, A2 => N64, Z => n563);
   U1386 : AOI22D1 port map( A1 => out_buf_208_port, A2 => n270, B1 => 
                           out_buf_144_port, B2 => n245, Z => n566);
   U1387 : NOR2M1D1 port map( A1 => n560, A2 => N62, Z => n689);
   U1388 : NOR2M1D1 port map( A1 => n561, A2 => N62, Z => n688);
   U1389 : AOI22D1 port map( A1 => out_buf_112_port, A2 => n689, B1 => 
                           out_buf_48_port, B2 => n688, Z => n565);
   U1390 : NOR2M1D1 port map( A1 => n562, A2 => N62, Z => n691);
   U1391 : NOR2M1D1 port map( A1 => n563, A2 => N62, Z => n690);
   U1392 : AOI22D1 port map( A1 => out_buf_240_port, A2 => n691, B1 => 
                           out_buf_176_port, B2 => n690, Z => n564);
   U1393 : NAN4D1 port map( A1 => n567, A2 => n566, A3 => n565, A4 => n564, Z 
                           => N2882);
   U1394 : AOI22D1 port map( A1 => out_buf_81_port, A2 => n269, B1 => 
                           out_buf_17_port, B2 => n244, Z => n571);
   U1395 : AOI22D1 port map( A1 => out_buf_209_port, A2 => n270, B1 => 
                           out_buf_145_port, B2 => n245, Z => n570);
   U1396 : AOI22D1 port map( A1 => out_buf_113_port, A2 => n689, B1 => 
                           out_buf_49_port, B2 => n688, Z => n569);
   U1397 : AOI22D1 port map( A1 => out_buf_241_port, A2 => n691, B1 => 
                           out_buf_177_port, B2 => n690, Z => n568);
   U1398 : NAN4D1 port map( A1 => n571, A2 => n570, A3 => n569, A4 => n568, Z 
                           => N2881);
   U1399 : AOI22D1 port map( A1 => out_buf_82_port, A2 => n269, B1 => 
                           out_buf_18_port, B2 => n244, Z => n575);
   U1400 : AOI22D1 port map( A1 => out_buf_210_port, A2 => n270, B1 => 
                           out_buf_146_port, B2 => n245, Z => n574);
   U1401 : AOI22D1 port map( A1 => out_buf_114_port, A2 => n689, B1 => 
                           out_buf_50_port, B2 => n688, Z => n573);
   U1402 : AOI22D1 port map( A1 => out_buf_242_port, A2 => n691, B1 => 
                           out_buf_178_port, B2 => n690, Z => n572);
   U1403 : NAN4D1 port map( A1 => n575, A2 => n574, A3 => n573, A4 => n572, Z 
                           => N2880);
   U1404 : AOI22D1 port map( A1 => out_buf_83_port, A2 => n269, B1 => 
                           out_buf_19_port, B2 => n244, Z => n579);
   U1405 : AOI22D1 port map( A1 => out_buf_211_port, A2 => n270, B1 => 
                           out_buf_147_port, B2 => n245, Z => n578);
   U1406 : AOI22D1 port map( A1 => out_buf_115_port, A2 => n689, B1 => 
                           out_buf_51_port, B2 => n688, Z => n577);
   U1407 : AOI22D1 port map( A1 => out_buf_243_port, A2 => n691, B1 => 
                           out_buf_179_port, B2 => n690, Z => n576);
   U1408 : NAN4D1 port map( A1 => n579, A2 => n578, A3 => n577, A4 => n576, Z 
                           => N2879);
   U1409 : AOI22D1 port map( A1 => out_buf_84_port, A2 => n269, B1 => 
                           out_buf_20_port, B2 => n244, Z => n583);
   U1410 : AOI22D1 port map( A1 => out_buf_212_port, A2 => n270, B1 => 
                           out_buf_148_port, B2 => n245, Z => n582);
   U1411 : AOI22D1 port map( A1 => out_buf_116_port, A2 => n689, B1 => 
                           out_buf_52_port, B2 => n688, Z => n581);
   U1412 : AOI22D1 port map( A1 => out_buf_244_port, A2 => n691, B1 => 
                           out_buf_180_port, B2 => n690, Z => n580);
   U1413 : NAN4D1 port map( A1 => n583, A2 => n582, A3 => n581, A4 => n580, Z 
                           => N2878);
   U1414 : AOI22D1 port map( A1 => out_buf_85_port, A2 => n269, B1 => 
                           out_buf_21_port, B2 => n244, Z => n587);
   U1415 : AOI22D1 port map( A1 => out_buf_213_port, A2 => n270, B1 => 
                           out_buf_149_port, B2 => n245, Z => n586);
   U1416 : AOI22D1 port map( A1 => out_buf_117_port, A2 => n689, B1 => 
                           out_buf_53_port, B2 => n688, Z => n585);
   U1417 : AOI22D1 port map( A1 => out_buf_245_port, A2 => n691, B1 => 
                           out_buf_181_port, B2 => n690, Z => n584);
   U1418 : NAN4D1 port map( A1 => n587, A2 => n586, A3 => n585, A4 => n584, Z 
                           => N2877);
   U1419 : AOI22D1 port map( A1 => out_buf_86_port, A2 => n269, B1 => 
                           out_buf_22_port, B2 => n244, Z => n591);
   U1420 : AOI22D1 port map( A1 => out_buf_214_port, A2 => n270, B1 => 
                           out_buf_150_port, B2 => n245, Z => n5901);
   U1421 : AOI22D1 port map( A1 => out_buf_118_port, A2 => n689, B1 => 
                           out_buf_54_port, B2 => n688, Z => n589);
   U1422 : AOI22D1 port map( A1 => out_buf_246_port, A2 => n691, B1 => 
                           out_buf_182_port, B2 => n690, Z => n588);
   U1423 : NAN4D1 port map( A1 => n591, A2 => n5901, A3 => n589, A4 => n588, Z 
                           => N2876);
   U1424 : AOI22D1 port map( A1 => out_buf_87_port, A2 => n269, B1 => 
                           out_buf_23_port, B2 => n244, Z => n595);
   U1425 : AOI22D1 port map( A1 => out_buf_215_port, A2 => n270, B1 => 
                           out_buf_151_port, B2 => n245, Z => n594);
   U1426 : AOI22D1 port map( A1 => out_buf_119_port, A2 => n689, B1 => 
                           out_buf_55_port, B2 => n688, Z => n593);
   U1427 : AOI22D1 port map( A1 => out_buf_247_port, A2 => n691, B1 => 
                           out_buf_183_port, B2 => n690, Z => n592);
   U1428 : NAN4D1 port map( A1 => n595, A2 => n594, A3 => n593, A4 => n592, Z 
                           => N2875);
   U1429 : AOI22D1 port map( A1 => out_buf_88_port, A2 => n269, B1 => 
                           out_buf_24_port, B2 => n244, Z => n599);
   U1430 : AOI22D1 port map( A1 => out_buf_216_port, A2 => n270, B1 => 
                           out_buf_152_port, B2 => n245, Z => n598);
   U1431 : AOI22D1 port map( A1 => out_buf_120_port, A2 => n689, B1 => 
                           out_buf_56_port, B2 => n688, Z => n597);
   U1432 : AOI22D1 port map( A1 => out_buf_248_port, A2 => n691, B1 => 
                           out_buf_184_port, B2 => n690, Z => n596);
   U1433 : NAN4D1 port map( A1 => n599, A2 => n598, A3 => n597, A4 => n596, Z 
                           => N2874);
   U1434 : AOI22D1 port map( A1 => out_buf_89_port, A2 => n269, B1 => 
                           out_buf_25_port, B2 => n244, Z => n603);
   U1435 : AOI22D1 port map( A1 => out_buf_217_port, A2 => n270, B1 => 
                           out_buf_153_port, B2 => n245, Z => n602);
   U1436 : AOI22D1 port map( A1 => out_buf_121_port, A2 => n689, B1 => 
                           out_buf_57_port, B2 => n688, Z => n601);
   U1437 : AOI22D1 port map( A1 => out_buf_249_port, A2 => n691, B1 => 
                           out_buf_185_port, B2 => n690, Z => n6001);
   U1438 : NAN4D1 port map( A1 => n603, A2 => n602, A3 => n601, A4 => n6001, Z 
                           => N2873);
   U1439 : AOI22D1 port map( A1 => out_buf_90_port, A2 => n269, B1 => 
                           out_buf_26_port, B2 => n244, Z => n607);
   U1440 : AOI22D1 port map( A1 => out_buf_218_port, A2 => n270, B1 => 
                           out_buf_154_port, B2 => n245, Z => n606);
   U1441 : AOI22D1 port map( A1 => out_buf_122_port, A2 => n689, B1 => 
                           out_buf_58_port, B2 => n688, Z => n605);
   U1442 : AOI22D1 port map( A1 => out_buf_250_port, A2 => n691, B1 => 
                           out_buf_186_port, B2 => n690, Z => n604);
   U1443 : NAN4D1 port map( A1 => n607, A2 => n606, A3 => n605, A4 => n604, Z 
                           => N2872);
   U1444 : AOI22D1 port map( A1 => out_buf_91_port, A2 => n269, B1 => 
                           out_buf_27_port, B2 => n244, Z => n611);
   U1445 : AOI22D1 port map( A1 => out_buf_219_port, A2 => n270, B1 => 
                           out_buf_155_port, B2 => n245, Z => n6101);
   U1446 : AOI22D1 port map( A1 => out_buf_123_port, A2 => n689, B1 => 
                           out_buf_59_port, B2 => n688, Z => n609);
   U1447 : AOI22D1 port map( A1 => out_buf_251_port, A2 => n691, B1 => 
                           out_buf_187_port, B2 => n690, Z => n608);
   U1448 : NAN4D1 port map( A1 => n611, A2 => n6101, A3 => n609, A4 => n608, Z 
                           => N2871);
   U1449 : AOI22D1 port map( A1 => out_buf_92_port, A2 => n269, B1 => 
                           out_buf_28_port, B2 => n244, Z => n615);
   U1450 : AOI22D1 port map( A1 => out_buf_220_port, A2 => n270, B1 => 
                           out_buf_156_port, B2 => n245, Z => n614);
   U1451 : AOI22D1 port map( A1 => out_buf_124_port, A2 => n689, B1 => 
                           out_buf_60_port, B2 => n688, Z => n613);
   U1452 : AOI22D1 port map( A1 => out_buf_252_port, A2 => n691, B1 => 
                           out_buf_188_port, B2 => n690, Z => n612);
   U1453 : NAN4D1 port map( A1 => n615, A2 => n614, A3 => n613, A4 => n612, Z 
                           => N2870);
   U1454 : AOI22D1 port map( A1 => out_buf_93_port, A2 => n269, B1 => 
                           out_buf_29_port, B2 => n244, Z => n619);
   U1455 : AOI22D1 port map( A1 => out_buf_221_port, A2 => n270, B1 => 
                           out_buf_157_port, B2 => n245, Z => n618);
   U1456 : AOI22D1 port map( A1 => out_buf_125_port, A2 => n689, B1 => 
                           out_buf_61_port, B2 => n688, Z => n617);
   U1457 : AOI22D1 port map( A1 => out_buf_253_port, A2 => n691, B1 => 
                           out_buf_189_port, B2 => n690, Z => n616);
   U1458 : NAN4D1 port map( A1 => n619, A2 => n618, A3 => n617, A4 => n616, Z 
                           => N2869);
   U1459 : AOI22D1 port map( A1 => out_buf_94_port, A2 => n269, B1 => 
                           out_buf_30_port, B2 => n244, Z => n623);
   U1460 : AOI22D1 port map( A1 => out_buf_222_port, A2 => n270, B1 => 
                           out_buf_158_port, B2 => n245, Z => n622);
   U1461 : AOI22D1 port map( A1 => out_buf_126_port, A2 => n689, B1 => 
                           out_buf_62_port, B2 => n688, Z => n621);
   U1462 : AOI22D1 port map( A1 => out_buf_254_port, A2 => n691, B1 => 
                           out_buf_190_port, B2 => n690, Z => n620);
   U1463 : NAN4D1 port map( A1 => n623, A2 => n622, A3 => n621, A4 => n620, Z 
                           => N2868);
   U1464 : AOI22D1 port map( A1 => out_buf_95_port, A2 => n269, B1 => 
                           out_buf_31_port, B2 => n244, Z => n627);
   U1465 : AOI22D1 port map( A1 => out_buf_223_port, A2 => n270, B1 => 
                           out_buf_159_port, B2 => n245, Z => n626);
   U1466 : AOI22D1 port map( A1 => out_buf_127_port, A2 => n689, B1 => 
                           out_buf_63_port, B2 => n688, Z => n625);
   U1467 : AOI22D1 port map( A1 => out_buf_255_port, A2 => n691, B1 => 
                           out_buf_191_port, B2 => n690, Z => n624);
   U1468 : NAN4D1 port map( A1 => n627, A2 => n626, A3 => n625, A4 => n624, Z 
                           => N2867);
   U1469 : AOI22D1 port map( A1 => out_buf_64_port, A2 => n269, B1 => 
                           out_buf_0_port, B2 => n244, Z => n631);
   U1470 : AOI22D1 port map( A1 => out_buf_192_port, A2 => n270, B1 => 
                           out_buf_128_port, B2 => n245, Z => n6301);
   U1471 : AOI22D1 port map( A1 => out_buf_96_port, A2 => n689, B1 => 
                           out_buf_32_port, B2 => n688, Z => n629);
   U1472 : AOI22D1 port map( A1 => out_buf_224_port, A2 => n691, B1 => 
                           out_buf_160_port, B2 => n690, Z => n628);
   U1473 : NAN4D1 port map( A1 => n631, A2 => n6301, A3 => n629, A4 => n628, Z 
                           => N2865);
   U1474 : AOI22D1 port map( A1 => out_buf_65_port, A2 => n269, B1 => 
                           out_buf_1_port, B2 => n244, Z => n635);
   U1475 : AOI22D1 port map( A1 => out_buf_193_port, A2 => n270, B1 => 
                           out_buf_129_port, B2 => n245, Z => n634);
   U1476 : AOI22D1 port map( A1 => out_buf_97_port, A2 => n689, B1 => 
                           out_buf_33_port, B2 => n688, Z => n633);
   U1477 : AOI22D1 port map( A1 => out_buf_225_port, A2 => n691, B1 => 
                           out_buf_161_port, B2 => n690, Z => n632);
   U1478 : NAN4D1 port map( A1 => n635, A2 => n634, A3 => n633, A4 => n632, Z 
                           => N2864);
   U1479 : AOI22D1 port map( A1 => out_buf_66_port, A2 => n269, B1 => 
                           out_buf_2_port, B2 => n244, Z => n639);
   U1480 : AOI22D1 port map( A1 => out_buf_194_port, A2 => n270, B1 => 
                           out_buf_130_port, B2 => n245, Z => n638);
   U1481 : AOI22D1 port map( A1 => out_buf_98_port, A2 => n689, B1 => 
                           out_buf_34_port, B2 => n688, Z => n637);
   U1482 : AOI22D1 port map( A1 => out_buf_226_port, A2 => n691, B1 => 
                           out_buf_162_port, B2 => n690, Z => n636);
   U1483 : NAN4D1 port map( A1 => n639, A2 => n638, A3 => n637, A4 => n636, Z 
                           => N2863);
   U1484 : AOI22D1 port map( A1 => out_buf_67_port, A2 => n269, B1 => 
                           out_buf_3_port, B2 => n244, Z => n643);
   U1485 : AOI22D1 port map( A1 => out_buf_195_port, A2 => n270, B1 => 
                           out_buf_131_port, B2 => n245, Z => n642);
   U1486 : AOI22D1 port map( A1 => out_buf_99_port, A2 => n689, B1 => 
                           out_buf_35_port, B2 => n688, Z => n641);
   U1487 : AOI22D1 port map( A1 => out_buf_227_port, A2 => n691, B1 => 
                           out_buf_163_port, B2 => n690, Z => n6401);
   U1488 : NAN4D1 port map( A1 => n643, A2 => n642, A3 => n641, A4 => n6401, Z 
                           => N2862);
   U1489 : AOI22D1 port map( A1 => out_buf_68_port, A2 => n269, B1 => 
                           out_buf_4_port, B2 => n244, Z => n647);
   U1490 : AOI22D1 port map( A1 => out_buf_196_port, A2 => n270, B1 => 
                           out_buf_132_port, B2 => n245, Z => n646);
   U1491 : AOI22D1 port map( A1 => out_buf_100_port, A2 => n689, B1 => 
                           out_buf_36_port, B2 => n688, Z => n645);
   U1492 : AOI22D1 port map( A1 => out_buf_228_port, A2 => n691, B1 => 
                           out_buf_164_port, B2 => n690, Z => n644);
   U1493 : NAN4D1 port map( A1 => n647, A2 => n646, A3 => n645, A4 => n644, Z 
                           => N2861);
   U1494 : AOI22D1 port map( A1 => out_buf_69_port, A2 => n269, B1 => 
                           out_buf_5_port, B2 => n244, Z => n651);
   U1495 : AOI22D1 port map( A1 => out_buf_197_port, A2 => n270, B1 => 
                           out_buf_133_port, B2 => n245, Z => n650);
   U1496 : AOI22D1 port map( A1 => out_buf_101_port, A2 => n689, B1 => 
                           out_buf_37_port, B2 => n688, Z => n649);
   U1497 : AOI22D1 port map( A1 => out_buf_229_port, A2 => n691, B1 => 
                           out_buf_165_port, B2 => n690, Z => n648);
   U1498 : NAN4D1 port map( A1 => n651, A2 => n650, A3 => n649, A4 => n648, Z 
                           => N2860);
   U1499 : AOI22D1 port map( A1 => out_buf_70_port, A2 => n269, B1 => 
                           out_buf_6_port, B2 => n244, Z => n655);
   U1500 : AOI22D1 port map( A1 => out_buf_198_port, A2 => n270, B1 => 
                           out_buf_134_port, B2 => n245, Z => n654);
   U1501 : AOI22D1 port map( A1 => out_buf_102_port, A2 => n689, B1 => 
                           out_buf_38_port, B2 => n688, Z => n653);
   U1502 : AOI22D1 port map( A1 => out_buf_230_port, A2 => n691, B1 => 
                           out_buf_166_port, B2 => n690, Z => n652);
   U1503 : NAN4D1 port map( A1 => n655, A2 => n654, A3 => n653, A4 => n652, Z 
                           => N2859);
   U1504 : AOI22D1 port map( A1 => out_buf_71_port, A2 => n269, B1 => 
                           out_buf_7_port, B2 => n244, Z => n659);
   U1505 : AOI22D1 port map( A1 => out_buf_199_port, A2 => n270, B1 => 
                           out_buf_135_port, B2 => n245, Z => n658);
   U1506 : AOI22D1 port map( A1 => out_buf_103_port, A2 => n689, B1 => 
                           out_buf_39_port, B2 => n688, Z => n657);
   U1507 : AOI22D1 port map( A1 => out_buf_231_port, A2 => n691, B1 => 
                           out_buf_167_port, B2 => n690, Z => n656);
   U1508 : NAN4D1 port map( A1 => n659, A2 => n658, A3 => n657, A4 => n656, Z 
                           => N2858);
   U1509 : AOI22D1 port map( A1 => out_buf_72_port, A2 => n269, B1 => 
                           out_buf_8_port, B2 => n244, Z => n663);
   U1510 : AOI22D1 port map( A1 => out_buf_200_port, A2 => n270, B1 => 
                           out_buf_136_port, B2 => n245, Z => n662);
   U1511 : AOI22D1 port map( A1 => out_buf_104_port, A2 => n689, B1 => 
                           out_buf_40_port, B2 => n688, Z => n661);
   U1512 : AOI22D1 port map( A1 => out_buf_232_port, A2 => n691, B1 => 
                           out_buf_168_port, B2 => n690, Z => n660);
   U1513 : NAN4D1 port map( A1 => n663, A2 => n662, A3 => n661, A4 => n660, Z 
                           => N2857);
   U1514 : AOI22D1 port map( A1 => out_buf_73_port, A2 => n269, B1 => 
                           out_buf_9_port, B2 => n244, Z => n667);
   U1515 : AOI22D1 port map( A1 => out_buf_201_port, A2 => n270, B1 => 
                           out_buf_137_port, B2 => n245, Z => n666);
   U1516 : AOI22D1 port map( A1 => out_buf_105_port, A2 => n689, B1 => 
                           out_buf_41_port, B2 => n688, Z => n665);
   U1517 : AOI22D1 port map( A1 => out_buf_233_port, A2 => n691, B1 => 
                           out_buf_169_port, B2 => n690, Z => n664);
   U1518 : NAN4D1 port map( A1 => n667, A2 => n666, A3 => n665, A4 => n664, Z 
                           => N2856);
   U1519 : AOI22D1 port map( A1 => out_buf_74_port, A2 => n269, B1 => 
                           out_buf_10_port, B2 => n244, Z => n671);
   U1520 : AOI22D1 port map( A1 => out_buf_202_port, A2 => n270, B1 => 
                           out_buf_138_port, B2 => n245, Z => n670);
   U1521 : AOI22D1 port map( A1 => out_buf_106_port, A2 => n689, B1 => 
                           out_buf_42_port, B2 => n688, Z => n669);
   U1522 : AOI22D1 port map( A1 => out_buf_234_port, A2 => n691, B1 => 
                           out_buf_170_port, B2 => n690, Z => n668);
   U1523 : NAN4D1 port map( A1 => n671, A2 => n670, A3 => n669, A4 => n668, Z 
                           => N2855);
   U1524 : AOI22D1 port map( A1 => out_buf_75_port, A2 => n269, B1 => 
                           out_buf_11_port, B2 => n244, Z => n675);
   U1525 : AOI22D1 port map( A1 => out_buf_203_port, A2 => n270, B1 => 
                           out_buf_139_port, B2 => n245, Z => n674);
   U1526 : AOI22D1 port map( A1 => out_buf_107_port, A2 => n689, B1 => 
                           out_buf_43_port, B2 => n688, Z => n673);
   U1527 : AOI22D1 port map( A1 => out_buf_235_port, A2 => n691, B1 => 
                           out_buf_171_port, B2 => n690, Z => n672);
   U1528 : NAN4D1 port map( A1 => n675, A2 => n674, A3 => n673, A4 => n672, Z 
                           => N2854);
   U1529 : AOI22D1 port map( A1 => out_buf_76_port, A2 => n269, B1 => 
                           out_buf_12_port, B2 => n244, Z => n679);
   U1530 : AOI22D1 port map( A1 => out_buf_204_port, A2 => n270, B1 => 
                           out_buf_140_port, B2 => n245, Z => n678);
   U1531 : AOI22D1 port map( A1 => out_buf_108_port, A2 => n689, B1 => 
                           out_buf_44_port, B2 => n688, Z => n677);
   U1532 : AOI22D1 port map( A1 => out_buf_236_port, A2 => n691, B1 => 
                           out_buf_172_port, B2 => n690, Z => n676);
   U1533 : NAN4D1 port map( A1 => n679, A2 => n678, A3 => n677, A4 => n676, Z 
                           => N2853);
   U1534 : AOI22D1 port map( A1 => out_buf_77_port, A2 => n269, B1 => 
                           out_buf_13_port, B2 => n244, Z => n683);
   U1535 : AOI22D1 port map( A1 => out_buf_205_port, A2 => n270, B1 => 
                           out_buf_141_port, B2 => n245, Z => n682);
   U1536 : AOI22D1 port map( A1 => out_buf_109_port, A2 => n689, B1 => 
                           out_buf_45_port, B2 => n688, Z => n681);
   U1537 : AOI22D1 port map( A1 => out_buf_237_port, A2 => n691, B1 => 
                           out_buf_173_port, B2 => n690, Z => n680);
   U1538 : NAN4D1 port map( A1 => n683, A2 => n682, A3 => n681, A4 => n680, Z 
                           => N2852);
   U1539 : AOI22D1 port map( A1 => out_buf_78_port, A2 => n269, B1 => 
                           out_buf_14_port, B2 => n244, Z => n687);
   U1540 : AOI22D1 port map( A1 => out_buf_206_port, A2 => n270, B1 => 
                           out_buf_142_port, B2 => n245, Z => n686);
   U1541 : AOI22D1 port map( A1 => out_buf_110_port, A2 => n689, B1 => 
                           out_buf_46_port, B2 => n688, Z => n685);
   U1542 : AOI22D1 port map( A1 => out_buf_238_port, A2 => n691, B1 => 
                           out_buf_174_port, B2 => n690, Z => n684);
   U1543 : NAN4D1 port map( A1 => n687, A2 => n686, A3 => n685, A4 => n684, Z 
                           => N2851);
   U1544 : AOI22D1 port map( A1 => out_buf_79_port, A2 => n269, B1 => 
                           out_buf_15_port, B2 => n244, Z => n695);
   U1545 : AOI22D1 port map( A1 => out_buf_207_port, A2 => n270, B1 => 
                           out_buf_143_port, B2 => n245, Z => n694);
   U1546 : AOI22D1 port map( A1 => out_buf_111_port, A2 => n689, B1 => 
                           out_buf_47_port, B2 => n688, Z => n693);
   U1547 : AOI22D1 port map( A1 => out_buf_239_port, A2 => n691, B1 => 
                           out_buf_175_port, B2 => n690, Z => n692);
   U1548 : NAN4D1 port map( A1 => n695, A2 => n694, A3 => n693, A4 => n692, Z 
                           => N2850);
   U1549 : NAN2D1 port map( A1 => n114, A2 => avs_addr(3), Z => n6400);
   U1550 : NAN3D1 port map( A1 => avs_write, A2 => n277, A3 => n795, Z => n178)
                           ;
   U1551 : NAN2D1 port map( A1 => operand_regs_255_port, A2 => n709, Z => n763)
                           ;
   U1552 : OAI21D1 port map( A1 => n713, A2 => n730, B => n763, Z => N3104);
   U1553 : NAN2D1 port map( A1 => operand_regs_254_port, A2 => n709, Z => n764)
                           ;
   U1554 : OAI21D1 port map( A1 => n706, A2 => n731, B => n764, Z => N3103);
   U1555 : NAN2D1 port map( A1 => operand_regs_253_port, A2 => n709, Z => n765)
                           ;
   U1556 : OAI21D1 port map( A1 => n708, A2 => n732, B => n765, Z => N3102);
   U1557 : NAN2D1 port map( A1 => operand_regs_252_port, A2 => n709, Z => n766)
                           ;
   U1558 : OAI21D1 port map( A1 => n706, A2 => n733, B => n766, Z => N3101);
   U1559 : NAN2D1 port map( A1 => operand_regs_251_port, A2 => n709, Z => n767)
                           ;
   U1560 : OAI21D1 port map( A1 => n706, A2 => n734, B => n767, Z => N3100);
   U1561 : NAN2D1 port map( A1 => operand_regs_250_port, A2 => n709, Z => n768)
                           ;
   U1562 : OAI21D1 port map( A1 => n713, A2 => n735, B => n768, Z => N3099);
   U1563 : NAN2D1 port map( A1 => operand_regs_249_port, A2 => n709, Z => n769)
                           ;
   U1564 : OAI21D1 port map( A1 => n707, A2 => n736, B => n769, Z => N3098);
   U1565 : NAN2D1 port map( A1 => operand_regs_248_port, A2 => n709, Z => n770)
                           ;
   U1566 : OAI21D1 port map( A1 => n708, A2 => n737, B => n770, Z => N3097);
   U1567 : NAN2D1 port map( A1 => operand_regs_247_port, A2 => n709, Z => n771)
                           ;
   U1568 : OAI21D1 port map( A1 => n707, A2 => n738, B => n771, Z => N3096);
   U1569 : NAN2D1 port map( A1 => operand_regs_246_port, A2 => n709, Z => n772)
                           ;
   U1570 : OAI21D1 port map( A1 => n713, A2 => n739, B => n772, Z => N3095);
   U1571 : NAN2D1 port map( A1 => operand_regs_245_port, A2 => n709, Z => n773)
                           ;
   U1572 : OAI21D1 port map( A1 => n707, A2 => n740, B => n773, Z => N3094);
   U1573 : NAN2D1 port map( A1 => operand_regs_244_port, A2 => n708, Z => n774)
                           ;
   U1574 : OAI21D1 port map( A1 => n707, A2 => n741, B => n774, Z => N3093);
   U1575 : NAN2D1 port map( A1 => operand_regs_243_port, A2 => n708, Z => n775)
                           ;
   U1576 : OAI21D1 port map( A1 => n707, A2 => n742, B => n775, Z => N3092);
   U1577 : NAN2D1 port map( A1 => operand_regs_242_port, A2 => n708, Z => n776)
                           ;
   U1578 : OAI21D1 port map( A1 => n707, A2 => n743, B => n776, Z => N3091);
   U1579 : NAN2D1 port map( A1 => operand_regs_241_port, A2 => n708, Z => n777)
                           ;
   U1580 : OAI21D1 port map( A1 => n708, A2 => n744, B => n777, Z => N3090);
   U1581 : NAN2D1 port map( A1 => operand_regs_240_port, A2 => n708, Z => n778)
                           ;
   U1582 : OAI21D1 port map( A1 => n706, A2 => n745, B => n778, Z => N3089);
   U1583 : NAN2D1 port map( A1 => operand_regs_239_port, A2 => n708, Z => n779)
                           ;
   U1584 : OAI21D1 port map( A1 => n708, A2 => n746, B => n779, Z => N3088);
   U1585 : NAN2D1 port map( A1 => operand_regs_238_port, A2 => n708, Z => n780)
                           ;
   U1586 : OAI21D1 port map( A1 => n706, A2 => n747, B => n780, Z => N3087);
   U1587 : NAN2D1 port map( A1 => operand_regs_237_port, A2 => n708, Z => n781)
                           ;
   U1588 : OAI21D1 port map( A1 => n708, A2 => n748, B => n781, Z => N3086);
   U1589 : NAN2D1 port map( A1 => operand_regs_236_port, A2 => n707, Z => n782)
                           ;
   U1590 : OAI21D1 port map( A1 => n708, A2 => n749, B => n782, Z => N3085);
   U1591 : NAN2D1 port map( A1 => operand_regs_235_port, A2 => n708, Z => n783)
                           ;
   U1592 : OAI21D1 port map( A1 => n713, A2 => n750, B => n783, Z => N3084);
   U1593 : NAN2D1 port map( A1 => operand_regs_234_port, A2 => n708, Z => n784)
                           ;
   U1594 : OAI21D1 port map( A1 => n708, A2 => n751, B => n784, Z => N3083);
   U1595 : NAN2D1 port map( A1 => operand_regs_233_port, A2 => n708, Z => n785)
                           ;
   U1596 : OAI21D1 port map( A1 => n713, A2 => n752, B => n785, Z => N3082);
   U1597 : NAN2D1 port map( A1 => operand_regs_232_port, A2 => n707, Z => n786)
                           ;
   U1598 : OAI21D1 port map( A1 => n708, A2 => n753, B => n786, Z => N3081);
   U1599 : NAN2D1 port map( A1 => operand_regs_231_port, A2 => n708, Z => n787)
                           ;
   U1600 : OAI21D1 port map( A1 => n706, A2 => n754, B => n787, Z => N3080);
   U1601 : NAN2D1 port map( A1 => operand_regs_230_port, A2 => n707, Z => n788)
                           ;
   U1602 : OAI21D1 port map( A1 => n706, A2 => n755, B => n788, Z => N3079);
   U1603 : NAN2D1 port map( A1 => operand_regs_229_port, A2 => n708, Z => n789)
                           ;
   U1604 : OAI21D1 port map( A1 => n706, A2 => n756, B => n789, Z => N3078);
   U1605 : NAN2D1 port map( A1 => operand_regs_228_port, A2 => n707, Z => n790)
                           ;
   U1606 : OAI21D1 port map( A1 => n706, A2 => n757, B => n790, Z => N3077);
   U1607 : NAN2D1 port map( A1 => operand_regs_227_port, A2 => n707, Z => n791)
                           ;
   U1608 : OAI21D1 port map( A1 => n706, A2 => n758, B => n791, Z => N3076);
   U1609 : NAN2D1 port map( A1 => operand_regs_226_port, A2 => n708, Z => n792)
                           ;
   U1610 : OAI21D1 port map( A1 => n706, A2 => n759, B => n792, Z => N3075);
   U1611 : NAN2D1 port map( A1 => operand_regs_225_port, A2 => n707, Z => n793)
                           ;
   U1612 : OAI21D1 port map( A1 => n706, A2 => n760, B => n793, Z => N3074);
   U1613 : NAN2D1 port map( A1 => operand_regs_224_port, A2 => n707, Z => n794)
                           ;
   U1614 : OAI21D1 port map( A1 => n706, A2 => n761, B => n794, Z => N3073);
   U1615 : OAI21M20D1 port map( A1 => operand_regs_159_port, A2 => n726, B => 
                           n763, Z => N3136);
   U1616 : OAI21M20D1 port map( A1 => operand_regs_158_port, A2 => n726, B => 
                           n764, Z => N3135);
   U1617 : OAI21M20D1 port map( A1 => operand_regs_157_port, A2 => n726, B => 
                           n765, Z => N3134);
   U1618 : OAI21M20D1 port map( A1 => operand_regs_156_port, A2 => n726, B => 
                           n766, Z => N3133);
   U1619 : OAI21M20D1 port map( A1 => operand_regs_155_port, A2 => n726, B => 
                           n767, Z => N3132);
   U1620 : OAI21M20D1 port map( A1 => operand_regs_154_port, A2 => n728, B => 
                           n768, Z => N3131);
   U1621 : OAI21M20D1 port map( A1 => operand_regs_153_port, A2 => n728, B => 
                           n769, Z => N3130);
   U1622 : OAI21M20D1 port map( A1 => operand_regs_152_port, A2 => n728, B => 
                           n770, Z => N3129);
   U1623 : OAI21M20D1 port map( A1 => operand_regs_151_port, A2 => n728, B => 
                           n771, Z => N3128);
   U1624 : OAI21M20D1 port map( A1 => operand_regs_150_port, A2 => n727, B => 
                           n772, Z => N3127);
   U1625 : OAI21M20D1 port map( A1 => operand_regs_149_port, A2 => n728, B => 
                           n773, Z => N3126);
   U1626 : OAI21M20D1 port map( A1 => operand_regs_148_port, A2 => n728, B => 
                           n774, Z => N3125);
   U1627 : OAI21M20D1 port map( A1 => operand_regs_147_port, A2 => n727, B => 
                           n775, Z => N3124);
   U1628 : OAI21M20D1 port map( A1 => operand_regs_146_port, A2 => n727, B => 
                           n776, Z => N3123);
   U1629 : OAI21M20D1 port map( A1 => operand_regs_145_port, A2 => n727, B => 
                           n777, Z => N3122);
   U1630 : OAI21M20D1 port map( A1 => operand_regs_144_port, A2 => n728, B => 
                           n778, Z => N3121);
   U1631 : OAI21M20D1 port map( A1 => operand_regs_143_port, A2 => n727, B => 
                           n779, Z => N3120);
   U1632 : OAI21M20D1 port map( A1 => operand_regs_142_port, A2 => n727, B => 
                           n780, Z => N3119);
   U1633 : OAI21M20D1 port map( A1 => operand_regs_141_port, A2 => n728, B => 
                           n781, Z => N3118);
   U1634 : OAI21M20D1 port map( A1 => operand_regs_140_port, A2 => n727, B => 
                           n782, Z => N3117);
   U1635 : OAI21M20D1 port map( A1 => operand_regs_139_port, A2 => n728, B => 
                           n783, Z => N3116);
   U1636 : OAI21M20D1 port map( A1 => operand_regs_138_port, A2 => n727, B => 
                           n784, Z => N3115);
   U1637 : OAI21M20D1 port map( A1 => operand_regs_137_port, A2 => n728, B => 
                           n785, Z => N3114);
   U1638 : OAI21M20D1 port map( A1 => operand_regs_136_port, A2 => n727, B => 
                           n786, Z => N3113);
   U1639 : OAI21M20D1 port map( A1 => operand_regs_135_port, A2 => n727, B => 
                           n787, Z => N3112);
   U1640 : OAI21M20D1 port map( A1 => operand_regs_134_port, A2 => n727, B => 
                           n788, Z => N3111);
   U1641 : OAI21M20D1 port map( A1 => operand_regs_133_port, A2 => n727, B => 
                           n789, Z => N3110);
   U1642 : OAI21M20D1 port map( A1 => operand_regs_132_port, A2 => n727, B => 
                           n790, Z => N3109);
   U1643 : OAI21M20D1 port map( A1 => operand_regs_131_port, A2 => n727, B => 
                           n791, Z => N3108);
   U1644 : OAI21M20D1 port map( A1 => operand_regs_130_port, A2 => n727, B => 
                           n792, Z => N3107);
   U1645 : OAI21M20D1 port map( A1 => operand_regs_129_port, A2 => n727, B => 
                           n793, Z => N3106);
   U1646 : OAI21M20D1 port map( A1 => operand_regs_128_port, A2 => n727, B => 
                           n794, Z => N3105);
   U1647 : OAI21M20D1 port map( A1 => operand_regs_95_port, A2 => n728, B => 
                           n763, Z => N3168);
   U1648 : OAI21M20D1 port map( A1 => operand_regs_94_port, A2 => n727, B => 
                           n764, Z => N3167);
   U1649 : OAI21M20D1 port map( A1 => operand_regs_93_port, A2 => n728, B => 
                           n765, Z => N3166);
   U1650 : OAI21M20D1 port map( A1 => operand_regs_92_port, A2 => n727, B => 
                           n766, Z => N3165);
   U1651 : OAI21M20D1 port map( A1 => operand_regs_91_port, A2 => n728, B => 
                           n767, Z => N3164);
   U1652 : OAI21M20D1 port map( A1 => operand_regs_90_port, A2 => n728, B => 
                           n768, Z => N3163);
   U1653 : OAI21M20D1 port map( A1 => operand_regs_89_port, A2 => n727, B => 
                           n769, Z => N3162);
   U1654 : OAI21M20D1 port map( A1 => operand_regs_88_port, A2 => n727, B => 
                           n770, Z => N3161);
   U1655 : OAI21M20D1 port map( A1 => operand_regs_87_port, A2 => n728, B => 
                           n771, Z => N3160);
   U1656 : OAI21M20D1 port map( A1 => operand_regs_86_port, A2 => n728, B => 
                           n772, Z => N3159);
   U1657 : OAI21M20D1 port map( A1 => operand_regs_85_port, A2 => n727, B => 
                           n773, Z => N3158);
   U1658 : OAI21M20D1 port map( A1 => operand_regs_84_port, A2 => n728, B => 
                           n774, Z => N3157);
   U1659 : OAI21M20D1 port map( A1 => operand_regs_83_port, A2 => n727, B => 
                           n775, Z => N3156);
   U1660 : OAI21M20D1 port map( A1 => operand_regs_82_port, A2 => n727, B => 
                           n776, Z => N3155);
   U1661 : OAI21M20D1 port map( A1 => operand_regs_81_port, A2 => n727, B => 
                           n777, Z => N3154);
   U1662 : OAI21M20D1 port map( A1 => operand_regs_80_port, A2 => n727, B => 
                           n778, Z => N3153);
   U1663 : OAI21M20D1 port map( A1 => operand_regs_79_port, A2 => n727, B => 
                           n779, Z => N3152);
   U1664 : OAI21M20D1 port map( A1 => operand_regs_78_port, A2 => n727, B => 
                           n780, Z => N3151);
   U1665 : OAI21M20D1 port map( A1 => operand_regs_77_port, A2 => n727, B => 
                           n781, Z => N3150);
   U1666 : OAI21M20D1 port map( A1 => operand_regs_76_port, A2 => n727, B => 
                           n782, Z => N3149);
   U1667 : OAI21M20D1 port map( A1 => operand_regs_75_port, A2 => n727, B => 
                           n783, Z => N3148);
   U1668 : OAI21M20D1 port map( A1 => operand_regs_74_port, A2 => n727, B => 
                           n784, Z => N3147);
   U1669 : OAI21M20D1 port map( A1 => operand_regs_73_port, A2 => n727, B => 
                           n785, Z => N3146);
   U1670 : OAI21M20D1 port map( A1 => operand_regs_72_port, A2 => n727, B => 
                           n786, Z => N3145);
   U1671 : OAI21M20D1 port map( A1 => operand_regs_71_port, A2 => n727, B => 
                           n787, Z => N3144);
   U1672 : OAI21M20D1 port map( A1 => operand_regs_70_port, A2 => n728, B => 
                           n788, Z => N3143);
   U1673 : OAI21M20D1 port map( A1 => operand_regs_69_port, A2 => n728, B => 
                           n789, Z => N3142);
   U1674 : OAI21M20D1 port map( A1 => operand_regs_68_port, A2 => n728, B => 
                           n790, Z => N3141);
   U1675 : OAI21M20D1 port map( A1 => operand_regs_67_port, A2 => n728, B => 
                           n791, Z => N3140);
   U1676 : OAI21M20D1 port map( A1 => operand_regs_66_port, A2 => n728, B => 
                           n792, Z => N3139);
   U1677 : OAI21M20D1 port map( A1 => operand_regs_65_port, A2 => n728, B => 
                           n793, Z => N3138);
   U1678 : OAI21M20D1 port map( A1 => operand_regs_64_port, A2 => n728, B => 
                           n794, Z => N3137);
   U1679 : NOR3D1 port map( A1 => avs_addr(3), A2 => avs_addr(5), A3 => 
                           avs_addr(4), Z => N66);

end hier_filter_none_5;
